//
// Conformal-LEC: Version 24.10-s400 (28-Apr-2025) (64 bit executable)
//
module WALLACE_CSA_DUMMY_OP4_group_359292(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, in_85, in_86, out_0);
input  in_47, in_55, in_58, in_76, in_84;
input   [4:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [6:0] in_4;
input   [1:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
input   [2:0] in_41;
input   [1:0] in_42;
input   [1:0] in_43;
input   [4:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [1:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [2:0] in_53;
input   [1:0] in_54;
input   [2:0] in_56;
input   [4:0] in_57;
input   [1:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [1:0] in_62;
input   [4:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [1:0] in_66;
input   [4:0] in_67;
input   [4:0] in_68;
input   [4:0] in_69;
input   [4:0] in_70;
input   [4:0] in_71;
input   [2:0] in_72;
input   [4:0] in_73;
input   [2:0] in_74;
input   [4:0] in_75;
input   [1:0] in_77;
input   [4:0] in_78;
input   [2:0] in_79;
input   [4:0] in_80;
input   [4:0] in_81;
input   [1:0] in_82;
input   [1:0] in_83;
input   [4:0] in_85;
input   [4:0] in_86;
output  [9:0] out_0;
wire  n_274, n_272, n_270, n_268, n_266, n_265, n_264, n_262, n_261, n_260, 
    n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, 
    n_249, n_248, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
    n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_218, 
    n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
    n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, 
    n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, 
    n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, 
    n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, 
    n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_84, 
    in_76, in_58, in_55, in_47;
wire   [9:0] out_0;
wire   [2:0] in_79;
wire   [2:0] in_74;
wire   [2:0] in_72;
wire   [2:0] in_56;
wire   [2:0] in_53;
wire   [2:0] in_41;
wire   [2:0] in_34;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [1:0] in_83;
wire   [1:0] in_82;
wire   [1:0] in_77;
wire   [1:0] in_66;
wire   [1:0] in_62;
wire   [1:0] in_61;
wire   [1:0] in_59;
wire   [1:0] in_54;
wire   [1:0] in_51;
wire   [1:0] in_48;
wire   [1:0] in_43;
wire   [1:0] in_42;
wire   [1:0] in_40;
wire   [1:0] in_36;
wire   [1:0] in_5;
wire   [6:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_86;
wire   [4:0] in_85;
wire   [4:0] in_81;
wire   [4:0] in_80;
wire   [4:0] in_78;
wire   [4:0] in_75;
wire   [4:0] in_73;
wire   [4:0] in_71;
wire   [4:0] in_70;
wire   [4:0] in_69;
wire   [4:0] in_68;
wire   [4:0] in_67;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_63;
wire   [4:0] in_60;
wire   [4:0] in_57;
wire   [4:0] in_52;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g8724(.Y(out_0[9]), .A(n_274));
  ADDFX1 g8725(.CO(n_274), .S(out_0[7]), .A(n_38), .B(n_256), .CI(n_272));
  ADDFX1 g8726(.CO(n_272), .S(out_0[6]), .A(n_257), .B(n_264), .CI(n_270));
  ADDFX1 g8727(.CO(n_270), .S(out_0[5]), .A(n_260), .B(n_265), .CI(n_268));
  ADDFX1 g8728(.CO(n_268), .S(out_0[4]), .A(n_258), .B(n_261), .CI(n_266));
  ADDFX1 g8729(.CO(n_266), .S(out_0[3]), .A(n_252), .B(n_262), .CI(n_259));
  ADDFX1 g8730(.CO(n_264), .S(n_265), .A(n_244), .B(n_254), .CI(n_249));
  ADDFX1 g8731(.CO(n_262), .S(out_0[2]), .A(n_239), .B(n_246), .CI(n_253));
  ADDFX1 g8732(.CO(n_260), .S(n_261), .A(n_250), .B(n_245), .CI(n_255));
  ADDFX1 g8733(.CO(n_258), .S(n_259), .A(n_231), .B(n_251), .CI(n_243));
  ADDFX1 g8734(.CO(n_256), .S(n_257), .A(n_228), .B(n_37), .CI(n_248));
  ADDFX1 g8735(.CO(n_254), .S(n_255), .A(n_235), .B(n_230), .CI(n_242));
  ADDFX1 g8736(.CO(n_252), .S(n_253), .A(n_236), .B(n_227), .CI(n_241));
  ADDFX1 g8737(.CO(n_250), .S(n_251), .A(n_226), .B(n_233), .CI(n_238));
  ADDFX1 g8738(.CO(n_248), .S(n_249), .A(n_204), .B(n_234), .CI(n_229));
  ADDFX1 g8739(.CO(n_246), .S(out_0[1]), .A(n_218), .B(n_237), .CI(n_209));
  ADDFX1 g8740(.CO(n_244), .S(n_245), .A(n_224), .B(n_232), .CI(n_205));
  ADDFX1 g8741(.CO(n_242), .S(n_243), .A(n_220), .B(n_225), .CI(n_240));
  ADDFX1 g8742(.CO(n_240), .S(n_241), .A(n_210), .B(n_202), .CI(n_223));
  ADDFX1 g8743(.CO(n_238), .S(n_239), .A(n_213), .B(n_208), .CI(n_221));
  ADDFX1 g8744(.CO(n_236), .S(n_237), .A(n_181), .B(n_211), .CI(n_203));
  ADDFX1 g8745(.CO(n_234), .S(n_235), .A(n_201), .B(n_216), .CI(n_206));
  ADDFX1 g8746(.CO(n_232), .S(n_233), .A(n_199), .B(n_217), .CI(n_222));
  ADDFX1 g8747(.CO(n_230), .S(n_231), .A(n_212), .B(n_214), .CI(n_207));
  ADDFX1 g8748(.CO(n_228), .S(n_229), .A(n_200), .B(n_0), .CI(in_3[5]));
  ADDFX1 g8749(.CO(n_226), .S(n_227), .A(n_180), .B(n_177), .CI(n_215));
  ADDFX1 g8750(.CO(n_224), .S(n_225), .A(n_178), .B(n_176), .CI(in_2[3]));
  ADDFX1 g8751(.CO(n_222), .S(n_223), .A(n_174), .B(n_196), .CI(in_2[2]));
  ADDFX1 g8752(.CO(n_220), .S(n_221), .A(n_171), .B(n_183), .CI(n_172));
  ADDFX1 g8753(.CO(n_218), .S(out_0[0]), .A(n_195), .B(n_189), .CI(n_127));
  ADDFX1 g8754(.CO(n_216), .S(n_217), .A(n_169), .B(n_184), .CI(n_187));
  ADDFX1 g8755(.CO(n_214), .S(n_215), .A(n_185), .B(n_192), .CI(in_3[2]));
  ADDFX1 g8756(.CO(n_212), .S(n_213), .A(n_167), .B(n_190), .CI(n_179));
  ADDFX1 g8757(.CO(n_210), .S(n_211), .A(n_197), .B(n_193), .CI(n_188));
  ADDFX1 g8758(.CO(n_208), .S(n_209), .A(n_194), .B(n_191), .CI(n_173));
  ADDFX1 g8759(.CO(n_206), .S(n_207), .A(n_170), .B(n_182), .CI(in_3[3]));
  ADDFX1 g8760(.CO(n_204), .S(n_205), .A(n_198), .B(in_2[4]), .CI(in_3[4]));
  ADDFX1 g8761(.CO(n_202), .S(n_203), .A(n_175), .B(in_2[1]), .CI(n_126));
  ADDFX1 g8762(.CO(n_200), .S(n_201), .A(n_114), .B(n_168), .CI(n_186));
  ADDFX1 g8763(.CO(n_198), .S(n_199), .A(n_156), .B(n_124), .CI(n_166));
  ADDFX1 g8764(.CO(n_196), .S(n_197), .A(n_160), .B(n_128), .CI(n_154));
  ADDFX1 g8765(.CO(n_194), .S(n_195), .A(n_129), .B(n_161), .CI(n_163));
  ADDFX1 g8766(.CO(n_192), .S(n_193), .A(n_123), .B(n_133), .CI(n_158));
  ADDFX1 g8767(.CO(n_190), .S(n_191), .A(n_147), .B(n_141), .CI(n_121));
  ADDFX1 g8768(.CO(n_188), .S(n_189), .A(n_159), .B(n_151), .CI(n_155));
  ADDFX1 g8769(.CO(n_186), .S(n_187), .A(n_118), .B(n_142), .CI(n_164));
  ADDFX1 g8770(.CO(n_184), .S(n_185), .A(n_148), .B(n_146), .CI(n_134));
  ADDFX1 g8771(.CO(n_182), .S(n_183), .A(n_143), .B(n_145), .CI(n_165));
  ADDFX1 g8772(.CO(n_180), .S(n_181), .A(n_162), .B(n_153), .CI(n_131));
  ADDFX1 g8773(.CO(n_178), .S(n_179), .A(n_132), .B(n_120), .CI(n_157));
  ADDFX1 g8774(.CO(n_176), .S(n_177), .A(n_152), .B(n_125), .CI(n_130));
  ADDFX1 g8775(.CO(n_174), .S(n_175), .A(n_149), .B(n_135), .CI(n_150));
  ADDFX1 g8776(.CO(n_172), .S(n_173), .A(n_137), .B(n_139), .CI(in_3[1]));
  ADDFX1 g8777(.CO(n_170), .S(n_171), .A(n_140), .B(n_138), .CI(n_136));
  ADDFX1 g8778(.CO(n_168), .S(n_169), .A(n_57), .B(n_115), .CI(n_144));
  ADDFX1 g8779(.CO(n_166), .S(n_167), .A(n_43), .B(n_122), .CI(n_119));
  ADDFX1 g8780(.CO(n_164), .S(n_165), .A(n_71), .B(n_91), .CI(n_89));
  ADDFX1 g8781(.CO(n_162), .S(n_163), .A(n_107), .B(n_102), .CI(n_117));
  ADDFX1 g8782(.CO(n_160), .S(n_161), .A(n_64), .B(n_100), .CI(n_98));
  ADDFX1 g8783(.CO(n_158), .S(n_159), .A(n_88), .B(n_60), .CI(n_86));
  ADDFX1 g8784(.CO(n_156), .S(n_157), .A(n_81), .B(n_113), .CI(n_75));
  ADDFX1 g8785(.CO(n_154), .S(n_155), .A(n_78), .B(n_68), .CI(n_111));
  ADDFX1 g8786(.CO(n_152), .S(n_153), .A(n_72), .B(n_76), .CI(n_116));
  ADDFX1 g8787(.CO(n_150), .S(n_151), .A(in_29[0]), .B(n_84), .CI(n_70));
  ADDFX1 g8788(.CO(n_148), .S(n_149), .A(n_106), .B(n_99), .CI(n_73));
  ADDFX1 g8789(.CO(n_146), .S(n_147), .A(n_30), .B(n_77), .CI(n_59));
  ADDFX1 g8790(.CO(n_144), .S(n_145), .A(n_53), .B(n_41), .CI(n_108));
  ADDFX1 g8791(.CO(n_142), .S(n_143), .A(n_79), .B(n_93), .CI(n_49));
  ADDFX1 g8792(.CO(n_140), .S(n_141), .A(n_69), .B(n_97), .CI(n_95));
  ADDFX1 g8793(.CO(n_138), .S(n_139), .A(n_94), .B(n_104), .CI(n_109));
  ADDFX1 g8794(.CO(n_136), .S(n_137), .A(n_50), .B(n_92), .CI(n_90));
  ADDFX1 g8795(.CO(n_134), .S(n_135), .A(n_67), .B(n_110), .CI(n_101));
  ADDFX1 g8796(.CO(n_132), .S(n_133), .A(n_87), .B(n_85), .CI(n_54));
  ADDFX1 g8797(.CO(n_130), .S(n_131), .A(n_61), .B(n_44), .CI(n_40));
  ADDFX1 g8798(.CO(n_128), .S(n_129), .A(n_96), .B(n_74), .CI(n_48));
  ADDFX1 g8799(.CO(n_126), .S(n_127), .A(n_62), .B(in_3[0]), .CI(in_2[0]));
  ADDFX1 g8800(.CO(n_124), .S(n_125), .A(n_35), .B(n_39), .CI(n_58));
  ADDFX1 g8801(.CO(n_122), .S(n_123), .A(n_63), .B(n_47), .CI(n_83));
  ADDFX1 g8802(.CO(n_120), .S(n_121), .A(n_82), .B(n_42), .CI(n_80));
  ADDFX1 g8803(.CO(n_118), .S(n_119), .A(n_3), .B(n_20), .CI(n_103));
  ADDFX1 g8804(.CO(n_116), .S(n_117), .A(in_14[0]), .B(n_33), .CI(in_13[0]));
  XNOR2X1 g8805(.Y(n_115), .A(n_31), .B(n_112));
  NOR2BX1 g8806(.Y(n_114), .AN(n_31), .B(n_112));
  INVX1 g8807(.Y(n_113), .A(n_105));
  ADDFX1 g8808(.CO(n_110), .S(n_111), .A(in_22[0]), .B(n_5), .CI(in_55));
  ADDFX1 g8809(.CO(n_108), .S(n_109), .A(in_8[1]), .B(n_10), .CI(in_56[0]));
  ADDFX1 g8810(.CO(n_106), .S(n_107), .A(n_1), .B(n_13), .CI(in_82[0]));
  ADDFX1 g8811(.CO(n_112), .S(n_105), .A(in_17[2]), .B(in_24[0]), .CI(in_69[0]));
  ADDFX1 g8812(.CO(n_103), .S(n_104), .A(in_4[1]), .B(in_61[1]), .CI(in_19[1]));
  ADDFX1 g8813(.CO(n_101), .S(n_102), .A(in_51[0]), .B(n_11), .CI(n_27));
  ADDFX1 g8814(.CO(n_99), .S(n_100), .A(in_23[0]), .B(n_28), .CI(n_8));
  ADDFX1 g8815(.CO(n_97), .S(n_98), .A(in_10[0]), .B(in_42[0]), .CI(n_14));
  ADDFX1 g8816(.CO(n_95), .S(n_96), .A(in_24[0]), .B(n_19), .CI(in_69[0]));
  ADDFX1 g8817(.CO(n_93), .S(n_94), .A(in_9[1]), .B(in_42[0]), .CI(n_25));
  ADDFX1 g8818(.CO(n_91), .S(n_92), .A(in_34[1]), .B(in_74[1]), .CI(in_72[1]));
  ADDFX1 g8819(.CO(n_89), .S(n_90), .A(in_48[1]), .B(in_59[1]), .CI(n_29));
  ADDFX1 g8820(.CO(n_87), .S(n_88), .A(in_58), .B(in_43[0]), .CI(in_65[0]));
  ADDFX1 g8821(.CO(n_85), .S(n_86), .A(in_66[0]), .B(n_16), .CI(in_76));
  INVX1 g8822(.Y(n_84), .A(n_66));
  INVX1 g8823(.Y(n_83), .A(n_65));
  INVX1 g8824(.Y(n_82), .A(n_56));
  INVX1 g8825(.Y(n_81), .A(n_55));
  INVX1 g8826(.Y(n_80), .A(n_52));
  INVX1 g8827(.Y(n_79), .A(n_51));
  INVX1 g8828(.Y(n_78), .A(n_46));
  INVX1 g8829(.Y(n_77), .A(n_45));
  ADDFX1 g8830(.CO(n_75), .S(n_76), .A(in_83[1]), .B(n_9), .CI(n_17));
  ADDFX1 g8831(.CO(n_73), .S(n_74), .A(in_15[0]), .B(n_12), .CI(in_84));
  ADDFX1 g8832(.CO(n_71), .S(n_72), .A(n_18), .B(n_2), .CI(in_79[1]));
  ADDFX1 g8833(.CO(n_69), .S(n_70), .A(in_5[0]), .B(in_26[0]), .CI(in_40[0]));
  ADDFX1 g8834(.CO(n_67), .S(n_68), .A(in_18[0]), .B(n_7), .CI(n_26));
  ADDFX1 g8835(.CO(n_65), .S(n_66), .A(in_73[0]), .B(in_20[0]), .CI(in_75[0]));
  ADDFX1 g8836(.CO(n_63), .S(n_64), .A(in_38[0]), .B(in_56[0]), .CI(in_77[0]));
  ADDFX1 g8837(.CO(n_61), .S(n_62), .A(in_19[0]), .B(in_7[0]), .CI(in_27[0]));
  ADDFX1 g8838(.CO(n_59), .S(n_60), .A(in_28[0]), .B(in_4[0]), .CI(in_47));
  ADDFX1 g8839(.CO(n_57), .S(n_58), .A(in_41[2]), .B(n_21), .CI(n_6));
  ADDFX1 g8840(.CO(n_55), .S(n_56), .A(in_70[1]), .B(in_80[1]), .CI(in_81[1]));
  ADDFX1 g8841(.CO(n_53), .S(n_54), .A(n_23), .B(n_4), .CI(in_62[1]));
  ADDFX1 g8842(.CO(n_51), .S(n_52), .A(in_49[1]), .B(in_78[1]), .CI(in_86[1]));
  ADDFX1 g8843(.CO(n_49), .S(n_50), .A(in_54[1]), .B(n_22), .CI(in_77[0]));
  ADDFX1 g8844(.CO(n_47), .S(n_48), .A(in_21[0]), .B(in_36[0]), .CI(n_15));
  ADDFX1 g8845(.CO(n_45), .S(n_46), .A(in_0[0]), .B(in_12[0]), .CI(in_32[0]));
  ADDFX1 g8846(.CO(n_43), .S(n_44), .A(in_14[1]), .B(in_15[1]), .CI(n_24));
  ADDFX1 g8847(.CO(n_41), .S(n_42), .A(in_22[1]), .B(in_18[0]), .CI(in_53[1]));
  ADDFX1 g8848(.CO(n_39), .S(n_40), .A(in_7[1]), .B(in_21[1]), .CI(in_10[1]));
  XNOR2X1 g8849(.Y(n_38), .A(n_34), .B(n_36));
  MX2XL g8850(.Y(n_37), .A(n_0), .B(in_2[5]), .S0(n_34));
  AOI22X1 g8851(.Y(n_36), .A0(in_3[6]), .A1(n_32), .B0(in_2[6]), .B1(in_2[5]));
  OAI21X1 g8852(.Y(n_35), .A0(in_65[0]), .A1(in_38[0]), .B0(n_31));
  XNOR2X1 g8853(.Y(n_34), .A(in_2[6]), .B(in_3[6]));
  XOR2XL g8854(.Y(n_33), .A(in_46[0]), .B(in_45[0]));
  OR2XL g8855(.Y(n_32), .A(in_2[6]), .B(in_2[5]));
  NAND2X1 g8856(.Y(n_31), .A(in_65[0]), .B(in_38[0]));
  NOR2X1 g8857(.Y(n_30), .A(in_46[0]), .B(in_45[0]));
  INVX1 g8858(.Y(n_29), .A(in_71[1]));
  INVX1 g8859(.Y(n_28), .A(in_67[0]));
  INVX1 g8860(.Y(n_27), .A(in_63[0]));
  INVX1 g8861(.Y(n_26), .A(in_25[0]));
  INVX1 g8862(.Y(n_25), .A(in_60[1]));
  INVX1 g8863(.Y(n_24), .A(in_29[1]));
  INVX1 g8864(.Y(n_23), .A(in_31[1]));
  INVX1 g8865(.Y(n_22), .A(in_33[1]));
  INVX1 g8866(.Y(n_21), .A(in_15[2]));
  INVX1 g8867(.Y(n_20), .A(in_10[2]));
  INVX1 g8868(.Y(n_19), .A(in_37[0]));
  INVX1 g8869(.Y(n_18), .A(in_64[1]));
  INVX1 g8870(.Y(n_17), .A(in_13[1]));
  INVX1 g8871(.Y(n_16), .A(in_68[0]));
  INVX1 g8872(.Y(n_15), .A(in_85[0]));
  INVX1 g8873(.Y(n_14), .A(in_50[0]));
  INVX1 g8874(.Y(n_13), .A(in_6[0]));
  INVX1 g8875(.Y(n_12), .A(in_30[0]));
  INVX1 g8876(.Y(n_11), .A(in_16[0]));
  INVX1 g8877(.Y(n_10), .A(in_35[1]));
  INVX1 g8878(.Y(n_9), .A(in_27[1]));
  INVX1 g8879(.Y(n_8), .A(in_44[0]));
  INVX1 g8880(.Y(n_7), .A(in_11[0]));
  INVX1 g8881(.Y(n_6), .A(in_7[2]));
  INVX1 g8882(.Y(n_5), .A(in_39[0]));
  INVX1 g8883(.Y(n_4), .A(in_57[1]));
  INVX1 g8884(.Y(n_3), .A(in_21[2]));
  INVX1 g8885(.Y(n_2), .A(in_52[1]));
  INVX1 g8886(.Y(n_1), .A(in_1[0]));
  INVX1 g8887(.Y(n_0), .A(in_2[5]));
endmodule

module WALLACE_CSA_DUMMY_OP8_group_359302(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, out_0);
input  in_11, in_12, in_15, in_17, in_21, in_25;
input   [4:0] in_0;
input   [5:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [4:0] in_4;
input   [2:0] in_5;
input   [4:0] in_6;
input   [2:0] in_7;
input   [4:0] in_8;
input   [1:0] in_9;
input   [1:0] in_10;
input   [1:0] in_13;
input   [1:0] in_14;
input   [2:0] in_16;
input   [1:0] in_18;
input   [2:0] in_19;
input   [1:0] in_20;
input   [2:0] in_22;
input   [4:0] in_23;
input   [1:0] in_24;
output  [9:0] out_0;
wire  n_59, n_56, n_54, n_53, n_52, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_43, n_42, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1, in_25, in_21, in_17, in_15, in_12, in_11;
wire   [9:0] out_0;
wire   [1:0] in_24;
wire   [1:0] in_20;
wire   [1:0] in_18;
wire   [1:0] in_14;
wire   [1:0] in_13;
wire   [1:0] in_10;
wire   [1:0] in_9;
wire   [2:0] in_22;
wire   [2:0] in_19;
wire   [2:0] in_16;
wire   [2:0] in_7;
wire   [2:0] in_5;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [5:0] in_1;
wire   [4:0] in_23;
wire   [4:0] in_8;
wire   [4:0] in_6;
wire   [4:0] in_4;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  AO21XL g1873(.Y(out_0[5]), .A0(n_29), .A1(n_59), .B0(out_0[9]));
  NOR2X1 g1874(.Y(out_0[9]), .A(n_29), .B(n_59));
  ADDFX1 g1875(.CO(n_59), .S(out_0[4]), .A(n_28), .B(n_48), .CI(n_56));
  ADDFX1 g1876(.CO(n_56), .S(out_0[3]), .A(n_49), .B(n_52), .CI(n_54));
  ADDFX1 g1877(.CO(n_54), .S(out_0[2]), .A(n_42), .B(n_53), .CI(n_50));
  ADDFX1 g1878(.CO(n_52), .S(n_53), .A(n_39), .B(n_47), .CI(n_44));
  ADDFX1 g1879(.CO(n_50), .S(out_0[1]), .A(n_40), .B(n_45), .CI(n_43));
  ADDFX1 g1880(.CO(n_48), .S(n_49), .A(n_28), .B(n_38), .CI(n_46));
  ADDFX1 g1881(.CO(n_46), .S(n_47), .A(n_36), .B(n_30), .CI(n_32));
  ADDFX1 g1882(.CO(n_44), .S(n_45), .A(n_16), .B(n_37), .CI(n_31));
  ADDFX1 g1883(.CO(n_42), .S(n_43), .A(n_25), .B(n_34), .CI(n_33));
  ADDFX1 g1884(.CO(n_40), .S(out_0[0]), .A(n_14), .B(n_26), .CI(n_35));
  ADDFX1 g1885(.CO(n_38), .S(n_39), .A(n_21), .B(n_15), .CI(n_27));
  ADDFX1 g1886(.CO(n_36), .S(n_37), .A(in_2[1]), .B(n_19), .CI(n_17));
  ADDFX1 g1887(.CO(n_34), .S(n_35), .A(n_18), .B(n_24), .CI(n_20));
  ADDFX1 g1888(.CO(n_32), .S(n_33), .A(n_12), .B(n_10), .CI(n_22));
  ADDFX1 g1889(.CO(n_30), .S(n_31), .A(n_7), .B(n_23), .CI(n_13));
  INVX1 g1890(.Y(n_28), .A(n_29));
  ADDHX1 g1891(.CO(n_29), .S(n_27), .A(n_11), .B(n_9));
  ADDFX1 g1892(.CO(n_25), .S(n_26), .A(in_11), .B(in_19[0]), .CI(n_8));
  ADDFX1 g1893(.CO(n_23), .S(n_24), .A(in_15), .B(in_25), .CI(n_3));
  ADDFX1 g1894(.CO(n_21), .S(n_22), .A(in_20[1]), .B(in_18[1]), .CI(in_24[1]));
  ADDFX1 g1895(.CO(n_19), .S(n_20), .A(in_9[0]), .B(in_21), .CI(n_6));
  ADDFX1 g1896(.CO(n_17), .S(n_18), .A(in_17), .B(in_7[0]), .CI(n_5));
  ADDFX1 g1897(.CO(n_15), .S(n_16), .A(in_10[0]), .B(in_13[1]), .CI(in_16[1]));
  ADDFX1 g1898(.CO(n_13), .S(n_14), .A(in_3[0]), .B(n_2), .CI(in_12));
  ADDFX1 g1899(.CO(n_11), .S(n_12), .A(in_14[1]), .B(in_19[0]), .CI(in_22[1]));
  ADDFX1 g1900(.CO(n_9), .S(n_10), .A(in_5[1]), .B(n_4), .CI(in_7[0]));
  OAI21X1 g1901(.Y(n_8), .A0(in_0[0]), .A1(n_1), .B0(n_7));
  NAND2X1 g1902(.Y(n_7), .A(in_0[0]), .B(n_1));
  INVX1 g1903(.Y(n_6), .A(in_8[0]));
  INVX1 g1904(.Y(n_5), .A(in_23[0]));
  INVX1 g1905(.Y(n_4), .A(in_1[1]));
  INVX1 g1906(.Y(n_3), .A(in_4[0]));
  INVX1 g1907(.Y(n_2), .A(in_6[0]));
  INVX1 g1908(.Y(n_1), .A(in_10[0]));
endmodule

module WALLACE_CSA_DUMMY_OP12_group_106221(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88, in_89, in_90
    , in_91, in_92, in_93, in_94, in_95, in_96, in_97, in_98, in_99, in_100, 
    in_101, in_102, in_103, out_0);
input  in_42, in_66, in_69, in_72, in_82, in_83, in_92, in_102, in_103;
input   [4:0] in_0;
input   [9:0] in_1;
input   [8:0] in_2;
input   [8:0] in_3;
input   [8:0] in_4;
input   [7:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [1:0] in_39;
input   [2:0] in_40;
input   [4:0] in_41;
input   [1:0] in_43;
input   [1:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [1:0] in_48;
input   [4:0] in_49;
input   [1:0] in_50;
input   [4:0] in_51;
input   [1:0] in_52;
input   [1:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [1:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [4:0] in_62;
input   [4:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [1:0] in_67;
input   [1:0] in_68;
input   [4:0] in_70;
input   [1:0] in_71;
input   [1:0] in_73;
input   [4:0] in_74;
input   [4:0] in_75;
input   [4:0] in_76;
input   [1:0] in_77;
input   [2:0] in_78;
input   [4:0] in_79;
input   [4:0] in_80;
input   [1:0] in_81;
input   [4:0] in_84;
input   [4:0] in_85;
input   [1:0] in_86;
input   [4:0] in_87;
input   [1:0] in_88;
input   [4:0] in_89;
input   [4:0] in_90;
input   [4:0] in_91;
input   [1:0] in_93;
input   [1:0] in_94;
input   [4:0] in_95;
input   [2:0] in_96;
input   [1:0] in_97;
input   [1:0] in_98;
input   [4:0] in_99;
input   [2:0] in_100;
input   [1:0] in_101;
output  [9:0] out_0;
wire  n_333, n_331, n_329, n_327, n_325, n_324, n_323, n_322, n_321, n_320, 
    n_319, n_318, n_317, n_315, n_314, n_313, n_312, n_311, n_310, n_309, 
    n_308, n_307, n_305, n_304, n_303, n_302, n_301, n_300, n_299, n_298, 
    n_297, n_296, n_295, n_294, n_293, n_292, n_291, n_290, n_289, n_288, 
    n_287, n_286, n_285, n_284, n_283, n_282, n_281, n_280, n_279, n_278, 
    n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, n_268, 
    n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
    n_257, n_256, n_255, n_254, n_253, n_251, n_250, n_249, n_248, n_247, 
    n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, n_237, 
    n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, n_227, 
    n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, n_218, n_217, 
    n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, n_207, 
    n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
    n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, n_187, 
    n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, 
    n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
    n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, 
    n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, 
    n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
    n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, 
    n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_103, 
    in_102, in_92, in_83, in_82, in_72, in_69, in_66, in_42;
wire   [9:0] out_0;
wire   [1:0] in_101;
wire   [1:0] in_98;
wire   [1:0] in_97;
wire   [1:0] in_94;
wire   [1:0] in_93;
wire   [1:0] in_88;
wire   [1:0] in_86;
wire   [1:0] in_81;
wire   [1:0] in_77;
wire   [1:0] in_73;
wire   [1:0] in_71;
wire   [1:0] in_68;
wire   [1:0] in_67;
wire   [1:0] in_61;
wire   [1:0] in_56;
wire   [1:0] in_53;
wire   [1:0] in_52;
wire   [1:0] in_50;
wire   [1:0] in_48;
wire   [1:0] in_44;
wire   [1:0] in_43;
wire   [1:0] in_39;
wire   [2:0] in_100;
wire   [2:0] in_96;
wire   [2:0] in_78;
wire   [2:0] in_40;
wire   [2:0] in_34;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [7:0] in_5;
wire   [8:0] in_4;
wire   [8:0] in_3;
wire   [8:0] in_2;
wire   [9:0] in_1;
wire   [4:0] in_99;
wire   [4:0] in_95;
wire   [4:0] in_91;
wire   [4:0] in_90;
wire   [4:0] in_89;
wire   [4:0] in_87;
wire   [4:0] in_85;
wire   [4:0] in_84;
wire   [4:0] in_80;
wire   [4:0] in_79;
wire   [4:0] in_76;
wire   [4:0] in_75;
wire   [4:0] in_74;
wire   [4:0] in_70;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_63;
wire   [4:0] in_62;
wire   [4:0] in_60;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_51;
wire   [4:0] in_49;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_41;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g10428(.Y(out_0[9]), .A(n_333));
  ADDFX1 g10429(.CO(n_333), .S(out_0[7]), .A(n_295), .B(n_319), .CI(n_331));
  ADDFX1 g10430(.CO(n_331), .S(out_0[6]), .A(n_320), .B(n_323), .CI(n_329));
  ADDFX1 g10431(.CO(n_329), .S(out_0[5]), .A(n_321), .B(n_327), .CI(n_324));
  ADDFX1 g10432(.CO(n_327), .S(out_0[4]), .A(n_317), .B(n_322), .CI(n_325));
  ADDFX1 g10433(.CO(n_325), .S(out_0[3]), .A(n_308), .B(n_318), .CI(n_315));
  ADDFX1 g10434(.CO(n_323), .S(n_324), .A(n_303), .B(n_311), .CI(n_314));
  ADDFX1 g10435(.CO(n_321), .S(n_322), .A(n_304), .B(n_307), .CI(n_312));
  ADDFX1 g10436(.CO(n_319), .S(n_320), .A(n_296), .B(n_299), .CI(n_313));
  ADDFX1 g10437(.CO(n_317), .S(n_318), .A(n_293), .B(n_302), .CI(n_309));
  ADDFX1 g10438(.CO(n_315), .S(out_0[2]), .A(n_294), .B(n_305), .CI(n_310));
  ADDFX1 g10439(.CO(n_313), .S(n_314), .A(n_297), .B(n_291), .CI(n_300));
  ADDFX1 g10440(.CO(n_311), .S(n_312), .A(n_301), .B(n_298), .CI(n_285));
  ADDFX1 g10441(.CO(n_309), .S(n_310), .A(n_288), .B(n_281), .CI(n_284));
  ADDFX1 g10442(.CO(n_307), .S(n_308), .A(n_290), .B(n_283), .CI(n_286));
  ADDFX1 g10443(.CO(n_305), .S(out_0[1]), .A(n_251), .B(n_244), .CI(n_282));
  ADDFX1 g10444(.CO(n_303), .S(n_304), .A(n_289), .B(n_292), .CI(n_278));
  ADDFX1 g10445(.CO(n_301), .S(n_302), .A(n_280), .B(n_287), .CI(n_273));
  ADDFX1 g10446(.CO(n_299), .S(n_300), .A(n_194), .B(n_277), .CI(n_276));
  ADDFX1 g10447(.CO(n_297), .S(n_298), .A(n_279), .B(n_258), .CI(n_269));
  ADDFX1 g10448(.CO(n_295), .S(n_296), .A(n_193), .B(n_34), .CI(n_275));
  ADDFX1 g10449(.CO(n_293), .S(n_294), .A(n_243), .B(n_246), .CI(n_274));
  ADDFX1 g10450(.CO(n_291), .S(n_292), .A(n_253), .B(n_247), .CI(n_271));
  ADDFX1 g10451(.CO(n_289), .S(n_290), .A(n_248), .B(n_245), .CI(n_267));
  ADDFX1 g10452(.CO(n_287), .S(n_288), .A(n_262), .B(n_265), .CI(n_250));
  ADDFX1 g10453(.CO(n_285), .S(n_286), .A(n_263), .B(n_270), .CI(n_272));
  ADDFX1 g10454(.CO(n_283), .S(n_284), .A(n_264), .B(n_255), .CI(n_268));
  ADDFX1 g10455(.CO(n_281), .S(n_282), .A(n_266), .B(n_260), .CI(n_256));
  ADDFX1 g10456(.CO(n_279), .S(n_280), .A(n_261), .B(n_254), .CI(n_249));
  ADDFX1 g10457(.CO(n_277), .S(n_278), .A(n_242), .B(n_239), .CI(in_1[4]));
  ADDFX1 g10458(.CO(n_275), .S(n_276), .A(n_241), .B(n_257), .CI(in_1[5]));
  ADDFX1 g10459(.CO(n_273), .S(n_274), .A(n_197), .B(n_259), .CI(n_225));
  ADDFX1 g10460(.CO(n_271), .S(n_272), .A(n_233), .B(n_232), .CI(in_1[3]));
  ADDFX1 g10461(.CO(n_269), .S(n_270), .A(n_229), .B(n_222), .CI(n_240));
  ADDFX1 g10462(.CO(n_267), .S(n_268), .A(n_237), .B(n_202), .CI(in_1[2]));
  ADDFX1 g10463(.CO(n_265), .S(n_266), .A(n_238), .B(n_191), .CI(n_208));
  ADDFX1 g10464(.CO(n_263), .S(n_264), .A(n_236), .B(n_234), .CI(n_230));
  ADDFX1 g10465(.CO(n_261), .S(n_262), .A(n_220), .B(n_215), .CI(n_207));
  ADDFX1 g10466(.CO(n_259), .S(n_260), .A(n_216), .B(n_223), .CI(n_210));
  ADDFX1 g10467(.CO(n_257), .S(n_258), .A(n_192), .B(n_213), .CI(n_221));
  ADDFX1 g10468(.CO(n_255), .S(n_256), .A(n_212), .B(n_203), .CI(n_226));
  ADDFX1 g10469(.CO(n_253), .S(n_254), .A(n_227), .B(n_201), .CI(n_214));
  ADDFX1 g10470(.CO(n_251), .S(out_0[0]), .A(n_204), .B(n_224), .CI(n_200));
  ADDFX1 g10471(.CO(n_249), .S(n_250), .A(n_228), .B(n_211), .CI(n_209));
  ADDFX1 g10472(.CO(n_247), .S(n_248), .A(n_235), .B(n_217), .CI(n_195));
  ADDFX1 g10473(.CO(n_245), .S(n_246), .A(n_205), .B(n_218), .CI(n_196));
  ADDFX1 g10474(.CO(n_243), .S(n_244), .A(n_206), .B(n_198), .CI(n_199));
  ADDFX1 g10475(.CO(n_241), .S(n_242), .A(n_231), .B(n_25), .CI(n_26));
  ADDFX1 g10476(.CO(n_239), .S(n_240), .A(n_173), .B(n_219), .CI(in_4[3]));
  ADDFX1 g10477(.CO(n_237), .S(n_238), .A(n_177), .B(n_188), .CI(n_140));
  ADDFX1 g10478(.CO(n_235), .S(n_236), .A(n_165), .B(n_137), .CI(n_163));
  ADDFX1 g10479(.CO(n_233), .S(n_234), .A(n_180), .B(n_185), .CI(n_146));
  ADDFX1 g10480(.CO(n_231), .S(n_232), .A(n_132), .B(n_164), .CI(n_7));
  ADDFX1 g10481(.CO(n_229), .S(n_230), .A(n_186), .B(n_159), .CI(n_190));
  ADDFX1 g10482(.CO(n_227), .S(n_228), .A(n_166), .B(n_160), .CI(n_133));
  ADDFX1 g10483(.CO(n_225), .S(n_226), .A(n_187), .B(n_153), .CI(in_1[1]));
  ADDFX1 g10484(.CO(n_223), .S(n_224), .A(n_175), .B(n_189), .CI(n_141));
  ADDFX1 g10485(.CO(n_221), .S(n_222), .A(n_162), .B(n_158), .CI(in_3[3]));
  ADDFX1 g10486(.CO(n_219), .S(n_220), .A(n_148), .B(n_134), .CI(n_176));
  ADDFX1 g10487(.CO(n_217), .S(n_218), .A(n_150), .B(n_182), .CI(in_2[2]));
  ADDFX1 g10488(.CO(n_215), .S(n_216), .A(n_161), .B(n_139), .CI(n_168));
  ADDFX1 g10489(.CO(n_213), .S(n_214), .A(n_136), .B(n_184), .CI(in_2[3]));
  ADDFX1 g10490(.CO(n_211), .S(n_212), .A(n_167), .B(n_157), .CI(n_144));
  ADDFX1 g10491(.CO(n_209), .S(n_210), .A(n_170), .B(n_154), .CI(in_3[1]));
  ADDFX1 g10492(.CO(n_207), .S(n_208), .A(n_149), .B(n_174), .CI(in_2[1]));
  ADDFX1 g10493(.CO(n_205), .S(n_206), .A(n_181), .B(n_151), .CI(n_183));
  ADDFX1 g10494(.CO(n_203), .S(n_204), .A(n_155), .B(n_169), .CI(n_145));
  ADDFX1 g10495(.CO(n_201), .S(n_202), .A(n_138), .B(n_156), .CI(in_5[2]));
  ADDFX1 g10496(.CO(n_199), .S(n_200), .A(n_171), .B(n_143), .CI(n_179));
  ADDFX1 g10497(.CO(n_197), .S(n_198), .A(n_147), .B(n_142), .CI(n_178));
  ADDFX1 g10498(.CO(n_195), .S(n_196), .A(n_152), .B(in_3[2]), .CI(in_4[2]));
  INVX1 g10499(.Y(n_194), .A(n_193));
  ADDFX1 g10500(.CO(n_193), .S(n_192), .A(n_0), .B(n_172), .CI(n_36));
  ADDFX1 g10501(.CO(n_190), .S(n_191), .A(n_66), .B(n_135), .CI(in_4[1]));
  ADDFX1 g10502(.CO(n_188), .S(n_189), .A(n_119), .B(n_65), .CI(n_127));
  ADDFX1 g10503(.CO(n_186), .S(n_187), .A(n_113), .B(n_125), .CI(n_123));
  ADDFX1 g10504(.CO(n_184), .S(n_185), .A(n_124), .B(n_80), .CI(n_114));
  ADDFX1 g10505(.CO(n_182), .S(n_183), .A(n_75), .B(n_97), .CI(in_5[1]));
  ADDFX1 g10506(.CO(n_180), .S(n_181), .A(n_72), .B(n_103), .CI(n_115));
  ADDFX1 g10507(.CO(n_178), .S(n_179), .A(n_57), .B(n_129), .CI(in_1[0]));
  ADDFX1 g10508(.CO(n_176), .S(n_177), .A(n_68), .B(n_126), .CI(n_108));
  ADDFX1 g10509(.CO(n_174), .S(n_175), .A(n_85), .B(n_109), .CI(n_101));
  ADDFX1 g10510(.CO(n_172), .S(n_173), .A(in_65[0]), .B(n_110), .CI(n_60));
  ADDFX1 g10511(.CO(n_170), .S(n_171), .A(n_73), .B(n_89), .CI(n_117));
  ADDFX1 g10512(.CO(n_168), .S(n_169), .A(n_63), .B(n_105), .CI(n_69));
  ADDFX1 g10513(.CO(n_166), .S(n_167), .A(n_88), .B(n_100), .CI(n_104));
  ADDFX1 g10514(.CO(n_164), .S(n_165), .A(n_50), .B(n_96), .CI(n_112));
  ADDFX1 g10515(.CO(n_162), .S(n_163), .A(n_76), .B(n_106), .CI(n_86));
  ADDFX1 g10516(.CO(n_160), .S(n_161), .A(n_98), .B(n_118), .CI(n_116));
  ADDFX1 g10517(.CO(n_158), .S(n_159), .A(n_111), .B(n_61), .CI(n_122));
  ADDFX1 g10518(.CO(n_156), .S(n_157), .A(n_70), .B(n_54), .CI(n_64));
  ADDFX1 g10519(.CO(n_154), .S(n_155), .A(n_79), .B(n_131), .CI(n_99));
  ADDFX1 g10520(.CO(n_152), .S(n_153), .A(n_59), .B(n_81), .CI(n_52));
  ADDFX1 g10521(.CO(n_150), .S(n_151), .A(n_107), .B(n_91), .CI(n_77));
  ADDFX1 g10522(.CO(n_148), .S(n_149), .A(n_78), .B(n_94), .CI(n_130));
  ADDFX1 g10523(.CO(n_146), .S(n_147), .A(n_56), .B(n_128), .CI(n_87));
  ADDFX1 g10524(.CO(n_144), .S(n_145), .A(n_55), .B(n_83), .CI(in_2[0]));
  ADDFX1 g10525(.CO(n_142), .S(n_143), .A(n_95), .B(n_67), .CI(in_3[0]));
  ADDFX1 g10526(.CO(n_140), .S(n_141), .A(n_71), .B(n_53), .CI(in_4[0]));
  ADDFX1 g10527(.CO(n_138), .S(n_139), .A(n_51), .B(n_62), .CI(n_82));
  ADDFX1 g10528(.CO(n_136), .S(n_137), .A(n_102), .B(n_90), .CI(n_74));
  ADDFX1 g10529(.CO(n_134), .S(n_135), .A(in_6[1]), .B(in_25[1]), .CI(n_84));
  ADDFX1 g10530(.CO(n_132), .S(n_133), .A(in_65[0]), .B(n_28), .CI(n_58));
  ADDFX1 g10531(.CO(n_130), .S(n_131), .A(in_39[0]), .B(n_20), .CI(n_9));
  ADDFX1 g10532(.CO(n_128), .S(n_129), .A(in_19[0]), .B(in_17[0]), .CI(in_14[0]));
  ADDFX1 g10533(.CO(n_126), .S(n_127), .A(in_21[0]), .B(in_31[0]), .CI(n_41));
  ADDFX1 g10534(.CO(n_124), .S(n_125), .A(in_97[1]), .B(n_29), .CI(in_98[1]));
  INVX1 g10535(.Y(n_123), .A(n_121));
  INVX1 g10536(.Y(n_122), .A(n_120));
  ADDFX1 g10537(.CO(n_120), .S(n_121), .A(in_28[1]), .B(in_20[1]), .CI(in_23[1]));
  ADDFX1 g10538(.CO(n_118), .S(n_119), .A(in_25[0]), .B(in_42), .CI(in_83));
  ADDFX1 g10539(.CO(n_116), .S(n_117), .A(in_56[0]), .B(n_12), .CI(in_90[0]));
  ADDFX1 g10540(.CO(n_114), .S(n_115), .A(in_40[1]), .B(in_67[0]), .CI(in_101[0]));
  ADDFX1 g10541(.CO(n_112), .S(n_113), .A(in_24[1]), .B(in_7[1]), .CI(in_78[1]));
  INVX1 g10542(.Y(n_111), .A(n_93));
  INVX1 g10543(.Y(n_110), .A(n_92));
  ADDFX1 g10544(.CO(n_108), .S(n_109), .A(in_38[0]), .B(in_50[0]), .CI(in_67[0]));
  ADDFX1 g10545(.CO(n_106), .S(n_107), .A(in_29[1]), .B(n_10), .CI(n_21));
  ADDFX1 g10546(.CO(n_104), .S(n_105), .A(in_66), .B(in_88[0]), .CI(in_101[0]));
  ADDFX1 g10547(.CO(n_102), .S(n_103), .A(n_15), .B(n_18), .CI(in_93[1]));
  ADDFX1 g10548(.CO(n_100), .S(n_101), .A(in_62[0]), .B(n_39), .CI(in_94[0]));
  ADDFX1 g10549(.CO(n_98), .S(n_99), .A(in_18[0]), .B(n_14), .CI(in_82));
  ADDFX1 g10550(.CO(n_96), .S(n_97), .A(in_15[1]), .B(n_38), .CI(n_42));
  ADDFX1 g10551(.CO(n_94), .S(n_95), .A(in_44[0]), .B(in_74[0]), .CI(n_19));
  ADDFX1 g10552(.CO(n_92), .S(n_93), .A(in_38[0]), .B(in_74[0]), .CI(in_90[0]));
  ADDFX1 g10553(.CO(n_90), .S(n_91), .A(in_96[1]), .B(n_40), .CI(n_22));
  ADDFX1 g10554(.CO(n_88), .S(n_89), .A(in_9[0]), .B(in_48[0]), .CI(n_35));
  ADDFX1 g10555(.CO(n_86), .S(n_87), .A(in_17[1]), .B(n_44), .CI(n_30));
  ADDFX1 g10556(.CO(n_84), .S(n_85), .A(n_8), .B(in_65[0]), .CI(in_72));
  ADDFX1 g10557(.CO(n_82), .S(n_83), .A(in_61[0]), .B(in_69), .CI(n_11));
  ADDFX1 g10558(.CO(n_80), .S(n_81), .A(in_68[1]), .B(n_6), .CI(n_43));
  ADDFX1 g10559(.CO(n_78), .S(n_79), .A(in_77[0]), .B(in_103), .CI(n_3));
  ADDFX1 g10560(.CO(n_76), .S(n_77), .A(n_13), .B(n_16), .CI(in_53[1]));
  ADDFX1 g10561(.CO(n_74), .S(n_75), .A(in_52[0]), .B(in_43[1]), .CI(n_23));
  ADDFX1 g10562(.CO(n_72), .S(n_73), .A(in_7[0]), .B(n_32), .CI(in_81[0]));
  ADDFX1 g10563(.CO(n_70), .S(n_71), .A(in_10[0]), .B(in_30[0]), .CI(n_31));
  ADDFX1 g10564(.CO(n_68), .S(n_69), .A(in_71[0]), .B(in_11[0]), .CI(in_102));
  ADDFX1 g10565(.CO(n_66), .S(n_67), .A(in_6[0]), .B(in_28[0]), .CI(in_5[0]));
  ADDFX1 g10566(.CO(n_64), .S(n_65), .A(in_52[0]), .B(n_27), .CI(in_92));
  ADDFX1 g10567(.CO(n_62), .S(n_63), .A(in_86[0]), .B(n_5), .CI(n_45));
  ADDFX1 g10568(.CO(n_60), .S(n_61), .A(n_1), .B(in_100[2]), .CI(n_33));
  ADDFX1 g10569(.CO(n_58), .S(n_59), .A(n_37), .B(in_34[1]), .CI(n_24));
  ADDFX1 g10570(.CO(n_56), .S(n_57), .A(n_17), .B(in_20[0]), .CI(in_23[0]));
  ADDFX1 g10571(.CO(n_54), .S(n_55), .A(in_33[0]), .B(n_4), .CI(n_46));
  XOR2XL g10572(.Y(n_53), .A(in_60[0]), .B(n_47));
  XOR2XL g10573(.Y(n_52), .A(in_26[1]), .B(n_47));
  OAI21X1 g10574(.Y(n_51), .A0(in_60[0]), .A1(n_2), .B0(n_48));
  OAI21X1 g10575(.Y(n_50), .A0(in_26[1]), .A1(n_2), .B0(n_49));
  OAI2BB1X1 g10576(.Y(n_49), .A0N(in_26[1]), .A1N(n_2), .B0(in_73[0]));
  OAI2BB1X1 g10577(.Y(n_48), .A0N(in_60[0]), .A1N(n_2), .B0(in_73[0]));
  MXI2XL g10578(.Y(n_47), .A(in_12[0]), .B(n_2), .S0(in_73[0]));
  INVX1 g10579(.Y(n_46), .A(in_89[0]));
  INVX1 g10580(.Y(n_45), .A(in_87[0]));
  INVX1 g10581(.Y(n_44), .A(in_19[1]));
  INVX1 g10582(.Y(n_43), .A(in_70[1]));
  INVX1 g10583(.Y(n_42), .A(in_85[1]));
  INVX1 g10584(.Y(n_41), .A(in_51[0]));
  INVX1 g10585(.Y(n_40), .A(in_37[1]));
  INVX1 g10586(.Y(n_39), .A(in_63[0]));
  INVX1 g10587(.Y(n_38), .A(in_75[1]));
  INVX1 g10588(.Y(n_37), .A(in_35[1]));
  INVX1 g10589(.Y(n_36), .A(in_2[4]));
  INVX1 g10590(.Y(n_35), .A(in_13[0]));
  INVX1 g10591(.Y(n_34), .A(in_1[6]));
  INVX1 g10592(.Y(n_33), .A(in_6[2]));
  INVX1 g10593(.Y(n_32), .A(in_49[0]));
  INVX1 g10594(.Y(n_31), .A(in_16[0]));
  INVX1 g10595(.Y(n_30), .A(in_14[1]));
  INVX1 g10596(.Y(n_29), .A(in_36[1]));
  INVX1 g10597(.Y(n_28), .A(in_25[2]));
  INVX1 g10598(.Y(n_27), .A(in_45[0]));
  INVX1 g10599(.Y(n_26), .A(in_4[4]));
  INVX1 g10600(.Y(n_25), .A(in_3[4]));
  INVX1 g10601(.Y(n_24), .A(in_84[1]));
  INVX1 g10602(.Y(n_23), .A(in_64[1]));
  INVX1 g10603(.Y(n_22), .A(in_99[1]));
  INVX1 g10604(.Y(n_21), .A(in_95[1]));
  INVX1 g10605(.Y(n_20), .A(in_76[0]));
  INVX1 g10606(.Y(n_19), .A(in_0[0]));
  INVX1 g10607(.Y(n_18), .A(in_58[1]));
  INVX1 g10608(.Y(n_17), .A(in_8[0]));
  INVX1 g10609(.Y(n_16), .A(in_46[1]));
  INVX1 g10610(.Y(n_15), .A(in_27[1]));
  INVX1 g10611(.Y(n_14), .A(in_32[0]));
  INVX1 g10612(.Y(n_13), .A(in_41[1]));
  INVX1 g10613(.Y(n_12), .A(in_79[0]));
  INVX1 g10614(.Y(n_11), .A(in_59[0]));
  INVX1 g10615(.Y(n_10), .A(in_55[1]));
  INVX1 g10616(.Y(n_9), .A(in_47[0]));
  INVX1 g10617(.Y(n_8), .A(in_22[0]));
  INVX1 g10618(.Y(n_7), .A(in_5[3]));
  INVX1 g10619(.Y(n_6), .A(in_57[1]));
  INVX1 g10620(.Y(n_5), .A(in_54[0]));
  INVX1 g10621(.Y(n_4), .A(in_80[0]));
  INVX1 g10622(.Y(n_3), .A(in_91[0]));
  INVX1 g10623(.Y(n_2), .A(in_12[0]));
  INVX1 g10624(.Y(n_1), .A(in_62[0]));
  INVX1 g10625(.Y(n_0), .A(in_65[0]));
endmodule

module WALLACE_CSA_DUMMY_OP17_group_106212(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, out_0);
input  in_28, in_29;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [9:0] in_3;
input   [9:0] in_4;
input   [9:0] in_5;
input   [6:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [4:0] in_25;
input   [2:0] in_26;
input   [1:0] in_27;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [1:0] in_42;
input   [1:0] in_43;
input   [4:0] in_44;
input   [4:0] in_45;
input   [2:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [1:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [1:0] in_59;
input   [4:0] in_60;
input   [4:0] in_61;
input   [2:0] in_62;
input   [2:0] in_63;
input   [4:0] in_64;
output  [9:0] out_0;
wire  n_225, n_223, n_221, n_219, n_217, n_216, n_215, n_214, n_213, n_211, 
    n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, 
    n_200, n_199, n_198, n_197, n_195, n_194, n_193, n_192, n_191, n_190, 
    n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, 
    n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, 
    n_169, n_168, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, 
    n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, 
    n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, 
    in_29, in_28;
wire   [9:0] out_0;
wire   [1:0] in_59;
wire   [1:0] in_51;
wire   [1:0] in_50;
wire   [1:0] in_43;
wire   [1:0] in_42;
wire   [1:0] in_34;
wire   [1:0] in_33;
wire   [1:0] in_27;
wire   [2:0] in_63;
wire   [2:0] in_62;
wire   [2:0] in_46;
wire   [2:0] in_26;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [6:0] in_6;
wire   [9:0] in_5;
wire   [9:0] in_4;
wire   [9:0] in_3;
wire   [4:0] in_64;
wire   [4:0] in_61;
wire   [4:0] in_60;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_25;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVXL g7078(.Y(out_0[9]), .A(n_225));
  ADDFX1 g7079(.CO(n_225), .S(out_0[7]), .A(n_168), .B(n_209), .CI(n_223));
  ADDFX1 g7080(.CO(n_223), .S(out_0[6]), .A(n_215), .B(n_210), .CI(n_221));
  ADDFX1 g7081(.CO(n_221), .S(out_0[5]), .A(n_213), .B(n_216), .CI(n_219));
  ADDFX1 g7082(.CO(n_219), .S(out_0[4]), .A(n_207), .B(n_214), .CI(n_217));
  ADDFX1 g7083(.CO(n_217), .S(out_0[3]), .A(n_201), .B(n_211), .CI(n_208));
  ADDFX1 g7084(.CO(n_215), .S(n_216), .A(n_165), .B(n_204), .CI(n_205));
  ADDFX1 g7085(.CO(n_213), .S(n_214), .A(n_199), .B(n_192), .CI(n_206));
  ADDFX1 g7086(.CO(n_211), .S(out_0[2]), .A(n_181), .B(n_195), .CI(n_202));
  ADDFX1 g7087(.CO(n_209), .S(n_210), .A(n_164), .B(n_203), .CI(n_156));
  ADDFX1 g7088(.CO(n_207), .S(n_208), .A(n_200), .B(n_193), .CI(n_198));
  ADDFX1 g7089(.CO(n_205), .S(n_206), .A(n_185), .B(n_197), .CI(n_190));
  ADDFX1 g7090(.CO(n_203), .S(n_204), .A(n_179), .B(n_189), .CI(n_191));
  ADDFX1 g7091(.CO(n_201), .S(n_202), .A(n_188), .B(n_172), .CI(n_194));
  ADDFX1 g7092(.CO(n_199), .S(n_200), .A(n_186), .B(n_187), .CI(n_170));
  ADDFX1 g7093(.CO(n_197), .S(n_198), .A(n_183), .B(n_176), .CI(n_171));
  ADDFX1 g7094(.CO(n_195), .S(out_0[1]), .A(n_174), .B(n_166), .CI(n_182));
  ADDFX1 g7095(.CO(n_193), .S(n_194), .A(n_160), .B(n_173), .CI(n_184));
  ADDFX1 g7096(.CO(n_191), .S(n_192), .A(n_180), .B(n_169), .CI(n_175));
  ADDFX1 g7097(.CO(n_189), .S(n_190), .A(n_177), .B(in_4[4]), .CI(in_3[4]));
  ADDFX1 g7098(.CO(n_187), .S(n_188), .A(n_159), .B(n_140), .CI(n_163));
  ADDFX1 g7099(.CO(n_185), .S(n_186), .A(n_158), .B(n_162), .CI(n_178));
  ADDFX1 g7100(.CO(n_183), .S(n_184), .A(n_150), .B(n_148), .CI(in_4[2]));
  ADDFX1 g7101(.CO(n_181), .S(n_182), .A(n_149), .B(n_161), .CI(n_131));
  ADDFX1 g7102(.CO(n_179), .S(n_180), .A(n_134), .B(n_154), .CI(n_127));
  ADDFX1 g7103(.CO(n_177), .S(n_178), .A(n_143), .B(n_141), .CI(in_5[3]));
  ADDFX1 g7104(.CO(n_175), .S(n_176), .A(n_135), .B(n_152), .CI(in_3[3]));
  ADDFX1 g7105(.CO(n_173), .S(n_174), .A(n_138), .B(n_151), .CI(n_133));
  ADDFX1 g7106(.CO(n_171), .S(n_172), .A(n_153), .B(in_3[2]), .CI(n_130));
  ADDFX1 g7107(.CO(n_169), .S(n_170), .A(n_155), .B(n_139), .CI(in_4[3]));
  XNOR2X1 g7108(.Y(n_168), .A(n_157), .B(n_88));
  ADDFX1 g7109(.CO(n_166), .S(out_0[0]), .A(n_112), .B(n_146), .CI(n_129));
  ADDFX1 g7110(.CO(n_164), .S(n_165), .A(n_147), .B(in_4[5]), .CI(in_3[5]));
  ADDFX1 g7111(.CO(n_162), .S(n_163), .A(n_144), .B(n_137), .CI(n_132));
  ADDFX1 g7112(.CO(n_160), .S(n_161), .A(n_145), .B(n_111), .CI(n_128));
  ADDFX1 g7113(.CO(n_158), .S(n_159), .A(n_117), .B(n_114), .CI(n_142));
  OAI21X1 g7114(.Y(n_157), .A0(n_136), .A1(n_27), .B0(n_28));
  XNOR2X1 g7115(.Y(n_156), .A(n_136), .B(n_29));
  ADDFX1 g7116(.CO(n_154), .S(n_155), .A(n_124), .B(n_121), .CI(n_113));
  ADDFX1 g7117(.CO(n_152), .S(n_153), .A(n_122), .B(n_125), .CI(n_105));
  ADDFX1 g7118(.CO(n_150), .S(n_151), .A(n_123), .B(n_95), .CI(n_97));
  ADDFX1 g7119(.CO(n_148), .S(n_149), .A(n_107), .B(n_106), .CI(n_118));
  AO21X1 g7120(.Y(n_147), .A0(in_5[5]), .A1(n_126), .B0(n_136));
  ADDFX1 g7121(.CO(n_145), .S(n_146), .A(n_108), .B(n_96), .CI(n_102));
  ADDFX1 g7122(.CO(n_143), .S(n_144), .A(n_92), .B(n_99), .CI(n_109));
  ADDFX1 g7123(.CO(n_141), .S(n_142), .A(n_62), .B(n_115), .CI(n_89));
  ADDFX1 g7124(.CO(n_139), .S(n_140), .A(n_94), .B(n_103), .CI(in_5[2]));
  ADDFX1 g7125(.CO(n_137), .S(n_138), .A(n_116), .B(n_110), .CI(n_101));
  NOR2X1 g7126(.Y(n_136), .A(in_5[5]), .B(n_126));
  ADDFX1 g7127(.CO(n_134), .S(n_135), .A(n_91), .B(n_61), .CI(n_93));
  ADDFX1 g7128(.CO(n_132), .S(n_133), .A(n_100), .B(n_90), .CI(in_5[1]));
  ADDFX1 g7129(.CO(n_130), .S(n_131), .A(n_104), .B(in_4[1]), .CI(in_3[1]));
  ADDFX1 g7130(.CO(n_128), .S(n_129), .A(n_98), .B(in_4[0]), .CI(in_3[0]));
  XNOR2X1 g7131(.Y(n_127), .A(n_120), .B(in_5[4]));
  NOR2BX1 g7132(.Y(n_126), .AN(in_5[4]), .B(n_120));
  ADDFX1 g7133(.CO(n_124), .S(n_125), .A(n_54), .B(n_67), .CI(n_65));
  ADDFX1 g7134(.CO(n_122), .S(n_123), .A(n_83), .B(n_38), .CI(n_64));
  INVX1 g7135(.Y(n_121), .A(n_119));
  ADDFX1 g7136(.CO(n_120), .S(n_119), .A(in_60[0]), .B(n_73), .CI(n_32));
  ADDFX1 g7137(.CO(n_117), .S(n_118), .A(n_68), .B(n_55), .CI(n_66));
  ADDFX1 g7138(.CO(n_115), .S(n_116), .A(n_22), .B(n_79), .CI(n_52));
  ADDFX1 g7139(.CO(n_113), .S(n_114), .A(n_85), .B(n_60), .CI(n_30));
  ADDFX1 g7140(.CO(n_111), .S(n_112), .A(n_76), .B(n_57), .CI(in_5[0]));
  ADDFX1 g7141(.CO(n_109), .S(n_110), .A(n_34), .B(n_77), .CI(n_71));
  ADDFX1 g7142(.CO(n_107), .S(n_108), .A(n_39), .B(n_37), .CI(n_35));
  ADDFX1 g7143(.CO(n_105), .S(n_106), .A(n_41), .B(n_47), .CI(n_70));
  ADDFX1 g7144(.CO(n_103), .S(n_104), .A(n_75), .B(n_31), .CI(n_56));
  ADDFX1 g7145(.CO(n_101), .S(n_102), .A(n_78), .B(n_80), .CI(n_87));
  ADDFX1 g7146(.CO(n_99), .S(n_100), .A(n_36), .B(n_48), .CI(n_44));
  ADDFX1 g7147(.CO(n_97), .S(n_98), .A(n_25), .B(n_49), .CI(n_84));
  ADDFX1 g7148(.CO(n_95), .S(n_96), .A(n_72), .B(n_45), .CI(n_53));
  ADDFX1 g7149(.CO(n_93), .S(n_94), .A(n_46), .B(n_69), .CI(n_63));
  ADDFX1 g7150(.CO(n_91), .S(n_92), .A(in_60[0]), .B(n_21), .CI(n_40));
  ADDFX1 g7151(.CO(n_89), .S(n_90), .A(n_24), .B(n_86), .CI(in_9[1]));
  XNOR2X1 g7152(.Y(n_88), .A(n_23), .B(n_29));
  INVX1 g7153(.Y(n_87), .A(n_82));
  INVX1 g7154(.Y(n_86), .A(n_81));
  INVX1 g7155(.Y(n_85), .A(n_74));
  ADDFX1 g7156(.CO(n_83), .S(n_84), .A(in_21[0]), .B(n_6), .CI(in_59[0]));
  ADDFX1 g7157(.CO(n_81), .S(n_82), .A(in_37[0]), .B(in_49[0]), .CI(in_2[0]));
  ADDFX1 g7158(.CO(n_79), .S(n_80), .A(in_8[0]), .B(n_15), .CI(in_33[0]));
  ADDFX1 g7159(.CO(n_77), .S(n_78), .A(in_11[0]), .B(in_50[0]), .CI(n_4));
  ADDFX1 g7160(.CO(n_75), .S(n_76), .A(in_15[0]), .B(in_13[0]), .CI(in_12[0]));
  ADDFX1 g7161(.CO(n_73), .S(n_74), .A(in_36[0]), .B(in_16[0]), .CI(in_58[0]));
  ADDFX1 g7162(.CO(n_71), .S(n_72), .A(in_7[0]), .B(n_1), .CI(in_58[0]));
  ADDFX1 g7163(.CO(n_69), .S(n_70), .A(in_19[1]), .B(n_5), .CI(n_9));
  ADDFX1 g7164(.CO(n_67), .S(n_68), .A(in_46[1]), .B(n_19), .CI(n_14));
  INVX1 g7165(.Y(n_66), .A(n_59));
  INVX1 g7166(.Y(n_65), .A(n_58));
  INVX1 g7167(.Y(n_64), .A(n_51));
  INVX1 g7168(.Y(n_63), .A(n_50));
  INVX1 g7169(.Y(n_62), .A(n_43));
  INVX1 g7170(.Y(n_61), .A(n_42));
  INVX1 g7171(.Y(n_60), .A(n_33));
  ADDFX1 g7172(.CO(n_58), .S(n_59), .A(in_15[1]), .B(in_13[1]), .CI(in_20[1]));
  ADDFX1 g7173(.CO(n_56), .S(n_57), .A(in_38[0]), .B(in_23[0]), .CI(in_20[0]));
  ADDFX1 g7174(.CO(n_54), .S(n_55), .A(in_26[1]), .B(n_13), .CI(n_11));
  ADDFX1 g7175(.CO(n_52), .S(n_53), .A(in_42[0]), .B(n_0), .CI(n_18));
  ADDFX1 g7176(.CO(n_50), .S(n_51), .A(in_39[1]), .B(in_41[1]), .CI(in_64[1]));
  ADDFX1 g7177(.CO(n_48), .S(n_49), .A(in_29), .B(n_7), .CI(in_60[0]));
  ADDFX1 g7178(.CO(n_46), .S(n_47), .A(n_17), .B(n_3), .CI(in_18[1]));
  ADDFX1 g7179(.CO(n_44), .S(n_45), .A(in_16[0]), .B(n_8), .CI(in_45[0]));
  ADDFX1 g7180(.CO(n_42), .S(n_43), .A(in_45[0]), .B(in_9[2]), .CI(in_12[2]));
  ADDFX1 g7181(.CO(n_40), .S(n_41), .A(n_16), .B(in_14[1]), .CI(in_62[1]));
  ADDFX1 g7182(.CO(n_38), .S(n_39), .A(in_36[0]), .B(in_43[0]), .CI(n_12));
  ADDFX1 g7183(.CO(n_36), .S(n_37), .A(in_9[0]), .B(in_28), .CI(n_10));
  ADDFX1 g7184(.CO(n_34), .S(n_35), .A(in_27[0]), .B(in_34[0]), .CI(in_51[0]));
  ADDFX1 g7185(.CO(n_32), .S(n_33), .A(in_11[0]), .B(in_8[0]), .CI(in_38[0]));
  ADDFX1 g7186(.CO(n_30), .S(n_31), .A(n_20), .B(n_2), .CI(in_12[1]));
  NOR2BX1 g7187(.Y(n_29), .AN(n_28), .B(n_27));
  NAND2BX1 g7188(.Y(n_28), .AN(n_26), .B(in_3[6]));
  NOR2BX1 g7189(.Y(n_27), .AN(n_26), .B(in_3[6]));
  OAI21X1 g7190(.Y(n_26), .A0(in_5[5]), .A1(in_4[6]), .B0(n_23));
  OAI21X1 g7191(.Y(n_25), .A0(in_17[0]), .A1(in_53[0]), .B0(n_22));
  XNOR2X1 g7192(.Y(n_24), .A(in_44[1]), .B(in_63[1]));
  NAND2X1 g7193(.Y(n_23), .A(in_5[5]), .B(in_4[6]));
  NAND2X1 g7194(.Y(n_22), .A(in_53[0]), .B(in_17[0]));
  NOR2BX1 g7195(.Y(n_21), .AN(in_63[1]), .B(in_44[1]));
  INVX1 g7196(.Y(n_20), .A(in_47[1]));
  INVX1 g7197(.Y(n_19), .A(in_57[1]));
  INVX1 g7198(.Y(n_18), .A(in_56[0]));
  INVX1 g7199(.Y(n_17), .A(in_1[1]));
  INVX1 g7200(.Y(n_16), .A(in_32[1]));
  INVX1 g7201(.Y(n_15), .A(in_22[0]));
  INVX1 g7202(.Y(n_14), .A(in_35[1]));
  INVX1 g7203(.Y(n_13), .A(in_55[1]));
  INVX1 g7204(.Y(n_12), .A(in_52[0]));
  INVX1 g7205(.Y(n_11), .A(in_61[1]));
  INVX1 g7206(.Y(n_10), .A(in_40[0]));
  INVX1 g7207(.Y(n_9), .A(in_48[1]));
  INVX1 g7208(.Y(n_8), .A(in_25[0]));
  INVX1 g7209(.Y(n_7), .A(in_30[0]));
  INVX1 g7210(.Y(n_6), .A(in_6[0]));
  INVX1 g7211(.Y(n_5), .A(in_31[1]));
  INVX1 g7212(.Y(n_4), .A(in_0[0]));
  INVX1 g7213(.Y(n_3), .A(in_10[1]));
  INVX1 g7214(.Y(n_2), .A(in_23[1]));
  INVX1 g7215(.Y(n_1), .A(in_24[0]));
  INVX1 g7216(.Y(n_0), .A(in_54[0]));
endmodule

module WALLACE_CSA_DUMMY_OP22_group_106194(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, out_0);
input  in_18, in_19;
input   [4:0] in_0;
input   [6:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [4:0] in_15;
input   [2:0] in_16;
input   [1:0] in_17;
input   [1:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [2:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [1:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
output  [9:0] out_0;
wire  n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
    n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, 
    n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_52, n_49, n_47, n_45, n_44, n_43, n_41, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_1, in_19, in_18;
wire   [9:0] out_0;
wire   [1:0] in_39;
wire   [1:0] in_22;
wire   [1:0] in_20;
wire   [1:0] in_17;
wire   [2:0] in_32;
wire   [2:0] in_29;
wire   [2:0] in_16;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [6:0] in_1;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_15;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_134), .S(n_133), .A(n_26), .B(n_10), .CI(n_25));
  ADDFX1 cdnfadd_000_1(.CO(n_108), .S(n_107), .A(n_33), .B(n_133), .CI(n_21));
  ADDFX1 cdnfadd_000_2(.CO(n_132), .S(n_131), .A(in_22[0]), .B(n_29), .CI(
    in_42[0]));
  ADDFX1 cdnfadd_000_3(.CO(n_130), .S(n_129), .A(n_5), .B(in_20[0]), .CI(in_3[0]));
  ADDFX1 cdnfadd_000_4(.CO(n_128), .S(n_127), .A(n_20), .B(n_4), .CI(in_39[0]));
  ADDFX1 cdnfadd_000_5(.CO(n_126), .S(n_125), .A(in_31[0]), .B(in_10[0]), .CI(
    n_16));
  ADDFX1 cdnfadd_000_6(.CO(n_124), .S(n_123), .A(in_18), .B(n_1), .CI(in_36[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_122), .S(n_121), .A(in_5[0]), .B(n_18), .CI(
    in_17[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_120), .S(n_119), .A(n_2), .B(in_19), .CI(in_8[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_89), .S(n_88), .A(in_12[0]), .B(in_11[0]), .CI(
    n_107));
  ADDFX1 cdnfadd_000_10(.CO(n_106), .S(n_135), .A(n_125), .B(n_127), .CI(n_131));
  ADDFX1 cdnfadd_000_11(.CO(n_105), .S(n_142), .A(n_123), .B(in_1[0]), .CI(n_129));
  ADDFX1 cdnfadd_000_12(.CO(n_74), .S(n_136), .A(n_121), .B(n_119), .CI(n_88));
  ADDFX1 cdnfadd_001_1(.CO(n_95), .S(n_104), .A(n_31), .B(n_134), .CI(n_32));
  ADDFX1 cdnfadd_001_2(.CO(n_94), .S(n_93), .A(n_104), .B(n_23), .CI(n_9));
  ADDFX1 cdnfadd_001_3(.CO(n_118), .S(n_117), .A(n_17), .B(n_28), .CI(in_32[1]));
  ADDFX1 cdnfadd_001_4(.CO(n_116), .S(n_115), .A(in_5[1]), .B(n_11), .CI(
    in_29[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_114), .S(n_113), .A(in_36[0]), .B(n_7), .CI(
    in_16[1]));
  ADDFX1 cdnfadd_001_6(.CO(n_112), .S(n_111), .A(n_19), .B(in_12[1]), .CI(n_8));
  ADDFX1 cdnfadd_001_7(.CO(n_103), .S(n_102), .A(n_6), .B(in_10[1]), .CI(n_122));
  ADDFX1 cdnfadd_001_8(.CO(n_87), .S(n_86), .A(n_132), .B(n_108), .CI(n_130));
  ADDFX1 cdnfadd_001_9(.CO(n_101), .S(n_100), .A(n_126), .B(n_124), .CI(n_128));
  ADDFX1 cdnfadd_001_10(.CO(n_80), .S(n_79), .A(n_113), .B(in_1[1]), .CI(n_93));
  ADDFX1 cdnfadd_001_11(.CO(n_99), .S(n_98), .A(n_117), .B(n_115), .CI(n_120));
  ADDFX1 cdnfadd_001_12(.CO(n_73), .S(n_72), .A(n_111), .B(n_89), .CI(n_102));
  ADDFX1 cdnfadd_001_13(.CO(n_85), .S(n_84), .A(n_105), .B(n_100), .CI(n_106));
  ADDFX1 cdnfadd_001_14(.CO(n_65), .S(n_143), .A(n_86), .B(n_98), .CI(n_79));
  ADDFX1 cdnfadd_001_15(.CO(n_144), .S(n_137), .A(n_74), .B(n_72), .CI(n_84));
  ADDFX1 cdnfadd_002_1(.CO(n_92), .S(n_91), .A(n_35), .B(n_12), .CI(n_15));
  ADDFX1 cdnfadd_002_2(.CO(n_110), .S(n_109), .A(n_14), .B(n_22), .CI(n_3));
  ADDFX1 cdnfadd_002_3(.CO(n_78), .S(n_77), .A(in_5[2]), .B(n_94), .CI(n_116));
  ADDFX1 cdnfadd_002_4(.CO(n_76), .S(n_75), .A(n_118), .B(n_114), .CI(n_91));
  ADDFX1 cdnfadd_002_5(.CO(n_97), .S(n_96), .A(n_112), .B(n_27), .CI(n_109));
  ADDFX1 cdnfadd_002_6(.CO(n_71), .S(n_70), .A(n_103), .B(n_101), .CI(n_87));
  ADDFX1 cdnfadd_002_7(.CO(n_69), .S(n_68), .A(n_80), .B(n_77), .CI(n_75));
  ADDFX1 cdnfadd_002_8(.CO(n_64), .S(n_63), .A(n_96), .B(n_99), .CI(n_73));
  ADDFX1 cdnfadd_002_9(.CO(n_59), .S(n_58), .A(n_85), .B(n_70), .CI(n_65));
  ADDFX1 cdnfadd_002_10(.CO(n_145), .S(n_138), .A(n_68), .B(n_63), .CI(n_58));
  ADDFX1 cdnfadd_003_0(.CO(n_83), .S(n_90), .A(n_13), .B(n_34), .CI(in_36[0]));
  ADDFX1 cdnfadd_003_1(.CO(n_82), .S(n_81), .A(n_24), .B(n_92), .CI(n_90));
  ADDFX1 cdnfadd_003_2(.CO(n_67), .S(n_66), .A(n_110), .B(n_78), .CI(n_76));
  ADDFX1 cdnfadd_003_3(.CO(n_62), .S(n_61), .A(n_81), .B(n_97), .CI(n_71));
  ADDFX1 cdnfadd_003_4(.CO(n_57), .S(n_56), .A(n_66), .B(n_69), .CI(n_64));
  ADDFX1 cdnfadd_003_5(.CO(n_146), .S(n_139), .A(n_61), .B(n_59), .CI(n_56));
  ADDFX1 cdnfadd_004_0(.CO(n_55), .S(n_60), .A(n_38), .B(n_82), .CI(n_67));
  ADDFX1 cdnfadd_004_1(.CO(n_141), .S(n_140), .A(n_62), .B(n_60), .CI(n_57));
  OA21X1 g328(.Y(out_0[6]), .A0(n_43), .A1(n_52), .B0(out_0[9]));
  NAND2X1 g329(.Y(out_0[9]), .A(n_43), .B(n_52));
  ADDFX1 g330(.CO(n_52), .S(out_0[5]), .A(n_44), .B(n_141), .CI(n_49));
  ADDFX1 g331(.CO(n_49), .S(out_0[4]), .A(n_146), .B(n_140), .CI(n_47));
  ADDFX1 g332(.CO(n_47), .S(out_0[3]), .A(n_145), .B(n_139), .CI(n_45));
  ADDFX1 g333(.CO(n_45), .S(out_0[2]), .A(n_144), .B(n_41), .CI(n_138));
  OAI2BB1X1 g334(.Y(n_44), .A0N(n_37), .A1N(n_55), .B0(n_43));
  OR2X1 g335(.Y(n_43), .A(n_37), .B(n_55));
  ADDFX1 g336(.CO(n_41), .S(out_0[1]), .A(n_39), .B(n_143), .CI(n_137));
  ADDFX1 g337(.CO(n_39), .S(out_0[0]), .A(n_135), .B(n_142), .CI(n_136));
  AOI21X1 g338(.Y(n_38), .A0(in_36[0]), .A1(n_36), .B0(n_37));
  NOR2X1 g339(.Y(n_37), .A(in_36[0]), .B(n_36));
  INVX1 g340(.Y(n_36), .A(n_83));
  OAI2BB1X1 g341(.Y(n_35), .A0N(n_30), .A1N(n_95), .B0(n_34));
  OR2X1 g342(.Y(n_34), .A(n_30), .B(n_95));
  AOI21X1 g343(.Y(n_33), .A0(in_7[0]), .A1(in_4[0]), .B0(n_31));
  OAI21X1 g344(.Y(n_32), .A0(in_9[1]), .A1(n_13), .B0(n_30));
  NOR2X1 g345(.Y(n_31), .A(in_7[0]), .B(in_4[0]));
  NAND2X1 g346(.Y(n_30), .A(in_9[1]), .B(n_13));
  INVX1 g347(.Y(n_29), .A(in_33[0]));
  INVX1 g348(.Y(n_28), .A(in_0[1]));
  INVX1 g349(.Y(n_27), .A(in_1[2]));
  INVX1 g350(.Y(n_26), .A(in_2[0]));
  INVX1 g351(.Y(n_25), .A(in_13[0]));
  INVX1 g352(.Y(n_24), .A(in_5[3]));
  INVX1 g353(.Y(n_23), .A(in_30[1]));
  INVX1 g354(.Y(n_22), .A(in_10[2]));
  INVX1 g355(.Y(n_21), .A(in_34[0]));
  INVX1 g356(.Y(n_20), .A(in_27[0]));
  INVX1 g357(.Y(n_19), .A(in_40[1]));
  INVX1 g358(.Y(n_18), .A(in_23[0]));
  INVX1 g359(.Y(n_17), .A(in_28[1]));
  INVX1 g360(.Y(n_16), .A(in_21[0]));
  INVX1 g361(.Y(n_15), .A(in_42[0]));
  INVX1 g362(.Y(n_14), .A(in_31[0]));
  INVX1 g363(.Y(n_13), .A(in_14[1]));
  INVX1 g364(.Y(n_12), .A(in_25[2]));
  INVX1 g365(.Y(n_11), .A(in_24[1]));
  INVX1 g366(.Y(n_10), .A(in_6[0]));
  INVX1 g367(.Y(n_9), .A(in_38[1]));
  INVX1 g368(.Y(n_8), .A(in_11[1]));
  INVX1 g369(.Y(n_7), .A(in_37[1]));
  INVX1 g370(.Y(n_6), .A(in_8[1]));
  INVX1 g371(.Y(n_5), .A(in_26[0]));
  INVX1 g372(.Y(n_4), .A(in_41[0]));
  INVX1 g373(.Y(n_3), .A(in_12[2]));
  INVX1 g374(.Y(n_2), .A(in_15[0]));
  INVX1 g375(.Y(n_1), .A(in_35[0]));
endmodule

module WALLACE_CSA_DUMMY_OP40_group_359279(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, out_0);
input  in_28, in_33, in_34;
input   [4:0] in_0;
input   [6:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [2:0] in_6;
input   [4:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [4:0] in_14;
input   [4:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [1:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [2:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [2:0] in_27;
input   [1:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
output  [9:0] out_0;
wire  n_124, n_121, n_119, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_103, n_102, n_101, n_100, n_99, 
    n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_34, 
    in_33, in_28;
wire   [9:0] out_0;
wire   [1:0] in_35;
wire   [1:0] in_29;
wire   [1:0] in_26;
wire   [1:0] in_19;
wire   [2:0] in_37;
wire   [2:0] in_27;
wire   [2:0] in_23;
wire   [2:0] in_6;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [6:0] in_1;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_15;
wire   [4:0] in_14;
wire   [4:0] in_7;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  OA21X1 g1474(.Y(out_0[6]), .A0(n_107), .A1(n_124), .B0(out_0[9]));
  NAND2X1 g1475(.Y(out_0[9]), .A(n_107), .B(n_124));
  ADDFX1 g1476(.CO(n_124), .S(out_0[5]), .A(n_110), .B(n_115), .CI(n_121));
  ADDFX1 g1477(.CO(n_121), .S(out_0[4]), .A(n_116), .B(n_113), .CI(n_119));
  ADDFX1 g1478(.CO(n_119), .S(out_0[3]), .A(n_108), .B(n_114), .CI(n_117));
  ADDFX1 g1479(.CO(n_117), .S(out_0[2]), .A(n_100), .B(n_103), .CI(n_109));
  ADDFX1 g1480(.CO(n_115), .S(n_116), .A(n_101), .B(n_105), .CI(n_111));
  ADDFX1 g1481(.CO(n_113), .S(n_114), .A(n_102), .B(n_99), .CI(n_112));
  ADDFX1 g1482(.CO(n_111), .S(n_112), .A(n_91), .B(n_98), .CI(n_95));
  OAI2BB1X1 g1483(.Y(n_110), .A0N(n_83), .A1N(n_106), .B0(n_107));
  ADDFX1 g1484(.CO(n_108), .S(n_109), .A(n_92), .B(n_96), .CI(n_89));
  OR2X1 g1485(.Y(n_107), .A(n_83), .B(n_106));
  ADDFX1 g1486(.CO(n_106), .S(n_105), .A(n_63), .B(n_88), .CI(n_97));
  ADDFX1 g1487(.CO(n_103), .S(out_0[1]), .A(n_86), .B(n_90), .CI(n_94));
  ADDFX1 g1488(.CO(n_101), .S(n_102), .A(n_64), .B(n_84), .CI(n_77));
  ADDFX1 g1489(.CO(n_99), .S(n_100), .A(n_78), .B(n_79), .CI(n_93));
  ADDFX1 g1490(.CO(n_97), .S(n_98), .A(n_61), .B(n_73), .CI(n_81));
  ADDFX1 g1491(.CO(n_95), .S(n_96), .A(n_71), .B(n_69), .CI(n_85));
  ADDFX1 g1492(.CO(n_93), .S(n_94), .A(n_65), .B(n_72), .CI(n_76));
  ADDFX1 g1493(.CO(n_91), .S(n_92), .A(n_62), .B(n_74), .CI(n_75));
  ADDFX1 g1494(.CO(n_89), .S(n_90), .A(n_58), .B(n_70), .CI(n_80));
  OAI2BB1X1 g1495(.Y(n_88), .A0N(n_52), .A1N(n_82), .B0(n_83));
  ADDFX1 g1496(.CO(n_86), .S(out_0[0]), .A(n_56), .B(n_68), .CI(n_66));
  ADDFX1 g1497(.CO(n_84), .S(n_85), .A(n_44), .B(n_26), .CI(n_60));
  OR2X1 g1498(.Y(n_83), .A(n_52), .B(n_82));
  ADDFX1 g1499(.CO(n_82), .S(n_81), .A(n_1), .B(n_53), .CI(n_59));
  ADDFX1 g1500(.CO(n_79), .S(n_80), .A(n_48), .B(n_67), .CI(n_24));
  ADDFX1 g1501(.CO(n_77), .S(n_78), .A(n_47), .B(n_23), .CI(n_57));
  ADDFX1 g1502(.CO(n_75), .S(n_76), .A(n_45), .B(n_41), .CI(n_54));
  ADDFX1 g1503(.CO(n_73), .S(n_74), .A(n_29), .B(in_2[2]), .CI(n_51));
  ADDFX1 g1504(.CO(n_71), .S(n_72), .A(n_35), .B(n_37), .CI(n_50));
  ADDFX1 g1505(.CO(n_69), .S(n_70), .A(n_30), .B(n_18), .CI(n_55));
  ADDFX1 g1506(.CO(n_67), .S(n_68), .A(n_38), .B(n_36), .CI(n_22));
  ADDFX1 g1507(.CO(n_65), .S(n_66), .A(n_42), .B(n_46), .CI(n_34));
  ADDFX1 g1508(.CO(n_63), .S(n_64), .A(n_43), .B(n_19), .CI(n_25));
  ADDFX1 g1509(.CO(n_61), .S(n_62), .A(n_17), .B(n_49), .CI(n_20));
  ADDFX1 g1510(.CO(n_59), .S(n_60), .A(n_9), .B(n_3), .CI(n_39));
  ADDFX1 g1511(.CO(n_57), .S(n_58), .A(n_33), .B(n_21), .CI(in_1[1]));
  ADDFX1 g1512(.CO(n_55), .S(n_56), .A(in_2[0]), .B(n_16), .CI(in_12[0]));
  OAI21X1 g1513(.Y(n_54), .A0(in_24[1]), .A1(n_40), .B0(n_51));
  XOR2XL g1514(.Y(n_53), .A(in_2[3]), .B(n_39));
  NOR2X1 g1515(.Y(n_52), .A(in_2[3]), .B(n_39));
  NAND2X1 g1516(.Y(n_51), .A(in_24[1]), .B(n_40));
  ADDFX1 g1517(.CO(n_49), .S(n_50), .A(in_6[1]), .B(in_37[1]), .CI(n_12));
  ADDFX1 g1518(.CO(n_47), .S(n_48), .A(n_15), .B(in_12[1]), .CI(in_10[1]));
  ADDFX1 g1519(.CO(n_45), .S(n_46), .A(in_19[0]), .B(in_17[0]), .CI(in_36[0]));
  ADDFX1 g1520(.CO(n_43), .S(n_44), .A(in_27[2]), .B(n_5), .CI(n_7));
  ADDFX1 g1521(.CO(n_41), .S(n_42), .A(in_28), .B(n_6), .CI(in_1[0]));
  ADDFX1 g1522(.CO(n_39), .S(n_40), .A(in_4[1]), .B(in_8[1]), .CI(in_9[1]));
  ADDFX1 g1523(.CO(n_37), .S(n_38), .A(in_10[0]), .B(in_26[0]), .CI(in_29[0]));
  ADDFX1 g1524(.CO(n_35), .S(n_36), .A(n_13), .B(in_35[0]), .CI(in_9[0]));
  INVX1 g1525(.Y(n_34), .A(n_32));
  INVX1 g1526(.Y(n_33), .A(n_31));
  ADDFX1 g1527(.CO(n_31), .S(n_32), .A(in_20[0]), .B(in_16[0]), .CI(in_32[0]));
  INVX1 g1528(.Y(n_30), .A(n_28));
  INVX1 g1529(.Y(n_29), .A(n_27));
  ADDFX1 g1530(.CO(n_27), .S(n_28), .A(in_15[1]), .B(in_25[1]), .CI(in_31[1]));
  ADDFX1 g1531(.CO(n_25), .S(n_26), .A(in_12[2]), .B(n_11), .CI(n_14));
  ADDFX1 g1532(.CO(n_23), .S(n_24), .A(n_8), .B(in_5[1]), .CI(in_2[1]));
  ADDFX1 g1533(.CO(n_21), .S(n_22), .A(in_5[0]), .B(in_33), .CI(in_34));
  ADDFX1 g1534(.CO(n_19), .S(n_20), .A(in_11[2]), .B(n_2), .CI(n_10));
  ADDFX1 g1535(.CO(n_17), .S(n_18), .A(in_13[1]), .B(in_23[1]), .CI(n_4));
  MXI2XL g1536(.Y(n_16), .A(in_18[0]), .B(n_9), .S0(in_3[0]));
  NOR2X1 g1537(.Y(n_15), .A(in_3[0]), .B(n_9));
  INVX1 g1538(.Y(n_14), .A(in_1[2]));
  INVX1 g1539(.Y(n_13), .A(in_30[0]));
  INVX1 g1540(.Y(n_12), .A(in_7[1]));
  INVX1 g1541(.Y(n_11), .A(in_10[2]));
  INVX1 g1542(.Y(n_10), .A(in_5[2]));
  INVX1 g1543(.Y(n_9), .A(in_18[0]));
  INVX1 g1544(.Y(n_8), .A(in_22[1]));
  INVX1 g1545(.Y(n_7), .A(in_38[2]));
  INVX1 g1546(.Y(n_6), .A(in_0[0]));
  INVX1 g1547(.Y(n_5), .A(in_21[2]));
  INVX1 g1548(.Y(n_4), .A(in_14[1]));
  INVX1 g1549(.Y(n_3), .A(in_36[0]));
  INVX1 g1550(.Y(n_2), .A(in_17[0]));
  INVX1 g1551(.Y(n_1), .A(in_12[1]));
endmodule

module WALLACE_CSA_DUMMY_OP43_group_359277(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    out_0);
input  in_25, in_31;
input   [4:0] in_0;
input   [6:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [4:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [4:0] in_11;
input   [4:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [1:0] in_24;
input   [4:0] in_26;
input   [2:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [1:0] in_30;
input   [2:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [4:0] in_37;
output  [9:0] out_0;
wire  n_118, n_116, n_114, n_112, n_111, n_110, n_108, n_107, n_106, n_105, 
    n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_94, n_93, 
    n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, 
    n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, 
    n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, 
    n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
    n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, 
    n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, 
    n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, 
    n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_31, in_25;
wire   [9:0] out_0;
wire   [2:0] in_36;
wire   [2:0] in_34;
wire   [2:0] in_32;
wire   [2:0] in_27;
wire   [1:0] in_30;
wire   [1:0] in_24;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [6:0] in_1;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_12;
wire   [4:0] in_11;
wire   [4:0] in_6;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3589(.Y(out_0[9]), .A(n_118));
  ADDFX1 g3590(.CO(n_118), .S(out_0[5]), .A(n_80), .B(n_104), .CI(n_116));
  ADDFX1 g3591(.CO(n_116), .S(out_0[4]), .A(n_105), .B(n_106), .CI(n_114));
  ADDFX1 g3592(.CO(n_114), .S(out_0[3]), .A(n_110), .B(n_107), .CI(n_112));
  ADDFX1 g3593(.CO(n_112), .S(out_0[2]), .A(n_102), .B(n_108), .CI(n_111));
  ADDFX1 g3594(.CO(n_110), .S(n_111), .A(n_97), .B(n_83), .CI(n_99));
  ADDFX1 g3595(.CO(n_108), .S(out_0[1]), .A(n_89), .B(n_94), .CI(n_103));
  ADDFX1 g3596(.CO(n_106), .S(n_107), .A(n_96), .B(n_98), .CI(n_101));
  ADDFX1 g3597(.CO(n_104), .S(n_105), .A(n_81), .B(n_92), .CI(n_100));
  ADDFX1 g3598(.CO(n_102), .S(n_103), .A(n_71), .B(n_85), .CI(n_87));
  ADDFX1 g3599(.CO(n_100), .S(n_101), .A(n_90), .B(n_82), .CI(n_93));
  ADDFX1 g3600(.CO(n_98), .S(n_99), .A(n_86), .B(n_88), .CI(n_84));
  ADDFX1 g3601(.CO(n_96), .S(n_97), .A(n_65), .B(n_62), .CI(n_91));
  ADDFX1 g3602(.CO(n_94), .S(out_0[0]), .A(n_74), .B(n_78), .CI(n_72));
  ADDFX1 g3603(.CO(n_92), .S(n_93), .A(n_61), .B(n_63), .CI(n_79));
  ADDFX1 g3604(.CO(n_90), .S(n_91), .A(n_75), .B(n_59), .CI(n_67));
  ADDFX1 g3605(.CO(n_88), .S(n_89), .A(n_76), .B(n_68), .CI(n_66));
  ADDFX1 g3606(.CO(n_86), .S(n_87), .A(n_60), .B(n_77), .CI(n_55));
  ADDFX1 g3607(.CO(n_84), .S(n_85), .A(n_28), .B(n_73), .CI(n_58));
  ADDFX1 g3608(.CO(n_82), .S(n_83), .A(n_70), .B(n_64), .CI(n_57));
  INVX1 g3609(.Y(n_81), .A(n_80));
  ADDFX1 g3610(.CO(n_80), .S(n_79), .A(n_45), .B(n_69), .CI(n_4));
  ADDFX1 g3611(.CO(n_77), .S(n_78), .A(n_48), .B(n_52), .CI(n_54));
  ADDFX1 g3612(.CO(n_75), .S(n_76), .A(n_31), .B(n_47), .CI(n_51));
  ADDFX1 g3613(.CO(n_73), .S(n_74), .A(n_32), .B(n_40), .CI(n_26));
  ADDFX1 g3614(.CO(n_71), .S(n_72), .A(n_22), .B(n_36), .CI(n_56));
  ADDFX1 g3615(.CO(n_69), .S(n_70), .A(in_36[1]), .B(n_41), .CI(n_49));
  ADDFX1 g3616(.CO(n_67), .S(n_68), .A(n_42), .B(n_20), .CI(n_30));
  ADDFX1 g3617(.CO(n_65), .S(n_66), .A(n_50), .B(n_34), .CI(n_35));
  ADDFX1 g3618(.CO(n_63), .S(n_64), .A(n_29), .B(n_33), .CI(in_2[2]));
  ADDFX1 g3619(.CO(n_61), .S(n_62), .A(n_46), .B(n_19), .CI(n_27));
  ADDFX1 g3620(.CO(n_59), .S(n_60), .A(n_53), .B(n_25), .CI(n_21));
  ADDFX1 g3621(.CO(n_57), .S(n_58), .A(n_43), .B(n_39), .CI(in_2[1]));
  ADDFX1 g3622(.CO(n_55), .S(n_56), .A(in_16[0]), .B(n_44), .CI(in_2[0]));
  ADDFX1 g3623(.CO(n_53), .S(n_54), .A(in_7[0]), .B(n_14), .CI(in_23[0]));
  ADDFX1 g3624(.CO(n_51), .S(n_52), .A(in_24[0]), .B(n_16), .CI(in_27[0]));
  ADDFX1 g3625(.CO(n_49), .S(n_50), .A(in_24[0]), .B(in_27[0]), .CI(in_1[0]));
  ADDFX1 g3626(.CO(n_47), .S(n_48), .A(in_8[0]), .B(in_25), .CI(n_11));
  INVX1 g3627(.Y(n_46), .A(n_38));
  INVX1 g3628(.Y(n_45), .A(n_37));
  INVX1 g3629(.Y(n_44), .A(n_24));
  INVX1 g3630(.Y(n_43), .A(n_23));
  ADDFX1 g3631(.CO(n_41), .S(n_42), .A(in_3[1]), .B(n_12), .CI(n_8));
  ADDFX1 g3632(.CO(n_39), .S(n_40), .A(in_17[0]), .B(n_18), .CI(in_1[0]));
  ADDFX1 g3633(.CO(n_37), .S(n_38), .A(in_5[0]), .B(in_23[0]), .CI(in_15[2]));
  ADDFX1 g3634(.CO(n_35), .S(n_36), .A(in_31), .B(in_34[0]), .CI(in_10[0]));
  ADDFX1 g3635(.CO(n_33), .S(n_34), .A(in_34[0]), .B(n_3), .CI(n_9));
  ADDFX1 g3636(.CO(n_31), .S(n_32), .A(n_7), .B(n_13), .CI(in_32[0]));
  ADDFX1 g3637(.CO(n_29), .S(n_30), .A(n_6), .B(n_15), .CI(in_32[0]));
  ADDFX1 g3638(.CO(n_27), .S(n_28), .A(n_10), .B(in_10[1]), .CI(in_15[1]));
  ADDFX1 g3639(.CO(n_25), .S(n_26), .A(in_9[0]), .B(n_5), .CI(n_17));
  ADDFX1 g3640(.CO(n_23), .S(n_24), .A(in_12[0]), .B(in_4[0]), .CI(in_37[0]));
  ADDFX1 g3641(.CO(n_21), .S(n_22), .A(n_1), .B(in_5[0]), .CI(in_15[0]));
  ADDFX1 g3642(.CO(n_19), .S(n_20), .A(n_2), .B(in_30[1]), .CI(in_16[1]));
  INVX1 g3643(.Y(n_18), .A(in_26[0]));
  INVX1 g3644(.Y(n_17), .A(in_33[0]));
  INVX1 g3645(.Y(n_16), .A(in_14[0]));
  INVX1 g3646(.Y(n_15), .A(in_29[1]));
  INVX1 g3647(.Y(n_14), .A(in_0[0]));
  INVX1 g3648(.Y(n_13), .A(in_22[0]));
  INVX1 g3649(.Y(n_12), .A(in_11[1]));
  INVX1 g3650(.Y(n_11), .A(in_19[0]));
  INVX1 g3651(.Y(n_10), .A(in_36[1]));
  INVX1 g3652(.Y(n_9), .A(in_35[1]));
  INVX1 g3653(.Y(n_8), .A(in_20[1]));
  INVX1 g3654(.Y(n_7), .A(in_21[0]));
  INVX1 g3655(.Y(n_6), .A(in_6[1]));
  INVX1 g3656(.Y(n_5), .A(in_18[0]));
  INVX1 g3657(.Y(n_4), .A(in_2[3]));
  INVX1 g3658(.Y(n_3), .A(in_9[1]));
  INVX1 g3659(.Y(n_2), .A(in_28[1]));
  INVX1 g3660(.Y(n_1), .A(in_13[0]));
endmodule

module WALLACE_CSA_DUMMY_OP50_group_359285(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, out_0);
input  in_18, in_33;
input   [4:0] in_0;
input   [5:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [4:0] in_15;
input   [1:0] in_16;
input   [4:0] in_17;
input   [1:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [1:0] in_26;
input   [4:0] in_27;
input   [2:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [1:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [2:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [2:0] in_43;
output  [9:0] out_0;
wire  n_118, n_116, n_114, n_113, n_112, n_110, n_109, n_108, n_106, n_105, 
    n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, 
    n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, 
    n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, 
    n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, 
    n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
    n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, 
    n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, 
    n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, 
    n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_33, in_18;
wire   [9:0] out_0;
wire   [2:0] in_43;
wire   [2:0] in_40;
wire   [2:0] in_39;
wire   [2:0] in_36;
wire   [2:0] in_28;
wire   [1:0] in_34;
wire   [1:0] in_31;
wire   [1:0] in_29;
wire   [1:0] in_26;
wire   [1:0] in_25;
wire   [1:0] in_19;
wire   [1:0] in_16;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [5:0] in_1;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_27;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_17;
wire   [4:0] in_15;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3619(.Y(out_0[9]), .A(n_118));
  ADDFX1 g3620(.CO(n_118), .S(out_0[5]), .A(n_81), .B(n_108), .CI(n_116));
  ADDFX1 g3621(.CO(n_116), .S(out_0[4]), .A(n_109), .B(n_112), .CI(n_114));
  ADDFX1 g3622(.CO(n_114), .S(out_0[3]), .A(n_104), .B(n_113), .CI(n_110));
  ADDFX1 g3623(.CO(n_112), .S(n_113), .A(n_96), .B(n_102), .CI(n_101));
  ADDFX1 g3624(.CO(n_110), .S(out_0[2]), .A(n_103), .B(n_106), .CI(n_105));
  ADDFX1 g3625(.CO(n_108), .S(n_109), .A(n_71), .B(n_90), .CI(n_100));
  ADDFX1 g3626(.CO(n_106), .S(out_0[1]), .A(n_92), .B(n_95), .CI(n_99));
  ADDFX1 g3627(.CO(n_104), .S(n_105), .A(n_89), .B(n_97), .CI(n_98));
  ADDFX1 g3628(.CO(n_102), .S(n_103), .A(n_87), .B(n_84), .CI(n_94));
  ADDFX1 g3629(.CO(n_100), .S(n_101), .A(n_86), .B(n_88), .CI(n_91));
  ADDFX1 g3630(.CO(n_98), .S(n_99), .A(n_76), .B(n_83), .CI(n_85));
  ADDFX1 g3631(.CO(n_96), .S(n_97), .A(n_66), .B(n_73), .CI(n_82));
  ADDFX1 g3632(.CO(n_94), .S(n_95), .A(n_58), .B(n_75), .CI(n_79));
  ADDFX1 g3633(.CO(n_92), .S(out_0[0]), .A(n_60), .B(n_70), .CI(n_77));
  ADDFX1 g3634(.CO(n_90), .S(n_91), .A(n_65), .B(n_72), .CI(n_80));
  ADDFX1 g3635(.CO(n_88), .S(n_89), .A(n_63), .B(n_74), .CI(n_78));
  ADDFX1 g3636(.CO(n_86), .S(n_87), .A(n_67), .B(n_57), .CI(n_61));
  ADDFX1 g3637(.CO(n_84), .S(n_85), .A(n_68), .B(n_69), .CI(n_59));
  ADDFX1 g3638(.CO(n_82), .S(n_83), .A(n_36), .B(n_55), .CI(n_62));
  INVX1 g3639(.Y(n_81), .A(n_71));
  XNOR2X1 g3640(.Y(n_80), .A(n_37), .B(n_64));
  ADDFX1 g3641(.CO(n_78), .S(n_79), .A(n_42), .B(n_46), .CI(n_50));
  ADDFX1 g3642(.CO(n_76), .S(n_77), .A(n_23), .B(n_54), .CI(n_56));
  ADDFX1 g3643(.CO(n_74), .S(n_75), .A(n_48), .B(n_40), .CI(n_27));
  ADDFX1 g3644(.CO(n_72), .S(n_73), .A(n_41), .B(n_38), .CI(n_35));
  NAND2BX1 g3645(.Y(n_71), .AN(n_37), .B(n_64));
  ADDFX1 g3646(.CO(n_69), .S(n_70), .A(n_15), .B(n_32), .CI(n_25));
  ADDFX1 g3647(.CO(n_67), .S(n_68), .A(n_53), .B(n_20), .CI(n_24));
  ADDFX1 g3648(.CO(n_65), .S(n_66), .A(n_45), .B(n_39), .CI(n_26));
  ADDFX1 g3649(.CO(n_64), .S(n_63), .A(n_6), .B(n_49), .CI(n_47));
  ADDFX1 g3650(.CO(n_61), .S(n_62), .A(n_43), .B(n_22), .CI(n_18));
  ADDFX1 g3651(.CO(n_59), .S(n_60), .A(n_44), .B(n_21), .CI(n_19));
  ADDFX1 g3652(.CO(n_57), .S(n_58), .A(n_29), .B(n_14), .CI(n_31));
  ADDFX1 g3653(.CO(n_55), .S(n_56), .A(in_6[0]), .B(in_8[0]), .CI(n_30));
  INVX1 g3654(.Y(n_54), .A(n_52));
  INVX1 g3655(.Y(n_53), .A(n_51));
  ADDFX1 g3656(.CO(n_51), .S(n_52), .A(in_22[0]), .B(in_32[0]), .CI(in_41[0]));
  ADDFX1 g3657(.CO(n_49), .S(n_50), .A(in_39[1]), .B(in_40[1]), .CI(n_3));
  ADDFX1 g3658(.CO(n_47), .S(n_48), .A(in_11[1]), .B(in_43[1]), .CI(in_36[0]));
  ADDFX1 g3659(.CO(n_45), .S(n_46), .A(n_4), .B(n_2), .CI(in_19[1]));
  ADDFX1 g3660(.CO(n_43), .S(n_44), .A(in_1[0]), .B(in_18), .CI(n_10));
  ADDFX1 g3661(.CO(n_41), .S(n_42), .A(in_28[0]), .B(n_12), .CI(in_34[1]));
  INVX1 g3662(.Y(n_40), .A(n_34));
  INVX1 g3663(.Y(n_39), .A(n_33));
  INVX1 g3664(.Y(n_38), .A(n_28));
  INVX1 g3665(.Y(n_36), .A(n_17));
  INVX1 g3666(.Y(n_35), .A(n_16));
  ADDFX1 g3667(.CO(n_33), .S(n_34), .A(in_5[1]), .B(in_35[1]), .CI(in_38[1]));
  ADDFX1 g3668(.CO(n_31), .S(n_32), .A(in_7[0]), .B(n_5), .CI(in_25[0]));
  ADDFX1 g3669(.CO(n_29), .S(n_30), .A(n_8), .B(n_11), .CI(in_31[0]));
  ADDFX1 g3670(.CO(n_37), .S(n_28), .A(in_23[2]), .B(in_21[2]), .CI(in_27[0]));
  ADDFX1 g3671(.CO(n_26), .S(n_27), .A(in_25[0]), .B(n_7), .CI(in_26[1]));
  ADDFX1 g3672(.CO(n_24), .S(n_25), .A(in_13[0]), .B(in_11[0]), .CI(in_27[0]));
  ADDFX1 g3673(.CO(n_22), .S(n_23), .A(in_4[0]), .B(n_1), .CI(n_13));
  ADDFX1 g3674(.CO(n_20), .S(n_21), .A(in_16[0]), .B(in_36[0]), .CI(n_9));
  ADDFX1 g3675(.CO(n_18), .S(n_19), .A(in_10[0]), .B(in_5[0]), .CI(in_29[0]));
  ADDFX1 g3676(.CO(n_16), .S(n_17), .A(in_12[1]), .B(in_8[1]), .CI(in_6[1]));
  ADDFX1 g3677(.CO(n_14), .S(n_15), .A(in_28[0]), .B(in_14[0]), .CI(in_33));
  INVX1 g3678(.Y(n_13), .A(in_15[0]));
  INVX1 g3679(.Y(n_12), .A(in_20[1]));
  INVX1 g3680(.Y(n_11), .A(in_30[0]));
  INVX1 g3681(.Y(n_10), .A(in_37[0]));
  INVX1 g3682(.Y(n_9), .A(in_42[0]));
  INVX1 g3683(.Y(n_8), .A(in_3[0]));
  INVX1 g3684(.Y(n_7), .A(in_1[1]));
  INVX1 g3685(.Y(n_6), .A(in_2[2]));
  INVX1 g3686(.Y(n_5), .A(in_24[0]));
  INVX1 g3687(.Y(n_4), .A(in_17[1]));
  INVX1 g3688(.Y(n_3), .A(in_0[1]));
  INVX1 g3689(.Y(n_2), .A(in_7[1]));
  INVX1 g3690(.Y(n_1), .A(in_9[0]));
endmodule

module WALLACE_CSA_DUMMY_OP58_group_109825_6338(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, in_39, in_40, in_41, out_0);
input  in_27, in_28, in_32, in_40;
input   [4:0] in_0;
input   [2:0] in_1;
input   [9:0] in_2;
input   [6:0] in_3;
input   [6:0] in_4;
input   [2:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [4:0] in_10;
input   [4:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [4:0] in_16;
input   [3:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [1:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [2:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [4:0] in_29;
input   [4:0] in_30;
input   [2:0] in_31;
input   [4:0] in_33;
input   [1:0] in_34;
input   [2:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [2:0] in_41;
output  [9:0] out_0;
wire  n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
    n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_42, n_40, n_38, n_36, 
    n_34, n_32, n_30, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, 
    n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
    n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_40, in_32, in_28, in_27;
wire   [9:0] out_0;
wire   [1:0] in_34;
wire   [1:0] in_26;
wire   [1:0] in_21;
wire   [1:0] in_20;
wire   [3:0] in_17;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_4;
wire   [6:0] in_3;
wire   [9:0] in_2;
wire   [2:0] in_41;
wire   [2:0] in_39;
wire   [2:0] in_37;
wire   [2:0] in_35;
wire   [2:0] in_31;
wire   [2:0] in_23;
wire   [2:0] in_5;
wire   [2:0] in_1;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_16;
wire   [4:0] in_11;
wire   [4:0] in_10;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_126), .S(n_125), .A(in_32), .B(in_37[0]), .CI(
    in_30[0]));
  ADDFX1 cdnfadd_000_1(.CO(n_124), .S(n_123), .A(in_26[0]), .B(in_20[0]), .CI(
    n_19));
  ADDFX1 cdnfadd_000_2(.CO(n_122), .S(n_121), .A(in_11[0]), .B(in_19[0]), .CI(
    n_5));
  ADDFX1 cdnfadd_000_3(.CO(n_120), .S(n_119), .A(in_21[0]), .B(n_15), .CI(
    in_10[0]));
  ADDFX1 cdnfadd_000_4(.CO(n_118), .S(n_117), .A(in_40), .B(in_27), .CI(n_16));
  ADDFX1 cdnfadd_000_5(.CO(n_116), .S(n_115), .A(n_17), .B(in_28), .CI(in_14[0]));
  ADDFX1 cdnfadd_000_6(.CO(n_114), .S(n_113), .A(n_2), .B(in_39[0]), .CI(in_3[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_112), .S(n_111), .A(in_23[0]), .B(in_34[0]), .CI(
    in_9[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_110), .S(n_109), .A(in_7[0]), .B(in_33[0]), .CI(
    in_12[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_108), .S(n_107), .A(in_6[0]), .B(in_8[0]), .CI(
    in_15[0]));
  ADDFX1 cdnfadd_000_10(.CO(n_92), .S(n_127), .A(n_119), .B(n_121), .CI(n_123));
  ADDFX1 cdnfadd_000_11(.CO(n_91), .S(n_90), .A(n_115), .B(n_117), .CI(n_125));
  ADDFX1 cdnfadd_000_12(.CO(n_89), .S(n_135), .A(n_113), .B(n_111), .CI(n_109));
  ADDFX1 cdnfadd_000_13(.CO(n_72), .S(n_128), .A(n_107), .B(in_2[0]), .CI(n_90));
  ADDFX1 cdnfadd_001_0(.CO(n_106), .S(n_105), .A(in_35[1]), .B(in_5[1]), .CI(n_6));
  ADDFX1 cdnfadd_001_1(.CO(n_104), .S(n_103), .A(in_3[1]), .B(n_8), .CI(in_14[1]));
  ADDFX1 cdnfadd_001_2(.CO(n_102), .S(n_101), .A(in_1[1]), .B(n_9), .CI(in_23[0]));
  ADDFX1 cdnfadd_001_3(.CO(n_100), .S(n_99), .A(in_37[0]), .B(n_7), .CI(n_3));
  ADDFX1 cdnfadd_001_4(.CO(n_98), .S(n_97), .A(n_20), .B(in_15[1]), .CI(n_18));
  ADDFX1 cdnfadd_001_5(.CO(n_96), .S(n_95), .A(n_4), .B(n_23), .CI(n_10));
  ADDFX1 cdnfadd_001_6(.CO(n_88), .S(n_87), .A(n_14), .B(n_120), .CI(n_126));
  ADDFX1 cdnfadd_001_7(.CO(n_86), .S(n_85), .A(n_124), .B(n_122), .CI(n_116));
  ADDFX1 cdnfadd_001_8(.CO(n_84), .S(n_83), .A(n_118), .B(n_114), .CI(n_103));
  ADDFX1 cdnfadd_001_9(.CO(n_82), .S(n_81), .A(n_105), .B(n_99), .CI(n_101));
  ADDFX1 cdnfadd_001_10(.CO(n_80), .S(n_79), .A(n_112), .B(n_110), .CI(n_97));
  ADDFX1 cdnfadd_001_11(.CO(n_71), .S(n_70), .A(n_108), .B(n_95), .CI(n_92));
  ADDFX1 cdnfadd_001_12(.CO(n_69), .S(n_68), .A(n_91), .B(n_83), .CI(n_87));
  ADDFX1 cdnfadd_001_13(.CO(n_67), .S(n_66), .A(n_85), .B(n_81), .CI(n_89));
  ADDFX1 cdnfadd_001_14(.CO(n_55), .S(n_136), .A(n_79), .B(in_2[1]), .CI(n_70));
  ADDFX1 cdnfadd_001_15(.CO(n_54), .S(n_129), .A(n_72), .B(n_68), .CI(n_66));
  ADDFX1 cdnfadd_002_1(.CO(n_94), .S(n_93), .A(n_1), .B(in_41[2]), .CI(n_13));
  ADDFX1 cdnfadd_002_2(.CO(n_78), .S(n_77), .A(n_21), .B(n_104), .CI(n_102));
  ADDFX1 cdnfadd_002_3(.CO(n_76), .S(n_75), .A(n_106), .B(n_100), .CI(n_93));
  ADDFX1 cdnfadd_002_4(.CO(n_74), .S(n_73), .A(n_98), .B(n_24), .CI(n_96));
  ADDFX1 cdnfadd_002_5(.CO(n_65), .S(n_64), .A(n_86), .B(n_88), .CI(n_84));
  ADDFX1 cdnfadd_002_6(.CO(n_63), .S(n_62), .A(n_82), .B(n_77), .CI(n_75));
  ADDFX1 cdnfadd_002_7(.CO(n_59), .S(n_58), .A(n_80), .B(n_73), .CI(n_69));
  ADDFX1 cdnfadd_002_8(.CO(n_53), .S(n_52), .A(n_71), .B(n_64), .CI(in_2[2]));
  ADDFX1 cdnfadd_002_9(.CO(n_45), .S(n_137), .A(n_62), .B(n_67), .CI(n_55));
  ADDFX1 cdnfadd_002_10(.CO(n_138), .S(n_130), .A(n_58), .B(n_52), .CI(n_54));
  ADDFX1 cdnfadd_003_0(.CO(n_60), .S(n_61), .A(n_94), .B(n_22), .CI(n_78));
  ADDFX1 cdnfadd_003_1(.CO(n_57), .S(n_56), .A(n_76), .B(n_74), .CI(n_61));
  ADDFX1 cdnfadd_003_2(.CO(n_51), .S(n_50), .A(n_65), .B(n_63), .CI(in_2[3]));
  ADDFX1 cdnfadd_003_3(.CO(n_49), .S(n_48), .A(n_56), .B(n_59), .CI(n_53));
  ADDFX1 cdnfadd_003_4(.CO(n_139), .S(n_131), .A(n_50), .B(n_45), .CI(n_48));
  ADDFX1 cdnfadd_004_1(.CO(n_47), .S(n_46), .A(n_57), .B(n_27), .CI(in_2[4]));
  ADDFX1 cdnfadd_004_2(.CO(n_133), .S(n_132), .A(n_51), .B(n_46), .CI(n_49));
  ADDFX1 cdnfadd_005_0(.CO(n_134), .S(n_140), .A(in_2[5]), .B(n_26), .CI(n_47));
  INVX1 g365(.Y(out_0[9]), .A(n_42));
  ADDFX1 g366(.CO(n_42), .S(out_0[7]), .A(n_12), .B(in_2[6]), .CI(n_40));
  ADDFX1 g367(.CO(n_40), .S(out_0[6]), .A(n_11), .B(n_134), .CI(n_38));
  ADDFX1 g368(.CO(n_38), .S(out_0[5]), .A(n_140), .B(n_133), .CI(n_36));
  ADDFX1 g369(.CO(n_36), .S(out_0[4]), .A(n_139), .B(n_132), .CI(n_34));
  ADDFX1 g370(.CO(n_34), .S(out_0[3]), .A(n_138), .B(n_131), .CI(n_32));
  ADDFX1 g371(.CO(n_32), .S(out_0[2]), .A(n_30), .B(n_137), .CI(n_130));
  ADDFX1 g372(.CO(n_30), .S(out_0[1]), .A(n_28), .B(n_129), .CI(n_136));
  ADDFX1 g373(.CO(n_28), .S(out_0[0]), .A(n_127), .B(n_135), .CI(n_128));
  OAI21X1 g374(.Y(n_27), .A0(n_22), .A1(n_25), .B0(n_26));
  NAND2X1 g375(.Y(n_26), .A(n_22), .B(n_25));
  INVX1 g376(.Y(n_25), .A(n_60));
  AO21XL g377(.Y(n_24), .A0(in_31[2]), .A1(in_17[2]), .B0(n_22));
  AOI21X1 g378(.Y(n_23), .A0(in_0[1]), .A1(n_0), .B0(n_21));
  NOR2X1 g379(.Y(n_22), .A(in_31[2]), .B(in_17[2]));
  NOR2X1 g380(.Y(n_21), .A(in_0[1]), .B(n_0));
  INVX1 g381(.Y(n_20), .A(in_7[1]));
  INVX1 g382(.Y(n_19), .A(in_29[0]));
  INVX1 g383(.Y(n_18), .A(in_9[1]));
  INVX1 g384(.Y(n_17), .A(in_16[0]));
  INVX1 g385(.Y(n_16), .A(in_4[0]));
  INVX1 g386(.Y(n_15), .A(in_38[0]));
  INVX1 g387(.Y(n_14), .A(in_33[0]));
  INVX1 g388(.Y(n_13), .A(in_30[0]));
  INVX1 g389(.Y(n_12), .A(in_2[7]));
  INVX1 g390(.Y(n_11), .A(in_2[6]));
  INVX1 g391(.Y(n_10), .A(in_8[1]));
  INVX1 g392(.Y(n_9), .A(in_22[1]));
  INVX1 g393(.Y(n_8), .A(in_36[1]));
  INVX1 g394(.Y(n_7), .A(in_24[1]));
  INVX1 g395(.Y(n_6), .A(in_18[1]));
  INVX1 g396(.Y(n_5), .A(in_25[0]));
  INVX1 g397(.Y(n_4), .A(in_12[1]));
  INVX1 g398(.Y(n_3), .A(in_6[1]));
  INVX1 g399(.Y(n_2), .A(in_13[0]));
  INVX1 g400(.Y(n_1), .A(in_19[0]));
  INVX1 g401(.Y(n_0), .A(in_39[0]));
endmodule

module WALLACE_CSA_DUMMY_OP58_group_109825(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, out_0);
input  in_20, in_27, in_41;
input   [4:0] in_0;
input   [4:0] in_1;
input   [2:0] in_2;
input   [6:0] in_3;
input   [6:0] in_4;
input   [4:0] in_5;
input   [4:0] in_6;
input   [4:0] in_7;
input   [4:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [1:0] in_19;
input   [1:0] in_21;
input   [4:0] in_22;
input   [2:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [1:0] in_26;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [2:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [1:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
output  [9:0] out_0;
wire  n_122, n_120, n_118, n_116, n_115, n_114, n_113, n_112, n_111, n_110, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_41, 
    in_27, in_20;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_35;
wire   [1:0] in_26;
wire   [1:0] in_25;
wire   [1:0] in_21;
wire   [1:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [6:0] in_4;
wire   [6:0] in_3;
wire   [2:0] in_37;
wire   [2:0] in_31;
wire   [2:0] in_23;
wire   [2:0] in_2;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_8;
wire   [4:0] in_7;
wire   [4:0] in_6;
wire   [4:0] in_5;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3776(.Y(out_0[9]), .A(n_122));
  ADDFX1 g3777(.CO(n_122), .S(out_0[5]), .A(n_96), .B(n_112), .CI(n_120));
  ADDFX1 g3778(.CO(n_120), .S(out_0[4]), .A(n_113), .B(n_114), .CI(n_118));
  ADDFX1 g3779(.CO(n_118), .S(out_0[3]), .A(n_110), .B(n_115), .CI(n_116));
  ADDFX1 g3780(.CO(n_116), .S(out_0[2]), .A(n_105), .B(n_108), .CI(n_111));
  ADDFX1 g3781(.CO(n_114), .S(n_115), .A(n_101), .B(n_104), .CI(n_107));
  ADDFX1 g3782(.CO(n_112), .S(n_113), .A(n_97), .B(n_100), .CI(n_106));
  ADDFX1 g3783(.CO(n_110), .S(n_111), .A(n_86), .B(n_99), .CI(n_102));
  ADDFX1 g3784(.CO(n_108), .S(out_0[1]), .A(n_84), .B(n_87), .CI(n_103));
  ADDFX1 g3785(.CO(n_106), .S(n_107), .A(n_91), .B(n_94), .CI(n_98));
  ADDFX1 g3786(.CO(n_104), .S(n_105), .A(n_88), .B(n_93), .CI(n_95));
  ADDFX1 g3787(.CO(n_102), .S(n_103), .A(n_66), .B(n_83), .CI(n_89));
  ADDFX1 g3788(.CO(n_100), .S(n_101), .A(n_64), .B(n_80), .CI(n_92));
  ADDFX1 g3789(.CO(n_98), .S(n_99), .A(n_65), .B(n_82), .CI(n_81));
  ADDHX1 g3790(.CO(n_96), .S(n_97), .A(n_60), .B(n_90));
  ADDFX1 g3791(.CO(n_94), .S(n_95), .A(n_78), .B(n_77), .CI(n_62));
  ADDFX1 g3792(.CO(n_92), .S(n_93), .A(n_58), .B(n_73), .CI(n_70));
  ADDFX1 g3793(.CO(n_90), .S(n_91), .A(n_76), .B(n_72), .CI(n_61));
  ADDFX1 g3794(.CO(n_88), .S(n_89), .A(n_54), .B(n_79), .CI(n_69));
  ADDFX1 g3795(.CO(n_86), .S(n_87), .A(n_74), .B(n_71), .CI(n_63));
  ADDFX1 g3796(.CO(n_84), .S(out_0[0]), .A(n_55), .B(n_75), .CI(n_67));
  ADDFX1 g3797(.CO(n_82), .S(n_83), .A(n_59), .B(n_36), .CI(n_57));
  ADDFX1 g3798(.CO(n_80), .S(n_81), .A(n_56), .B(n_53), .CI(n_68));
  ADDFX1 g3799(.CO(n_78), .S(n_79), .A(n_42), .B(n_28), .CI(n_25));
  ADDFX1 g3800(.CO(n_76), .S(n_77), .A(n_19), .B(n_26), .CI(n_32));
  ADDFX1 g3801(.CO(n_74), .S(n_75), .A(n_29), .B(n_47), .CI(n_43));
  ADDFX1 g3802(.CO(n_72), .S(n_73), .A(n_24), .B(n_44), .CI(n_34));
  ADDFX1 g3803(.CO(n_70), .S(n_71), .A(n_27), .B(n_41), .CI(n_45));
  ADDFX1 g3804(.CO(n_68), .S(n_69), .A(n_22), .B(n_30), .CI(n_38));
  ADDFX1 g3805(.CO(n_66), .S(n_67), .A(n_31), .B(n_23), .CI(n_37));
  ADDFX1 g3806(.CO(n_64), .S(n_65), .A(n_21), .B(n_40), .CI(n_48));
  ADDFX1 g3807(.CO(n_62), .S(n_63), .A(n_35), .B(n_33), .CI(n_49));
  ADDFX1 g3808(.CO(n_60), .S(n_61), .A(n_9), .B(n_18), .CI(n_52));
  ADDFX1 g3809(.CO(n_58), .S(n_59), .A(n_10), .B(in_3[1]), .CI(n_46));
  ADDFX1 g3810(.CO(n_56), .S(n_57), .A(n_3), .B(n_20), .CI(in_15[1]));
  ADDFX1 g3811(.CO(n_54), .S(n_55), .A(in_1[0]), .B(in_18[0]), .CI(n_39));
  INVX1 g3812(.Y(n_53), .A(n_51));
  INVX1 g3813(.Y(n_52), .A(n_50));
  ADDFX1 g3814(.CO(n_50), .S(n_51), .A(in_6[0]), .B(in_15[2]), .CI(in_3[2]));
  ADDFX1 g3815(.CO(n_48), .S(n_49), .A(in_14[1]), .B(n_8), .CI(n_14));
  ADDFX1 g3816(.CO(n_46), .S(n_47), .A(in_13[0]), .B(in_27), .CI(in_41));
  ADDFX1 g3817(.CO(n_44), .S(n_45), .A(in_19[0]), .B(in_40[1]), .CI(n_2));
  ADDFX1 g3818(.CO(n_42), .S(n_43), .A(in_20), .B(n_16), .CI(in_26[0]));
  ADDFX1 g3819(.CO(n_40), .S(n_41), .A(in_26[0]), .B(n_6), .CI(n_17));
  ADDFX1 g3820(.CO(n_38), .S(n_39), .A(in_19[0]), .B(n_1), .CI(n_7));
  ADDFX1 g3821(.CO(n_36), .S(n_37), .A(in_11[0]), .B(in_3[0]), .CI(in_9[0]));
  ADDFX1 g3822(.CO(n_34), .S(n_35), .A(in_32[0]), .B(n_5), .CI(in_37[1]));
  ADDFX1 g3823(.CO(n_32), .S(n_33), .A(in_2[1]), .B(n_12), .CI(in_31[1]));
  ADDFX1 g3824(.CO(n_30), .S(n_31), .A(in_24[0]), .B(n_4), .CI(in_35[0]));
  ADDFX1 g3825(.CO(n_28), .S(n_29), .A(in_15[0]), .B(in_6[0]), .CI(in_21[0]));
  ADDFX1 g3826(.CO(n_26), .S(n_27), .A(n_15), .B(in_23[1]), .CI(n_11));
  ADDFX1 g3827(.CO(n_24), .S(n_25), .A(in_10[1]), .B(n_13), .CI(in_17[1]));
  ADDFX1 g3828(.CO(n_22), .S(n_23), .A(in_25[0]), .B(in_16[0]), .CI(in_32[0]));
  OAI21X1 g3829(.Y(n_21), .A0(in_36[2]), .A1(in_24[0]), .B0(n_18));
  XOR2XL g3830(.Y(n_20), .A(in_7[1]), .B(in_30[1]));
  NOR2X1 g3831(.Y(n_19), .A(in_30[1]), .B(in_7[1]));
  NAND2X1 g3832(.Y(n_18), .A(in_36[2]), .B(in_24[0]));
  INVX1 g3833(.Y(n_17), .A(in_39[1]));
  INVX1 g3834(.Y(n_16), .A(in_0[0]));
  INVX1 g3835(.Y(n_15), .A(in_5[1]));
  INVX1 g3836(.Y(n_14), .A(in_11[1]));
  INVX1 g3837(.Y(n_13), .A(in_8[1]));
  INVX1 g3838(.Y(n_12), .A(in_4[1]));
  INVX1 g3839(.Y(n_11), .A(in_12[1]));
  INVX1 g3840(.Y(n_10), .A(in_1[0]));
  INVX1 g3841(.Y(n_9), .A(in_32[0]));
  INVX1 g3842(.Y(n_8), .A(in_18[1]));
  INVX1 g3843(.Y(n_7), .A(in_33[0]));
  INVX1 g3844(.Y(n_6), .A(in_38[1]));
  INVX1 g3845(.Y(n_5), .A(in_34[1]));
  INVX1 g3846(.Y(n_4), .A(in_29[0]));
  INVX1 g3847(.Y(n_3), .A(in_9[1]));
  INVX1 g3848(.Y(n_2), .A(in_22[1]));
  INVX1 g3849(.Y(n_1), .A(in_28[0]));
endmodule

module WALLACE_CSA_DUMMY_OP61_group_359287(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, out_0);
input  in_3, in_4, in_21, in_32;
input   [4:0] in_0;
input   [5:0] in_1;
input   [5:0] in_2;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [1:0] in_9;
input   [4:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [1:0] in_20;
input   [1:0] in_22;
input   [4:0] in_23;
input   [2:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [1:0] in_30;
input   [1:0] in_31;
input   [4:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [2:0] in_40;
input   [2:0] in_41;
input   [4:0] in_42;
input   [3:0] in_43;
input   [4:0] in_44;
output  [9:0] out_0;
wire  n_120, n_118, n_116, n_115, n_114, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_84, n_83, 
    n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, 
    n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, 
    n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, 
    n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, 
    n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, 
    n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_32, in_21, in_4, 
    in_3;
wire   [9:0] out_0;
wire   [3:0] in_43;
wire   [2:0] in_41;
wire   [2:0] in_40;
wire   [2:0] in_24;
wire   [1:0] in_34;
wire   [1:0] in_31;
wire   [1:0] in_30;
wire   [1:0] in_29;
wire   [1:0] in_22;
wire   [1:0] in_20;
wire   [1:0] in_9;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_2;
wire   [5:0] in_1;
wire   [4:0] in_44;
wire   [4:0] in_42;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_23;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_10;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1386(.Y(out_0[9]), .A(n_120));
  ADDFX1 g1387(.CO(n_120), .S(out_0[5]), .A(n_83), .B(n_110), .CI(n_118));
  ADDFX1 g1388(.CO(n_118), .S(out_0[4]), .A(n_111), .B(n_114), .CI(n_116));
  ADDFX1 g1389(.CO(n_116), .S(out_0[3]), .A(n_108), .B(n_112), .CI(n_115));
  ADDFX1 g1390(.CO(n_114), .S(n_115), .A(n_92), .B(n_102), .CI(n_107));
  ADDFX1 g1391(.CO(n_112), .S(out_0[2]), .A(n_96), .B(n_104), .CI(n_109));
  ADDFX1 g1392(.CO(n_110), .S(n_111), .A(n_77), .B(n_100), .CI(n_106));
  ADDFX1 g1393(.CO(n_108), .S(n_109), .A(n_93), .B(n_99), .CI(n_103));
  ADDFX1 g1394(.CO(n_106), .S(n_107), .A(n_90), .B(n_98), .CI(n_101));
  ADDFX1 g1395(.CO(n_104), .S(out_0[1]), .A(n_84), .B(n_97), .CI(n_95));
  ADDFX1 g1396(.CO(n_102), .S(n_103), .A(n_91), .B(n_88), .CI(n_94));
  ADDFX1 g1397(.CO(n_100), .S(n_101), .A(n_69), .B(n_80), .CI(n_86));
  ADDFX1 g1398(.CO(n_98), .S(n_99), .A(n_67), .B(n_81), .CI(n_87));
  ADDFX1 g1399(.CO(n_96), .S(n_97), .A(n_71), .B(n_79), .CI(n_89));
  ADDFX1 g1400(.CO(n_94), .S(n_95), .A(n_63), .B(n_58), .CI(n_82));
  ADDFX1 g1401(.CO(n_92), .S(n_93), .A(n_70), .B(n_57), .CI(n_78));
  ADDFX1 g1402(.CO(n_90), .S(n_91), .A(n_39), .B(n_59), .CI(n_73));
  ADDFX1 g1403(.CO(n_88), .S(n_89), .A(n_60), .B(n_74), .CI(n_65));
  ADDFX1 g1404(.CO(n_86), .S(n_87), .A(n_31), .B(n_61), .CI(n_75));
  ADDFX1 g1405(.CO(n_84), .S(out_0[0]), .A(n_66), .B(n_64), .CI(n_72));
  INVX1 g1406(.Y(n_83), .A(n_77));
  ADDFX1 g1407(.CO(n_81), .S(n_82), .A(n_45), .B(n_32), .CI(n_62));
  OAI2BB1X1 g1408(.Y(n_80), .A0N(n_56), .A1N(n_76), .B0(n_83));
  ADDFX1 g1409(.CO(n_78), .S(n_79), .A(n_42), .B(n_53), .CI(n_68));
  NOR2X1 g1411(.Y(n_77), .A(n_56), .B(n_76));
  ADDFX1 g1412(.CO(n_76), .S(n_75), .A(n_8), .B(in_43[2]), .CI(n_55));
  ADDFX1 g1413(.CO(n_73), .S(n_74), .A(n_49), .B(n_35), .CI(n_37));
  ADDFX1 g1414(.CO(n_71), .S(n_72), .A(n_44), .B(n_38), .CI(n_54));
  ADDFX1 g1415(.CO(n_69), .S(n_70), .A(n_41), .B(n_25), .CI(n_23));
  ADDFX1 g1416(.CO(n_67), .S(n_68), .A(n_33), .B(n_29), .CI(n_43));
  ADDFX1 g1417(.CO(n_65), .S(n_66), .A(n_36), .B(n_30), .CI(n_46));
  ADDFX1 g1418(.CO(n_63), .S(n_64), .A(n_34), .B(n_28), .CI(n_52));
  ADDFX1 g1419(.CO(n_61), .S(n_62), .A(in_31[1]), .B(n_9), .CI(n_22));
  ADDFX1 g1420(.CO(n_59), .S(n_60), .A(n_4), .B(n_27), .CI(n_51));
  ADDFX1 g1421(.CO(n_57), .S(n_58), .A(n_26), .B(n_24), .CI(n_40));
  ADDHX1 g1422(.CO(n_56), .S(n_55), .A(n_19), .B(n_21));
  ADDFX1 g1423(.CO(n_53), .S(n_54), .A(in_13[0]), .B(in_6[0]), .CI(n_50));
  ADDFX1 g1424(.CO(n_51), .S(n_52), .A(in_7[0]), .B(n_1), .CI(n_6));
  INVX1 g1425(.Y(n_50), .A(n_48));
  INVX1 g1426(.Y(n_49), .A(n_47));
  ADDFX1 g1427(.CO(n_47), .S(n_48), .A(in_11[0]), .B(in_5[0]), .CI(in_18[0]));
  ADDFX1 g1428(.CO(n_45), .S(n_46), .A(in_4), .B(n_12), .CI(n_18));
  ADDFX1 g1429(.CO(n_43), .S(n_44), .A(in_9[0]), .B(n_10), .CI(in_22[0]));
  ADDFX1 g1430(.CO(n_41), .S(n_42), .A(in_1[1]), .B(n_11), .CI(in_41[0]));
  ADDFX1 g1431(.CO(n_39), .S(n_40), .A(in_24[1]), .B(n_7), .CI(in_13[1]));
  ADDFX1 g1432(.CO(n_37), .S(n_38), .A(n_14), .B(in_1[0]), .CI(n_15));
  ADDFX1 g1433(.CO(n_35), .S(n_36), .A(in_3), .B(in_12[0]), .CI(in_20[0]));
  ADDFX1 g1434(.CO(n_33), .S(n_34), .A(in_21), .B(n_2), .CI(in_32));
  ADDFX1 g1435(.CO(n_31), .S(n_32), .A(in_29[1]), .B(in_30[1]), .CI(n_13));
  ADDFX1 g1436(.CO(n_29), .S(n_30), .A(in_2[0]), .B(in_34[0]), .CI(in_41[0]));
  ADDFX1 g1437(.CO(n_27), .S(n_28), .A(in_15[0]), .B(in_17[0]), .CI(n_16));
  ADDFX1 g1438(.CO(n_25), .S(n_26), .A(in_22[0]), .B(in_40[1]), .CI(n_17));
  ADDFX1 g1439(.CO(n_23), .S(n_24), .A(in_2[0]), .B(n_3), .CI(n_5));
  XNOR2X1 g1440(.Y(n_22), .A(in_8[1]), .B(n_20));
  NAND2X1 g1441(.Y(n_21), .A(in_8[1]), .B(n_20));
  XNOR2X1 g1442(.Y(n_20), .A(in_14[1]), .B(in_16[1]));
  NOR2XL g1443(.Y(n_19), .A(in_14[1]), .B(in_16[1]));
  INVX1 g1444(.Y(n_18), .A(in_42[0]));
  INVX1 g1445(.Y(n_17), .A(in_44[1]));
  INVX1 g1446(.Y(n_16), .A(in_27[0]));
  INVX1 g1447(.Y(n_15), .A(in_36[0]));
  INVX1 g1448(.Y(n_14), .A(in_19[0]));
  INVX1 g1449(.Y(n_13), .A(in_10[1]));
  INVX1 g1450(.Y(n_12), .A(in_25[0]));
  INVX1 g1451(.Y(n_11), .A(in_28[1]));
  INVX1 g1452(.Y(n_10), .A(in_0[0]));
  INVX1 g1453(.Y(n_9), .A(in_26[1]));
  INVX1 g1454(.Y(n_8), .A(in_17[0]));
  INVX1 g1455(.Y(n_7), .A(in_33[1]));
  INVX1 g1456(.Y(n_6), .A(in_38[0]));
  INVX1 g1457(.Y(n_5), .A(in_39[1]));
  INVX1 g1458(.Y(n_4), .A(in_6[1]));
  INVX1 g1459(.Y(n_3), .A(in_35[1]));
  INVX1 g1460(.Y(n_2), .A(in_23[0]));
  INVX1 g1461(.Y(n_1), .A(in_37[0]));
endmodule

module WALLACE_CSA_DUMMY_OP62_group_359293(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88, out_0);
input  in_5, in_49, in_67, in_68, in_85;
input   [4:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [1:0] in_4;
input   [4:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [1:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
input   [1:0] in_41;
input   [4:0] in_42;
input   [1:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [2:0] in_48;
input   [1:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [1:0] in_53;
input   [4:0] in_54;
input   [2:0] in_55;
input   [4:0] in_56;
input   [1:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [1:0] in_60;
input   [1:0] in_61;
input   [1:0] in_62;
input   [4:0] in_63;
input   [1:0] in_64;
input   [1:0] in_65;
input   [4:0] in_66;
input   [1:0] in_69;
input   [4:0] in_70;
input   [4:0] in_71;
input   [4:0] in_72;
input   [4:0] in_73;
input   [4:0] in_74;
input   [4:0] in_75;
input   [4:0] in_76;
input   [4:0] in_77;
input   [4:0] in_78;
input   [4:0] in_79;
input   [4:0] in_80;
input   [4:0] in_81;
input   [4:0] in_82;
input   [4:0] in_83;
input   [1:0] in_84;
input   [1:0] in_86;
input   [4:0] in_87;
input   [4:0] in_88;
output  [9:0] out_0;
wire  n_274, n_272, n_270, n_268, n_266, n_264, n_263, n_262, n_261, n_260, 
    n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, 
    n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
    n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, 
    n_218, n_217, n_216, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
    n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, 
    n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, 
    n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, 
    n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, 
    n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_85, 
    in_68, in_67, in_49, in_5;
wire   [9:0] out_0;
wire   [2:0] in_55;
wire   [2:0] in_48;
wire   [2:0] in_37;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [1:0] in_86;
wire   [1:0] in_84;
wire   [1:0] in_69;
wire   [1:0] in_65;
wire   [1:0] in_64;
wire   [1:0] in_62;
wire   [1:0] in_61;
wire   [1:0] in_60;
wire   [1:0] in_57;
wire   [1:0] in_53;
wire   [1:0] in_51;
wire   [1:0] in_50;
wire   [1:0] in_45;
wire   [1:0] in_43;
wire   [1:0] in_41;
wire   [1:0] in_40;
wire   [1:0] in_34;
wire   [1:0] in_10;
wire   [1:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_88;
wire   [4:0] in_87;
wire   [4:0] in_83;
wire   [4:0] in_82;
wire   [4:0] in_81;
wire   [4:0] in_80;
wire   [4:0] in_79;
wire   [4:0] in_78;
wire   [4:0] in_77;
wire   [4:0] in_76;
wire   [4:0] in_75;
wire   [4:0] in_74;
wire   [4:0] in_73;
wire   [4:0] in_72;
wire   [4:0] in_71;
wire   [4:0] in_70;
wire   [4:0] in_66;
wire   [4:0] in_63;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_56;
wire   [4:0] in_54;
wire   [4:0] in_52;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_44;
wire   [4:0] in_42;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_6;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g8854(.Y(out_0[9]), .A(n_274));
  ADDFX1 g8855(.CO(n_274), .S(out_0[7]), .A(n_228), .B(n_256), .CI(n_272));
  ADDFX1 g8856(.CO(n_272), .S(out_0[6]), .A(n_257), .B(n_260), .CI(n_270));
  ADDFX1 g8857(.CO(n_270), .S(out_0[5]), .A(n_262), .B(n_261), .CI(n_268));
  ADDFX1 g8858(.CO(n_268), .S(out_0[4]), .A(n_258), .B(n_263), .CI(n_266));
  ADDFX1 g8859(.CO(n_266), .S(out_0[3]), .A(n_251), .B(n_259), .CI(n_264));
  ADDFX1 g8860(.CO(n_264), .S(out_0[2]), .A(n_235), .B(n_248), .CI(n_253));
  ADDFX1 g8861(.CO(n_262), .S(n_263), .A(n_242), .B(n_250), .CI(n_255));
  ADDFX1 g8862(.CO(n_260), .S(n_261), .A(n_244), .B(n_247), .CI(n_254));
  ADDFX1 g8863(.CO(n_258), .S(n_259), .A(n_237), .B(n_243), .CI(n_252));
  ADDFX1 g8864(.CO(n_256), .S(n_257), .A(n_222), .B(n_229), .CI(n_246));
  ADDFX1 g8865(.CO(n_254), .S(n_255), .A(n_230), .B(n_236), .CI(n_245));
  ADDFX1 g8866(.CO(n_252), .S(n_253), .A(n_225), .B(n_238), .CI(n_241));
  ADDFX1 g8867(.CO(n_250), .S(n_251), .A(n_231), .B(n_234), .CI(n_240));
  ADDFX1 g8868(.CO(n_248), .S(out_0[1]), .A(n_214), .B(n_207), .CI(n_239));
  ADDFX1 g8869(.CO(n_246), .S(n_247), .A(n_232), .B(n_200), .CI(n_223));
  ADDFX1 g8870(.CO(n_244), .S(n_245), .A(n_233), .B(n_202), .CI(n_201));
  ADDFX1 g8871(.CO(n_242), .S(n_243), .A(n_218), .B(n_224), .CI(n_203));
  ADDFX1 g8872(.CO(n_240), .S(n_241), .A(n_208), .B(n_211), .CI(n_221));
  ADDFX1 g8873(.CO(n_238), .S(n_239), .A(n_209), .B(n_217), .CI(n_186));
  ADDFX1 g8874(.CO(n_236), .S(n_237), .A(n_199), .B(n_210), .CI(n_220));
  ADDFX1 g8875(.CO(n_234), .S(n_235), .A(n_219), .B(n_216), .CI(n_206));
  ADDFX1 g8876(.CO(n_232), .S(n_233), .A(n_195), .B(n_204), .CI(n_198));
  ADDFX1 g8877(.CO(n_230), .S(n_231), .A(n_205), .B(n_179), .CI(n_212));
  INVX1 g8878(.Y(n_229), .A(n_227));
  INVX1 g8879(.Y(n_228), .A(n_226));
  ADDFX1 g8880(.CO(n_226), .S(n_227), .A(n_0), .B(in_3[6]), .CI(in_2[6]));
  ADDFX1 g8881(.CO(n_224), .S(n_225), .A(n_213), .B(n_187), .CI(n_185));
  ADDFX1 g8882(.CO(n_222), .S(n_223), .A(n_197), .B(in_3[5]), .CI(in_2[5]));
  ADDFX1 g8883(.CO(n_220), .S(n_221), .A(n_194), .B(n_173), .CI(in_2[2]));
  ADDFX1 g8884(.CO(n_218), .S(n_219), .A(n_168), .B(n_184), .CI(n_180));
  ADDFX1 g8885(.CO(n_216), .S(n_217), .A(n_190), .B(n_171), .CI(n_163));
  ADDFX1 g8886(.CO(n_214), .S(out_0[0]), .A(n_172), .B(n_192), .CI(n_164));
  ADDFX1 g8887(.CO(n_212), .S(n_213), .A(n_161), .B(n_181), .CI(n_170));
  ADDFX1 g8888(.CO(n_210), .S(n_211), .A(n_177), .B(n_189), .CI(in_3[2]));
  ADDFX1 g8889(.CO(n_208), .S(n_209), .A(n_162), .B(n_174), .CI(n_182));
  ADDFX1 g8890(.CO(n_206), .S(n_207), .A(n_178), .B(n_191), .CI(n_188));
  ADDFX1 g8891(.CO(n_204), .S(n_205), .A(n_131), .B(n_193), .CI(n_169));
  ADDFX1 g8892(.CO(n_202), .S(n_203), .A(n_183), .B(n_176), .CI(in_2[3]));
  ADDFX1 g8893(.CO(n_200), .S(n_201), .A(n_175), .B(in_3[4]), .CI(in_2[4]));
  ADDFX1 g8894(.CO(n_198), .S(n_199), .A(n_166), .B(n_167), .CI(in_3[3]));
  XNOR2X1 g8895(.Y(n_197), .A(n_78), .B(n_196));
  ADDFX1 g8897(.CO(n_196), .S(n_195), .A(n_78), .B(n_121), .CI(n_165));
  ADDFX1 g8898(.CO(n_193), .S(n_194), .A(n_151), .B(n_147), .CI(n_145));
  ADDFX1 g8899(.CO(n_191), .S(n_192), .A(n_158), .B(n_114), .CI(n_140));
  ADDFX1 g8900(.CO(n_189), .S(n_190), .A(n_155), .B(n_157), .CI(n_146));
  ADDFX1 g8901(.CO(n_187), .S(n_188), .A(n_154), .B(n_128), .CI(in_2[1]));
  ADDFX1 g8902(.CO(n_185), .S(n_186), .A(n_139), .B(n_130), .CI(in_3[1]));
  ADDFX1 g8903(.CO(n_183), .S(n_184), .A(n_144), .B(n_160), .CI(n_153));
  ADDFX1 g8904(.CO(n_181), .S(n_182), .A(n_152), .B(n_111), .CI(n_113));
  ADDFX1 g8905(.CO(n_179), .S(n_180), .A(n_129), .B(n_150), .CI(n_132));
  ADDFX1 g8906(.CO(n_177), .S(n_178), .A(n_125), .B(n_116), .CI(n_141));
  ADDFX1 g8907(.CO(n_175), .S(n_176), .A(n_143), .B(n_122), .CI(n_149));
  ADDFX1 g8908(.CO(n_173), .S(n_174), .A(n_134), .B(n_148), .CI(n_118));
  ADDFX1 g8909(.CO(n_171), .S(n_172), .A(n_142), .B(n_126), .CI(n_112));
  ADDFX1 g8910(.CO(n_169), .S(n_170), .A(n_115), .B(n_117), .CI(n_133));
  ADDFX1 g8911(.CO(n_167), .S(n_168), .A(n_123), .B(n_138), .CI(n_127));
  ADDFX1 g8912(.CO(n_165), .S(n_166), .A(n_78), .B(n_159), .CI(n_137));
  ADDFX1 g8913(.CO(n_163), .S(n_164), .A(n_156), .B(in_2[0]), .CI(in_3[0]));
  ADDFX1 g8914(.CO(n_161), .S(n_162), .A(n_108), .B(n_109), .CI(n_124));
  ADDFX1 g8915(.CO(n_159), .S(n_160), .A(n_69), .B(n_92), .CI(n_63));
  ADDFX1 g8916(.CO(n_157), .S(n_158), .A(n_91), .B(n_37), .CI(n_83));
  ADDFX1 g8917(.CO(n_155), .S(n_156), .A(n_68), .B(n_103), .CI(n_101));
  ADDFX1 g8918(.CO(n_153), .S(n_154), .A(n_70), .B(n_97), .CI(n_93));
  ADDFX1 g8919(.CO(n_151), .S(n_152), .A(n_90), .B(n_56), .CI(n_61));
  INVX1 g8920(.Y(n_150), .A(n_136));
  INVX1 g8921(.Y(n_149), .A(n_135));
  ADDFX1 g8922(.CO(n_147), .S(n_148), .A(n_44), .B(n_80), .CI(n_100));
  ADDFX1 g8923(.CO(n_145), .S(n_146), .A(in_31[1]), .B(n_42), .CI(n_102));
  ADDFX1 g8924(.CO(n_143), .S(n_144), .A(n_96), .B(n_98), .CI(n_84));
  ADDFX1 g8925(.CO(n_141), .S(n_142), .A(n_62), .B(n_43), .CI(n_66));
  ADDFX1 g8926(.CO(n_139), .S(n_140), .A(n_55), .B(n_72), .CI(n_110));
  ADDFX1 g8927(.CO(n_137), .S(n_138), .A(in_48[0]), .B(n_104), .CI(n_38));
  ADDFX1 g8928(.CO(n_135), .S(n_136), .A(n_35), .B(n_51), .CI(n_94));
  ADDFX1 g8929(.CO(n_133), .S(n_134), .A(n_40), .B(n_86), .CI(n_75));
  ADDFX1 g8930(.CO(n_131), .S(n_132), .A(n_79), .B(n_77), .CI(n_107));
  ADDFX1 g8931(.CO(n_129), .S(n_130), .A(n_39), .B(n_71), .CI(n_106));
  ADDFX1 g8932(.CO(n_127), .S(n_128), .A(n_64), .B(n_105), .CI(n_99));
  ADDFX1 g8933(.CO(n_125), .S(n_126), .A(n_47), .B(n_76), .CI(n_41));
  ADDFX1 g8934(.CO(n_123), .S(n_124), .A(n_46), .B(n_67), .CI(n_85));
  INVX1 g8935(.Y(n_122), .A(n_120));
  INVX1 g8936(.Y(n_121), .A(n_119));
  ADDFX1 g8937(.CO(n_119), .S(n_120), .A(n_33), .B(n_50), .CI(n_48));
  ADDFX1 g8938(.CO(n_117), .S(n_118), .A(n_82), .B(n_65), .CI(n_52));
  ADDFX1 g8939(.CO(n_115), .S(n_116), .A(n_54), .B(n_36), .CI(n_59));
  ADDFX1 g8940(.CO(n_113), .S(n_114), .A(n_81), .B(n_87), .CI(n_57));
  ADDFX1 g8941(.CO(n_111), .S(n_112), .A(n_60), .B(n_53), .CI(n_45));
  ADDFX1 g8942(.CO(n_109), .S(n_110), .A(in_32[0]), .B(n_34), .CI(in_25[0]));
  ADDFX1 g8943(.CO(n_107), .S(n_108), .A(n_15), .B(n_32), .CI(in_19[1]));
  INVX1 g8944(.Y(n_106), .A(n_95));
  INVX1 g8945(.Y(n_105), .A(n_89));
  INVX1 g8946(.Y(n_104), .A(n_88));
  ADDFX1 g8947(.CO(n_102), .S(n_103), .A(in_23[0]), .B(n_5), .CI(in_84[0]));
  ADDFX1 g8948(.CO(n_100), .S(n_101), .A(in_29[0]), .B(n_31), .CI(n_21));
  ADDFX1 g8949(.CO(n_98), .S(n_99), .A(in_37[1]), .B(n_22), .CI(in_62[1]));
  ADDFX1 g8950(.CO(n_96), .S(n_97), .A(in_61[1]), .B(n_13), .CI(n_4));
  ADDFX1 g8951(.CO(n_94), .S(n_95), .A(in_32[1]), .B(in_25[1]), .CI(in_20[1]));
  ADDFX1 g8952(.CO(n_92), .S(n_93), .A(in_4[1]), .B(n_25), .CI(n_7));
  ADDFX1 g8953(.CO(n_90), .S(n_91), .A(in_12[0]), .B(in_22[0]), .CI(in_31[0]));
  ADDFX1 g8954(.CO(n_88), .S(n_89), .A(in_30[1]), .B(in_44[1]), .CI(in_82[1]));
  ADDFX1 g8955(.CO(n_86), .S(n_87), .A(in_19[0]), .B(in_51[0]), .CI(in_53[0]));
  ADDFX1 g8956(.CO(n_84), .S(n_85), .A(in_55[1]), .B(n_28), .CI(n_17));
  ADDFX1 g8957(.CO(n_82), .S(n_83), .A(in_57[0]), .B(in_34[0]), .CI(in_65[0]));
  INVX1 g8958(.Y(n_81), .A(n_74));
  INVX1 g8959(.Y(n_80), .A(n_73));
  INVX1 g8960(.Y(n_79), .A(n_58));
  INVX1 g8962(.Y(n_77), .A(n_49));
  ADDFX1 g8963(.CO(n_75), .S(n_76), .A(in_64[0]), .B(n_6), .CI(n_27));
  ADDFX1 g8964(.CO(n_73), .S(n_74), .A(in_17[0]), .B(in_33[0]), .CI(in_63[0]));
  ADDFX1 g8965(.CO(n_71), .S(n_72), .A(in_50[0]), .B(in_74[0]), .CI(in_20[0]));
  ADDFX1 g8966(.CO(n_69), .S(n_70), .A(in_21[1]), .B(in_84[0]), .CI(n_10));
  ADDFX1 g8967(.CO(n_67), .S(n_68), .A(n_20), .B(in_40[0]), .CI(n_12));
  ADDFX1 g8968(.CO(n_65), .S(n_66), .A(in_5), .B(n_18), .CI(in_66[0]));
  ADDFX1 g8969(.CO(n_63), .S(n_64), .A(in_50[0]), .B(n_3), .CI(n_29));
  ADDFX1 g8970(.CO(n_61), .S(n_62), .A(in_59[0]), .B(in_49), .CI(n_26));
  ADDFX1 g8971(.CO(n_59), .S(n_60), .A(in_43[0]), .B(n_1), .CI(n_30));
  ADDFX1 g8972(.CO(n_78), .S(n_58), .A(in_27[0]), .B(in_74[0]), .CI(in_75[0]));
  ADDFX1 g8973(.CO(n_56), .S(n_57), .A(in_24[0]), .B(n_24), .CI(in_58[0]));
  ADDFX1 g8974(.CO(n_54), .S(n_55), .A(in_67), .B(in_48[0]), .CI(in_68));
  ADDFX1 g8975(.CO(n_52), .S(n_53), .A(in_27[0]), .B(n_8), .CI(in_69[0]));
  ADDFX1 g8976(.CO(n_50), .S(n_51), .A(in_47[0]), .B(in_58[0]), .CI(in_59[0]));
  ADDFX1 g8977(.CO(n_48), .S(n_49), .A(in_66[0]), .B(in_31[2]), .CI(in_19[2]));
  ADDFX1 g8978(.CO(n_46), .S(n_47), .A(in_9[0]), .B(in_85), .CI(n_9));
  ADDFX1 g8979(.CO(n_44), .S(n_45), .A(in_41[0]), .B(n_19), .CI(in_45[0]));
  ADDFX1 g8980(.CO(n_42), .S(n_43), .A(in_75[0]), .B(in_10[0]), .CI(n_11));
  ADDFX1 g8981(.CO(n_40), .S(n_41), .A(in_15[0]), .B(in_6[0]), .CI(in_47[0]));
  ADDFX1 g8982(.CO(n_38), .S(n_39), .A(in_16[1]), .B(n_2), .CI(n_14));
  ADDFX1 g8983(.CO(n_36), .S(n_37), .A(in_60[0]), .B(n_23), .CI(in_86[0]));
  AOI21X1 g8984(.Y(n_35), .A0(in_26[2]), .A1(n_16), .B0(n_33));
  XOR2XL g8985(.Y(n_34), .A(in_72[0]), .B(in_0[0]));
  NOR2X1 g8986(.Y(n_33), .A(in_26[2]), .B(n_16));
  NOR2X1 g8987(.Y(n_32), .A(in_72[0]), .B(in_0[0]));
  INVX1 g8988(.Y(n_31), .A(in_52[0]));
  INVX1 g8989(.Y(n_30), .A(in_46[0]));
  INVX1 g8990(.Y(n_29), .A(in_83[1]));
  INVX1 g8991(.Y(n_28), .A(in_78[1]));
  INVX1 g8992(.Y(n_27), .A(in_79[0]));
  INVX1 g8993(.Y(n_26), .A(in_77[0]));
  INVX1 g8994(.Y(n_25), .A(in_38[1]));
  INVX1 g8995(.Y(n_24), .A(in_13[0]));
  INVX1 g8996(.Y(n_23), .A(in_35[0]));
  INVX1 g8997(.Y(n_22), .A(in_1[1]));
  INVX1 g8998(.Y(n_21), .A(in_8[0]));
  INVX1 g8999(.Y(n_20), .A(in_76[0]));
  INVX1 g9000(.Y(n_19), .A(in_7[0]));
  INVX1 g9001(.Y(n_18), .A(in_14[0]));
  INVX1 g9002(.Y(n_17), .A(in_56[1]));
  INVX1 g9003(.Y(n_16), .A(in_6[0]));
  INVX1 g9004(.Y(n_15), .A(in_48[0]));
  INVX1 g9005(.Y(n_14), .A(in_88[1]));
  INVX1 g9006(.Y(n_13), .A(in_73[1]));
  INVX1 g9007(.Y(n_12), .A(in_80[0]));
  INVX1 g9008(.Y(n_11), .A(in_81[0]));
  INVX1 g9009(.Y(n_10), .A(in_87[1]));
  INVX1 g9010(.Y(n_9), .A(in_36[0]));
  INVX1 g9011(.Y(n_8), .A(in_39[0]));
  INVX1 g9012(.Y(n_7), .A(in_11[1]));
  INVX1 g9013(.Y(n_6), .A(in_28[0]));
  INVX1 g9014(.Y(n_5), .A(in_18[0]));
  INVX1 g9015(.Y(n_4), .A(in_54[1]));
  INVX1 g9016(.Y(n_3), .A(in_71[1]));
  INVX1 g9017(.Y(n_2), .A(in_70[1]));
  INVX1 g9018(.Y(n_1), .A(in_42[0]));
  NAND2BX1 g2(.Y(n_0), .AN(n_78), .B(n_196));
endmodule

module WALLACE_CSA_DUMMY_OP70_group_106217(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, out_0);
input  in_32, in_33, in_34, in_62, in_64;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [9:0] in_4;
input   [9:0] in_5;
input   [8:0] in_6;
input   [6:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [1:0] in_30;
input   [4:0] in_31;
input   [1:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [2:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [1:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [3:0] in_51;
input   [1:0] in_52;
input   [4:0] in_53;
input   [1:0] in_54;
input   [1:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [1:0] in_63;
input   [4:0] in_65;
input   [4:0] in_66;
input   [1:0] in_67;
input   [4:0] in_68;
input   [4:0] in_69;
input   [4:0] in_70;
input   [4:0] in_71;
input   [4:0] in_72;
input   [4:0] in_73;
input   [4:0] in_74;
input   [4:0] in_75;
input   [4:0] in_76;
input   [4:0] in_77;
input   [4:0] in_78;
input   [1:0] in_79;
input   [3:0] in_80;
input   [4:0] in_81;
output  [9:0] out_0;
wire  n_300, n_298, n_296, n_294, n_292, n_290, n_289, n_288, n_287, n_286, 
    n_284, n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, 
    n_274, n_273, n_272, n_271, n_270, n_268, n_267, n_266, n_265, n_264, 
    n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
    n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, 
    n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, 
    n_223, n_222, n_221, n_219, n_218, n_217, n_216, n_215, n_214, n_213, 
    n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, 
    n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, 
    n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
    n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, 
    n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
    n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, 
    n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
    n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
    n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, 
    n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, 
    n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1, n_0, in_64, in_62, in_34, in_33, in_32;
wire   [9:0] out_0;
wire   [3:0] in_80;
wire   [3:0] in_51;
wire   [1:0] in_79;
wire   [1:0] in_67;
wire   [1:0] in_63;
wire   [1:0] in_61;
wire   [1:0] in_55;
wire   [1:0] in_54;
wire   [1:0] in_52;
wire   [1:0] in_46;
wire   [1:0] in_45;
wire   [1:0] in_35;
wire   [1:0] in_30;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_7;
wire   [8:0] in_6;
wire   [9:0] in_5;
wire   [9:0] in_4;
wire   [4:0] in_81;
wire   [4:0] in_78;
wire   [4:0] in_77;
wire   [4:0] in_76;
wire   [4:0] in_75;
wire   [4:0] in_74;
wire   [4:0] in_73;
wire   [4:0] in_72;
wire   [4:0] in_71;
wire   [4:0] in_70;
wire   [4:0] in_69;
wire   [4:0] in_68;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_60;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_53;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_41;
wire   [2:0] in_0;
  INVX1 g9592(.Y(out_0[9]), .A(n_300));
  ADDFX1 g9593(.CO(n_300), .S(out_0[8]), .A(n_47), .B(n_274), .CI(n_298));
  ADDFX1 g9594(.CO(n_298), .S(out_0[7]), .A(n_275), .B(n_282), .CI(n_296));
  ADDFX1 g9595(.CO(n_296), .S(out_0[6]), .A(n_288), .B(n_283), .CI(n_294));
  ADDFX1 g9596(.CO(n_294), .S(out_0[5]), .A(n_286), .B(n_289), .CI(n_292));
  ADDFX1 g9597(.CO(n_292), .S(out_0[4]), .A(n_280), .B(n_287), .CI(n_290));
  ADDFX1 g9598(.CO(n_290), .S(out_0[3]), .A(n_272), .B(n_281), .CI(n_284));
  ADDFX1 g9599(.CO(n_288), .S(n_289), .A(n_270), .B(n_276), .CI(n_279));
  ADDFX1 g9600(.CO(n_286), .S(n_287), .A(n_271), .B(n_266), .CI(n_277));
  ADDFX1 g9601(.CO(n_284), .S(out_0[2]), .A(n_247), .B(n_268), .CI(n_273));
  ADDFX1 g9602(.CO(n_282), .S(n_283), .A(n_260), .B(n_278), .CI(n_263));
  ADDFX1 g9603(.CO(n_280), .S(n_281), .A(n_246), .B(n_267), .CI(n_265));
  ADDFX1 g9604(.CO(n_278), .S(n_279), .A(n_245), .B(n_261), .CI(n_258));
  ADDFX1 g9605(.CO(n_276), .S(n_277), .A(n_256), .B(n_264), .CI(n_259));
  ADDFX1 g9606(.CO(n_274), .S(n_275), .A(n_216), .B(n_43), .CI(n_262));
  ADDFX1 g9607(.CO(n_272), .S(n_273), .A(n_255), .B(n_252), .CI(n_243));
  ADDFX1 g9608(.CO(n_270), .S(n_271), .A(n_248), .B(n_251), .CI(n_239));
  ADDFX1 g9609(.CO(n_268), .S(out_0[1]), .A(n_219), .B(n_213), .CI(n_253));
  ADDFX1 g9610(.CO(n_266), .S(n_267), .A(n_249), .B(n_242), .CI(n_257));
  ADDFX1 g9611(.CO(n_264), .S(n_265), .A(n_241), .B(n_254), .CI(n_228));
  ADDFX1 g9612(.CO(n_262), .S(n_263), .A(n_229), .B(in_5[6]), .CI(n_244));
  ADDFX1 g9613(.CO(n_260), .S(n_261), .A(n_210), .B(n_250), .CI(n_238));
  ADDFX1 g9614(.CO(n_258), .S(n_259), .A(n_240), .B(in_5[4]), .CI(n_227));
  ADDFX1 g9615(.CO(n_256), .S(n_257), .A(n_218), .B(n_234), .CI(n_236));
  ADDFX1 g9616(.CO(n_254), .S(n_255), .A(n_226), .B(n_233), .CI(n_212));
  ADDFX1 g9617(.CO(n_252), .S(n_253), .A(n_231), .B(n_195), .CI(n_224));
  ADDFX1 g9618(.CO(n_250), .S(n_251), .A(n_221), .B(n_215), .CI(n_217));
  ADDFX1 g9619(.CO(n_248), .S(n_249), .A(n_222), .B(n_225), .CI(n_232));
  ADDFX1 g9620(.CO(n_246), .S(n_247), .A(n_230), .B(n_235), .CI(n_237));
  ADDFX1 g9621(.CO(n_244), .S(n_245), .A(n_214), .B(in_4[5]), .CI(in_5[5]));
  ADDFX1 g9622(.CO(n_242), .S(n_243), .A(n_194), .B(in_5[2]), .CI(n_223));
  ADDFX1 g9623(.CO(n_240), .S(n_241), .A(n_185), .B(n_205), .CI(n_208));
  ADDFX1 g9624(.CO(n_238), .S(n_239), .A(n_204), .B(n_187), .CI(in_4[4]));
  ADDFX1 g9625(.CO(n_236), .S(n_237), .A(n_201), .B(n_188), .CI(in_4[2]));
  ADDFX1 g9626(.CO(n_234), .S(n_235), .A(n_191), .B(n_203), .CI(n_209));
  ADDFX1 g9627(.CO(n_232), .S(n_233), .A(n_183), .B(n_206), .CI(n_176));
  ADDFX1 g9628(.CO(n_230), .S(n_231), .A(n_207), .B(n_189), .CI(n_192));
  OAI2BB1X1 g9629(.Y(n_229), .A0N(n_211), .A1N(in_4[6]), .B0(n_216));
  ADDFX1 g9630(.CO(n_227), .S(n_228), .A(n_202), .B(in_4[3]), .CI(in_5[3]));
  ADDFX1 g9631(.CO(n_225), .S(n_226), .A(n_179), .B(n_196), .CI(n_198));
  ADDFX1 g9632(.CO(n_223), .S(n_224), .A(n_199), .B(n_180), .CI(in_5[1]));
  ADDFX1 g9633(.CO(n_221), .S(n_222), .A(n_182), .B(n_173), .CI(n_200));
  ADDFX1 g9634(.CO(n_219), .S(out_0[0]), .A(n_181), .B(n_175), .CI(n_193));
  ADDFX1 g9635(.CO(n_217), .S(n_218), .A(n_178), .B(n_190), .CI(in_6[3]));
  OR2X1 g9636(.Y(n_216), .A(n_211), .B(in_4[6]));
  ADDFX1 g9637(.CO(n_214), .S(n_215), .A(n_172), .B(n_184), .CI(in_6[4]));
  ADDFX1 g9638(.CO(n_212), .S(n_213), .A(n_197), .B(n_174), .CI(n_177));
  ADDFX1 g9639(.CO(n_211), .S(n_210), .A(n_124), .B(n_186), .CI(n_26));
  ADDFX1 g9640(.CO(n_208), .S(n_209), .A(n_163), .B(n_141), .CI(in_6[2]));
  ADDFX1 g9641(.CO(n_206), .S(n_207), .A(n_168), .B(n_131), .CI(n_170));
  ADDFX1 g9642(.CO(n_204), .S(n_205), .A(n_162), .B(n_147), .CI(n_140));
  ADDFX1 g9643(.CO(n_202), .S(n_203), .A(n_149), .B(n_136), .CI(n_158));
  ADDFX1 g9644(.CO(n_200), .S(n_201), .A(n_156), .B(n_166), .CI(n_116));
  ADDFX1 g9645(.CO(n_198), .S(n_199), .A(n_126), .B(n_154), .CI(n_164));
  ADDFX1 g9646(.CO(n_196), .S(n_197), .A(n_167), .B(n_151), .CI(n_142));
  ADDFX1 g9647(.CO(n_194), .S(n_195), .A(n_161), .B(n_159), .CI(in_4[1]));
  ADDFX1 g9648(.CO(n_192), .S(n_193), .A(n_143), .B(n_171), .CI(in_4[0]));
  ADDFX1 g9649(.CO(n_190), .S(n_191), .A(n_139), .B(n_153), .CI(n_160));
  ADDFX1 g9650(.CO(n_188), .S(n_189), .A(n_157), .B(n_137), .CI(n_145));
  ADDFX1 g9651(.CO(n_186), .S(n_187), .A(n_128), .B(n_127), .CI(n_146));
  ADDFX1 g9652(.CO(n_184), .S(n_185), .A(n_138), .B(n_152), .CI(n_129));
  ADDFX1 g9653(.CO(n_182), .S(n_183), .A(n_99), .B(n_134), .CI(n_150));
  ADDFX1 g9654(.CO(n_180), .S(n_181), .A(n_133), .B(n_155), .CI(n_165));
  ADDFX1 g9655(.CO(n_178), .S(n_179), .A(n_125), .B(n_130), .CI(n_144));
  ADDFX1 g9656(.CO(n_176), .S(n_177), .A(n_135), .B(n_132), .CI(in_6[1]));
  ADDFX1 g9657(.CO(n_174), .S(n_175), .A(n_52), .B(n_169), .CI(in_5[0]));
  ADDFX1 g9658(.CO(n_172), .S(n_173), .A(n_48), .B(n_148), .CI(n_115));
  ADDFX1 g9659(.CO(n_170), .S(n_171), .A(n_78), .B(n_94), .CI(n_58));
  ADDFX1 g9660(.CO(n_168), .S(n_169), .A(in_9[0]), .B(n_98), .CI(n_62));
  ADDFX1 g9661(.CO(n_166), .S(n_167), .A(n_77), .B(n_107), .CI(n_119));
  ADDFX1 g9662(.CO(n_164), .S(n_165), .A(n_108), .B(n_64), .CI(in_6[0]));
  ADDFX1 g9663(.CO(n_162), .S(n_163), .A(n_111), .B(n_102), .CI(n_118));
  ADDFX1 g9664(.CO(n_160), .S(n_161), .A(n_88), .B(n_112), .CI(n_76));
  ADDFX1 g9665(.CO(n_158), .S(n_159), .A(n_66), .B(n_100), .CI(n_51));
  ADDFX1 g9666(.CO(n_156), .S(n_157), .A(n_73), .B(n_109), .CI(n_97));
  ADDFX1 g9667(.CO(n_154), .S(n_155), .A(n_54), .B(n_96), .CI(n_74));
  ADDFX1 g9668(.CO(n_152), .S(n_153), .A(n_83), .B(n_79), .CI(n_105));
  ADDFX1 g9669(.CO(n_150), .S(n_151), .A(n_63), .B(n_95), .CI(n_93));
  ADDFX1 g9670(.CO(n_148), .S(n_149), .A(n_65), .B(n_55), .CI(n_59));
  ADDFX1 g9671(.CO(n_146), .S(n_147), .A(n_117), .B(n_101), .CI(n_69));
  ADDFX1 g9672(.CO(n_144), .S(n_145), .A(n_80), .B(n_84), .CI(n_106));
  ADDFX1 g9673(.CO(n_142), .S(n_143), .A(n_86), .B(n_90), .CI(n_120));
  ADDFX1 g9674(.CO(n_140), .S(n_141), .A(n_122), .B(n_67), .CI(n_70));
  ADDFX1 g9675(.CO(n_138), .S(n_139), .A(n_45), .B(n_75), .CI(n_87));
  ADDFX1 g9676(.CO(n_136), .S(n_137), .A(n_56), .B(n_60), .CI(n_68));
  ADDFX1 g9677(.CO(n_134), .S(n_135), .A(n_85), .B(n_57), .CI(n_61));
  ADDFX1 g9678(.CO(n_132), .S(n_133), .A(n_110), .B(n_72), .CI(n_50));
  ADDFX1 g9679(.CO(n_130), .S(n_131), .A(n_89), .B(n_53), .CI(n_49));
  ADDFX1 g9680(.CO(n_128), .S(n_129), .A(n_39), .B(n_0), .CI(n_121));
  OAI2BB1X1 g9681(.Y(n_127), .A0N(n_41), .A1N(n_123), .B0(n_124));
  ADDFX1 g9682(.CO(n_125), .S(n_126), .A(in_7[1]), .B(in_19[1]), .CI(n_71));
  OR2X1 g9683(.Y(n_124), .A(n_41), .B(n_123));
  OAI21X1 g9684(.Y(n_123), .A0(in_12[3]), .A1(n_46), .B0(n_42));
  INVX1 g9685(.Y(n_122), .A(n_114));
  INVX1 g9686(.Y(n_121), .A(n_113));
  INVX1 g9687(.Y(n_120), .A(n_104));
  INVX1 g9688(.Y(n_119), .A(n_103));
  INVX1 g9689(.Y(n_118), .A(n_92));
  INVX1 g9690(.Y(n_117), .A(n_91));
  ADDFX1 g9691(.CO(n_115), .S(n_116), .A(n_40), .B(n_6), .CI(in_12[2]));
  ADDFX1 g9692(.CO(n_113), .S(n_114), .A(in_42[0]), .B(in_71[0]), .CI(in_28[0]));
  ADDFX1 g9693(.CO(n_111), .S(n_112), .A(in_61[1]), .B(n_31), .CI(in_63[1]));
  ADDFX1 g9694(.CO(n_109), .S(n_110), .A(in_67[0]), .B(n_38), .CI(n_22));
  ADDFX1 g9695(.CO(n_107), .S(n_108), .A(in_25[0]), .B(in_42[0]), .CI(n_17));
  ADDFX1 g9696(.CO(n_105), .S(n_106), .A(in_46[1]), .B(n_13), .CI(in_73[0]));
  ADDFX1 g9697(.CO(n_103), .S(n_104), .A(in_1[0]), .B(in_22[0]), .CI(in_47[0]));
  ADDFX1 g9698(.CO(n_101), .S(n_102), .A(n_19), .B(in_80[2]), .CI(n_20));
  ADDFX1 g9699(.CO(n_99), .S(n_100), .A(in_26[1]), .B(n_27), .CI(n_44));
  ADDFX1 g9700(.CO(n_97), .S(n_98), .A(in_11[0]), .B(n_32), .CI(n_18));
  ADDFX1 g9701(.CO(n_95), .S(n_96), .A(in_19[0]), .B(in_53[0]), .CI(n_36));
  ADDFX1 g9702(.CO(n_93), .S(n_94), .A(in_12[0]), .B(in_2[0]), .CI(in_59[0]));
  ADDFX1 g9703(.CO(n_91), .S(n_92), .A(in_18[0]), .B(in_2[0]), .CI(in_36[0]));
  ADDFX1 g9704(.CO(n_89), .S(n_90), .A(in_28[0]), .B(n_34), .CI(n_12));
  ADDFX1 g9705(.CO(n_87), .S(n_88), .A(in_12[1]), .B(n_23), .CI(n_35));
  ADDFX1 g9706(.CO(n_85), .S(n_86), .A(n_9), .B(n_28), .CI(in_34));
  INVX1 g9707(.Y(n_84), .A(n_82));
  INVX1 g9708(.Y(n_83), .A(n_81));
  ADDFX1 g9709(.CO(n_81), .S(n_82), .A(in_57[1]), .B(in_39[1]), .CI(in_81[1]));
  ADDFX1 g9710(.CO(n_79), .S(n_80), .A(in_21[1]), .B(in_55[1]), .CI(n_15));
  ADDFX1 g9711(.CO(n_77), .S(n_78), .A(in_18[0]), .B(in_52[0]), .CI(in_62));
  ADDFX1 g9712(.CO(n_75), .S(n_76), .A(n_21), .B(n_10), .CI(in_77[0]));
  ADDFX1 g9713(.CO(n_73), .S(n_74), .A(in_23[0]), .B(in_64), .CI(n_11));
  ADDFX1 g9714(.CO(n_71), .S(n_72), .A(in_16[0]), .B(n_24), .CI(n_33));
  ADDFX1 g9715(.CO(n_69), .S(n_70), .A(in_51[2]), .B(n_2), .CI(n_25));
  ADDFX1 g9716(.CO(n_67), .S(n_68), .A(in_0[1]), .B(in_59[0]), .CI(n_8));
  ADDFX1 g9717(.CO(n_65), .S(n_66), .A(in_54[1]), .B(in_41[0]), .CI(n_37));
  ADDFX1 g9718(.CO(n_63), .S(n_64), .A(in_32), .B(n_4), .CI(in_41[0]));
  ADDFX1 g9719(.CO(n_61), .S(n_62), .A(n_3), .B(n_5), .CI(in_77[0]));
  ADDFX1 g9720(.CO(n_59), .S(n_60), .A(in_35[1]), .B(n_14), .CI(n_30));
  ADDFX1 g9721(.CO(n_57), .S(n_58), .A(in_71[0]), .B(in_73[0]), .CI(in_79[0]));
  ADDFX1 g9722(.CO(n_55), .S(n_56), .A(in_45[1]), .B(n_29), .CI(n_16));
  ADDFX1 g9723(.CO(n_53), .S(n_54), .A(in_24[0]), .B(in_30[0]), .CI(n_7));
  ADDFX1 g9724(.CO(n_51), .S(n_52), .A(in_58[0]), .B(in_26[0]), .CI(in_14[0]));
  ADDFX1 g9725(.CO(n_49), .S(n_50), .A(in_33), .B(in_15[0]), .CI(in_36[0]));
  XOR2XL g9726(.Y(n_48), .A(in_12[3]), .B(n_46));
  NOR2X1 g9727(.Y(n_47), .A(in_5[7]), .B(n_43));
  OAI2BB1X1 g9728(.Y(n_46), .A0N(in_73[0]), .A1N(in_77[0]), .B0(n_42));
  XNOR2X1 g9729(.Y(n_45), .A(in_8[2]), .B(in_16[0]));
  XNOR2X1 g9730(.Y(n_44), .A(in_58[0]), .B(in_3[1]));
  CLKXOR2X1 g9732(.Y(n_43), .A(in_4[6]), .B(in_5[7]));
  OR2XL g9733(.Y(n_42), .A(in_73[0]), .B(in_77[0]));
  NOR2XL g9734(.Y(n_41), .A(in_58[0]), .B(in_59[0]));
  NOR2X1 g9735(.Y(n_40), .A(in_3[1]), .B(n_1));
  NOR2BX1 g9736(.Y(n_39), .AN(in_8[2]), .B(in_16[0]));
  INVX1 g9737(.Y(n_38), .A(in_72[0]));
  INVX1 g9738(.Y(n_37), .A(in_65[1]));
  INVX1 g9739(.Y(n_36), .A(in_68[0]));
  INVX1 g9740(.Y(n_35), .A(in_56[1]));
  INVX1 g9741(.Y(n_34), .A(in_60[0]));
  INVX1 g9742(.Y(n_33), .A(in_74[0]));
  INVX1 g9743(.Y(n_32), .A(in_44[0]));
  INVX1 g9744(.Y(n_31), .A(in_29[1]));
  INVX1 g9745(.Y(n_30), .A(in_43[1]));
  INVX1 g9746(.Y(n_29), .A(in_24[1]));
  INVX1 g9747(.Y(n_28), .A(in_27[0]));
  INVX1 g9748(.Y(n_27), .A(in_9[1]));
  INVX1 g9749(.Y(n_26), .A(in_6[5]));
  INVX1 g9750(.Y(n_25), .A(in_19[2]));
  INVX1 g9751(.Y(n_24), .A(in_40[0]));
  INVX1 g9752(.Y(n_23), .A(in_25[1]));
  INVX1 g9753(.Y(n_22), .A(in_70[0]));
  INVX1 g9754(.Y(n_21), .A(in_50[1]));
  INVX1 g9755(.Y(n_20), .A(in_53[0]));
  INVX1 g9756(.Y(n_19), .A(in_23[0]));
  INVX1 g9758(.Y(n_18), .A(in_75[0]));
  INVX1 g9759(.Y(n_17), .A(in_76[0]));
  INVX1 g9760(.Y(n_16), .A(in_49[1]));
  INVX1 g9761(.Y(n_15), .A(in_66[1]));
  INVX1 g9762(.Y(n_14), .A(in_78[1]));
  INVX1 g9763(.Y(n_13), .A(in_48[1]));
  INVX1 g9764(.Y(n_12), .A(in_20[0]));
  INVX1 g9765(.Y(n_11), .A(in_10[0]));
  INVX1 g9766(.Y(n_10), .A(in_69[1]));
  INVX1 g9767(.Y(n_9), .A(in_13[0]));
  INVX1 g9768(.Y(n_8), .A(in_14[1]));
  INVX1 g9769(.Y(n_7), .A(in_17[0]));
  INVX1 g9770(.Y(n_6), .A(in_26[2]));
  INVX1 g9771(.Y(n_5), .A(in_38[0]));
  INVX1 g9772(.Y(n_4), .A(in_37[0]));
  INVX1 g9773(.Y(n_3), .A(in_31[0]));
  INVX1 g9774(.Y(n_2), .A(in_7[2]));
  INVX1 g9775(.Y(n_1), .A(in_58[0]));
  MXI2XL g2(.Y(n_0), .A(n_1), .B(in_58[0]), .S0(in_59[0]));
endmodule

module WALLACE_CSA_DUMMY_OP74_group_109823(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, out_0);
input  in_37, in_38;
input   [2:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [1:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [4:0] in_27;
input   [2:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [2:0] in_33;
input   [4:0] in_34;
input   [1:0] in_35;
input   [4:0] in_36;
input   [4:0] in_39;
input   [1:0] in_40;
output  [9:0] out_0;
wire  n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_35, n_33, 
    n_31, n_29, n_27, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, in_38, in_37;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_35;
wire   [1:0] in_26;
wire   [1:0] in_24;
wire   [1:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_39;
wire   [4:0] in_36;
wire   [4:0] in_34;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_25;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_1;
wire   [2:0] in_33;
wire   [2:0] in_32;
wire   [2:0] in_30;
wire   [2:0] in_28;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  ADDFX1 cdnfadd_000_1(.CO(n_113), .S(n_112), .A(n_20), .B(n_2), .CI(in_21[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_111), .S(n_110), .A(in_37), .B(n_4), .CI(in_8[0]));
  ADDFX1 cdnfadd_000_3(.CO(n_109), .S(n_108), .A(in_17[0]), .B(in_24[0]), .CI(
    n_9));
  ADDFX1 cdnfadd_000_4(.CO(n_107), .S(n_106), .A(in_26[0]), .B(n_8), .CI(
    in_40[0]));
  ADDFX1 cdnfadd_000_5(.CO(n_105), .S(n_104), .A(n_15), .B(in_15[0]), .CI(n_16));
  ADDFX1 cdnfadd_000_6(.CO(n_103), .S(n_102), .A(n_19), .B(in_10[0]), .CI(
    in_35[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_101), .S(n_100), .A(n_3), .B(in_30[0]), .CI(
    in_20[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_99), .S(n_98), .A(in_38), .B(in_19[0]), .CI(in_5[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_97), .S(n_96), .A(in_7[0]), .B(in_3[0]), .CI(
    in_14[0]));
  ADDFX1 cdnfadd_000_10(.CO(n_83), .S(n_82), .A(n_110), .B(n_108), .CI(n_106));
  ADDFX1 cdnfadd_000_11(.CO(n_81), .S(n_114), .A(n_100), .B(n_104), .CI(n_112));
  ADDFX1 cdnfadd_000_12(.CO(n_80), .S(n_122), .A(n_23), .B(n_102), .CI(n_96));
  ADDFX1 cdnfadd_000_13(.CO(n_63), .S(n_115), .A(n_98), .B(in_2[0]), .CI(n_82));
  ADDFX1 cdnfadd_001_0(.CO(n_95), .S(n_94), .A(in_0[1]), .B(in_12[1]), .CI(
    in_11[1]));
  ADDFX1 cdnfadd_001_1(.CO(n_93), .S(n_92), .A(n_6), .B(in_32[1]), .CI(n_10));
  ADDFX1 cdnfadd_001_2(.CO(n_91), .S(n_90), .A(in_28[1]), .B(n_14), .CI(in_33[1]));
  ADDFX1 cdnfadd_001_3(.CO(n_89), .S(n_88), .A(n_21), .B(in_7[1]), .CI(n_7));
  ADDFX1 cdnfadd_001_4(.CO(n_87), .S(n_86), .A(n_17), .B(n_1), .CI(in_9[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_79), .S(n_78), .A(n_11), .B(in_18[1]), .CI(n_103));
  ADDFX1 cdnfadd_001_6(.CO(n_77), .S(n_76), .A(n_109), .B(n_113), .CI(n_101));
  ADDFX1 cdnfadd_001_7(.CO(n_75), .S(n_74), .A(n_22), .B(n_111), .CI(n_107));
  ADDFX1 cdnfadd_001_8(.CO(n_73), .S(n_72), .A(n_105), .B(n_94), .CI(n_90));
  ADDFX1 cdnfadd_001_9(.CO(n_71), .S(n_70), .A(n_92), .B(n_99), .CI(n_86));
  ADDFX1 cdnfadd_001_10(.CO(n_65), .S(n_64), .A(n_88), .B(n_97), .CI(n_78));
  ADDFX1 cdnfadd_001_11(.CO(n_62), .S(n_61), .A(n_76), .B(n_74), .CI(n_81));
  ADDFX1 cdnfadd_001_12(.CO(n_60), .S(n_59), .A(n_83), .B(n_72), .CI(n_80));
  ADDFX1 cdnfadd_001_13(.CO(n_46), .S(n_123), .A(n_64), .B(n_70), .CI(in_2[1]));
  ADDFX1 cdnfadd_001_14(.CO(n_43), .S(n_116), .A(n_61), .B(n_63), .CI(n_59));
  ADDFX1 cdnfadd_002_0(.CO(n_85), .S(n_84), .A(n_13), .B(n_18), .CI(n_5));
  ADDFX1 cdnfadd_002_1(.CO(n_69), .S(n_68), .A(in_30[0]), .B(n_91), .CI(n_95));
  ADDFX1 cdnfadd_002_2(.CO(n_67), .S(n_66), .A(n_93), .B(n_89), .CI(n_84));
  ADDFX1 cdnfadd_002_3(.CO(n_58), .S(n_57), .A(n_87), .B(n_79), .CI(n_77));
  ADDFX1 cdnfadd_002_4(.CO(n_56), .S(n_55), .A(n_75), .B(n_68), .CI(n_73));
  ADDFX1 cdnfadd_002_5(.CO(n_45), .S(n_44), .A(n_66), .B(n_71), .CI(n_65));
  ADDFX1 cdnfadd_002_6(.CO(n_52), .S(n_51), .A(n_62), .B(n_57), .CI(n_55));
  ADDFX1 cdnfadd_002_7(.CO(n_42), .S(n_124), .A(in_2[2]), .B(n_44), .CI(n_60));
  ADDFX1 cdnfadd_002_8(.CO(n_125), .S(n_117), .A(n_46), .B(n_51), .CI(n_43));
  ADDFX1 cdnfadd_003_0(.CO(n_54), .S(n_53), .A(n_69), .B(n_24), .CI(n_67));
  ADDFX1 cdnfadd_003_1(.CO(n_50), .S(n_49), .A(n_58), .B(n_56), .CI(n_53));
  ADDFX1 cdnfadd_003_2(.CO(n_41), .S(n_40), .A(n_45), .B(in_2[3]), .CI(n_52));
  ADDFX1 cdnfadd_003_3(.CO(n_126), .S(n_118), .A(n_49), .B(n_42), .CI(n_40));
  ADDFX1 cdnfadd_004_0(.CO(n_48), .S(n_47), .A(n_24), .B(n_54), .CI(in_2[4]));
  ADDFX1 cdnfadd_004_1(.CO(n_120), .S(n_119), .A(n_50), .B(n_47), .CI(n_41));
  ADDFX1 cdnfadd_005_0(.CO(n_121), .S(n_127), .A(n_85), .B(in_2[5]), .CI(n_48));
  INVX1 g302(.Y(out_0[9]), .A(n_37));
  ADDFX1 g303(.CO(n_37), .S(out_0[6]), .A(n_12), .B(n_121), .CI(n_35));
  ADDFX1 g304(.CO(n_35), .S(out_0[5]), .A(n_127), .B(n_120), .CI(n_33));
  ADDFX1 g305(.CO(n_33), .S(out_0[4]), .A(n_126), .B(n_119), .CI(n_31));
  ADDFX1 g306(.CO(n_31), .S(out_0[3]), .A(n_125), .B(n_29), .CI(n_118));
  ADDFX1 g307(.CO(n_29), .S(out_0[2]), .A(n_27), .B(n_117), .CI(n_124));
  ADDFX1 g308(.CO(n_27), .S(out_0[1]), .A(n_25), .B(n_116), .CI(n_123));
  ADDFX1 g309(.CO(n_25), .S(out_0[0]), .A(n_114), .B(n_122), .CI(n_115));
  INVX1 g310(.Y(n_24), .A(n_85));
  OAI21X1 g311(.Y(n_23), .A0(in_39[0]), .A1(in_22[0]), .B0(n_22));
  NAND2X1 g312(.Y(n_22), .A(in_39[0]), .B(in_22[0]));
  INVX1 g313(.Y(n_21), .A(in_19[1]));
  INVX1 g314(.Y(n_20), .A(in_25[0]));
  INVX1 g315(.Y(n_19), .A(in_34[0]));
  INVX1 g316(.Y(n_18), .A(in_9[2]));
  INVX1 g317(.Y(n_17), .A(in_5[1]));
  INVX1 g318(.Y(n_16), .A(in_27[0]));
  INVX1 g319(.Y(n_15), .A(in_6[0]));
  INVX1 g320(.Y(n_14), .A(in_36[1]));
  INVX1 g321(.Y(n_13), .A(in_8[0]));
  INVX1 g322(.Y(n_12), .A(in_2[6]));
  INVX1 g323(.Y(n_11), .A(in_30[0]));
  INVX1 g324(.Y(n_10), .A(in_13[1]));
  INVX1 g325(.Y(n_9), .A(in_23[0]));
  INVX1 g326(.Y(n_8), .A(in_31[0]));
  INVX1 g327(.Y(n_7), .A(in_3[1]));
  INVX1 g328(.Y(n_6), .A(in_4[1]));
  INVX1 g329(.Y(n_5), .A(in_18[2]));
  INVX1 g330(.Y(n_4), .A(in_29[0]));
  INVX1 g331(.Y(n_3), .A(in_1[0]));
  INVX1 g332(.Y(n_2), .A(in_16[0]));
  INVX1 g333(.Y(n_1), .A(in_14[1]));
endmodule

module WALLACE_CSA_DUMMY_OP75_group_109813_6325(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, out_0);
input  in_37;
input   [4:0] in_0;
input   [6:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [4:0] in_6;
input   [4:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [2:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [1:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [1:0] in_38;
output  [9:0] out_0;
wire  n_123, n_121, n_119, n_117, n_116, n_115, n_113, n_112, n_111, n_110, 
    n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, 
    n_98, n_97, n_96, n_95, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_37;
wire   [9:0] out_0;
wire   [1:0] in_38;
wire   [1:0] in_33;
wire   [1:0] in_30;
wire   [1:0] in_29;
wire   [2:0] in_36;
wire   [2:0] in_25;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [6:0] in_1;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_7;
wire   [4:0] in_6;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1432(.Y(out_0[9]), .A(n_123));
  ADDFX1 g1433(.CO(n_123), .S(out_0[5]), .A(n_87), .B(n_109), .CI(n_121));
  ADDFX1 g1434(.CO(n_121), .S(out_0[4]), .A(n_110), .B(n_115), .CI(n_119));
  ADDFX1 g1435(.CO(n_119), .S(out_0[3]), .A(n_111), .B(n_116), .CI(n_117));
  ADDFX1 g1436(.CO(n_117), .S(out_0[2]), .A(n_108), .B(n_112), .CI(n_113));
  ADDFX1 g1437(.CO(n_115), .S(n_116), .A(n_101), .B(n_107), .CI(n_104));
  ADDFX1 g1438(.CO(n_113), .S(out_0[1]), .A(n_96), .B(n_93), .CI(n_106));
  ADDFX1 g1439(.CO(n_111), .S(n_112), .A(n_95), .B(n_102), .CI(n_105));
  ADDFX1 g1440(.CO(n_109), .S(n_110), .A(n_88), .B(n_91), .CI(n_103));
  ADDFX1 g1441(.CO(n_107), .S(n_108), .A(n_97), .B(n_99), .CI(n_90));
  ADDFX1 g1442(.CO(n_105), .S(n_106), .A(n_79), .B(n_98), .CI(n_100));
  ADDFX1 g1443(.CO(n_103), .S(n_104), .A(n_85), .B(n_89), .CI(n_92));
  ADDFX1 g1444(.CO(n_101), .S(n_102), .A(n_69), .B(n_66), .CI(n_86));
  ADDFX1 g1445(.CO(n_99), .S(n_100), .A(n_54), .B(n_74), .CI(n_76));
  ADDFX1 g1446(.CO(n_97), .S(n_98), .A(n_59), .B(n_63), .CI(n_81));
  ADDFX1 g1447(.CO(n_95), .S(n_96), .A(n_72), .B(n_62), .CI(n_70));
  ADDFX1 g1448(.CO(n_93), .S(out_0[0]), .A(n_82), .B(n_64), .CI(n_80));
  ADDFX1 g1449(.CO(n_91), .S(n_92), .A(n_67), .B(n_84), .CI(n_65));
  ADDFX1 g1450(.CO(n_89), .S(n_90), .A(n_71), .B(n_68), .CI(n_61));
  ADDHX1 g1451(.CO(n_87), .S(n_88), .A(n_16), .B(n_83));
  ADDFX1 g1452(.CO(n_85), .S(n_86), .A(n_73), .B(n_75), .CI(n_78));
  ADDFX1 g1453(.CO(n_83), .S(n_84), .A(n_20), .B(n_25), .CI(n_77));
  ADDFX1 g1454(.CO(n_81), .S(n_82), .A(n_48), .B(n_34), .CI(n_50));
  ADDFX1 g1455(.CO(n_79), .S(n_80), .A(n_60), .B(n_56), .CI(n_28));
  ADDFX1 g1456(.CO(n_77), .S(n_78), .A(n_17), .B(n_31), .CI(n_57));
  ADDFX1 g1457(.CO(n_75), .S(n_76), .A(n_49), .B(n_51), .CI(n_35));
  ADDFX1 g1458(.CO(n_73), .S(n_74), .A(n_33), .B(n_39), .CI(n_47));
  ADDFX1 g1459(.CO(n_71), .S(n_72), .A(n_19), .B(n_29), .CI(n_58));
  ADDFX1 g1460(.CO(n_69), .S(n_70), .A(n_27), .B(n_44), .CI(n_55));
  ADDFX1 g1461(.CO(n_67), .S(n_68), .A(n_18), .B(n_45), .CI(n_23));
  ADDFX1 g1462(.CO(n_65), .S(n_66), .A(n_43), .B(n_53), .CI(n_26));
  ADDFX1 g1463(.CO(n_63), .S(n_64), .A(n_36), .B(n_40), .CI(n_30));
  ADDFX1 g1464(.CO(n_61), .S(n_62), .A(n_32), .B(n_46), .CI(n_24));
  ADDFX1 g1465(.CO(n_59), .S(n_60), .A(in_34[0]), .B(in_11[0]), .CI(n_52));
  ADDFX1 g1466(.CO(n_57), .S(n_58), .A(n_3), .B(n_13), .CI(in_25[0]));
  ADDFX1 g1467(.CO(n_55), .S(n_56), .A(in_12[0]), .B(in_15[0]), .CI(in_19[0]));
  ADDFX1 g1468(.CO(n_53), .S(n_54), .A(n_1), .B(n_12), .CI(in_2[1]));
  ADDFX1 g1469(.CO(n_51), .S(n_52), .A(in_8[0]), .B(in_2[0]), .CI(n_14));
  ADDFX1 g1470(.CO(n_49), .S(n_50), .A(in_20[0]), .B(in_29[0]), .CI(n_9));
  INVX1 g1471(.Y(n_48), .A(n_42));
  INVX1 g1472(.Y(n_47), .A(n_41));
  INVX1 g1473(.Y(n_46), .A(n_38));
  INVX1 g1474(.Y(n_45), .A(n_37));
  INVX1 g1475(.Y(n_44), .A(n_22));
  INVX1 g1476(.Y(n_43), .A(n_21));
  ADDFX1 g1477(.CO(n_41), .S(n_42), .A(in_0[0]), .B(in_22[0]), .CI(in_28[0]));
  ADDFX1 g1478(.CO(n_39), .S(n_40), .A(n_2), .B(n_6), .CI(in_30[0]));
  ADDFX1 g1479(.CO(n_37), .S(n_38), .A(in_18[1]), .B(in_26[1]), .CI(in_35[1]));
  ADDFX1 g1480(.CO(n_35), .S(n_36), .A(in_16[0]), .B(in_21[0]), .CI(in_25[0]));
  ADDFX1 g1481(.CO(n_33), .S(n_34), .A(n_10), .B(in_37), .CI(n_4));
  ADDFX1 g1482(.CO(n_31), .S(n_32), .A(in_17[1]), .B(n_11), .CI(in_36[0]));
  ADDFX1 g1483(.CO(n_29), .S(n_30), .A(in_33[0]), .B(n_8), .CI(in_36[0]));
  ADDFX1 g1484(.CO(n_27), .S(n_28), .A(in_4[0]), .B(in_13[0]), .CI(in_5[0]));
  ADDFX1 g1485(.CO(n_25), .S(n_26), .A(in_19[2]), .B(n_7), .CI(n_5));
  ADDFX1 g1486(.CO(n_23), .S(n_24), .A(in_12[1]), .B(in_11[1]), .CI(in_19[1]));
  ADDFX1 g1487(.CO(n_21), .S(n_22), .A(in_5[1]), .B(in_4[1]), .CI(in_15[1]));
  INVX1 g1488(.Y(n_20), .A(n_16));
  OAI2BB1X1 g1489(.Y(n_19), .A0N(in_38[1]), .A1N(n_15), .B0(n_17));
  OAI21X1 g1490(.Y(n_18), .A0(in_31[2]), .A1(in_21[0]), .B0(n_16));
  OR2X1 g1491(.Y(n_17), .A(in_38[1]), .B(n_15));
  NAND2X1 g1492(.Y(n_16), .A(in_31[2]), .B(in_21[0]));
  INVX1 g1493(.Y(n_15), .A(in_1[1]));
  INVX1 g1494(.Y(n_14), .A(in_32[0]));
  INVX1 g1495(.Y(n_13), .A(in_14[1]));
  INVX1 g1496(.Y(n_12), .A(in_13[1]));
  INVX1 g1497(.Y(n_11), .A(in_7[1]));
  INVX1 g1498(.Y(n_10), .A(in_24[0]));
  INVX1 g1499(.Y(n_9), .A(in_23[0]));
  INVX1 g1500(.Y(n_8), .A(in_9[0]));
  INVX1 g1501(.Y(n_7), .A(in_12[2]));
  INVX1 g1502(.Y(n_6), .A(in_3[0]));
  INVX1 g1503(.Y(n_5), .A(in_2[2]));
  INVX1 g1504(.Y(n_4), .A(in_6[0]));
  INVX1 g1505(.Y(n_3), .A(in_10[1]));
  INVX1 g1506(.Y(n_2), .A(in_27[0]));
  INVX1 g1507(.Y(n_1), .A(in_34[0]));
endmodule

module WALLACE_CSA_DUMMY_OP75_group_109813(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, out_0);
input   [2:0] in_0;
input   [4:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [1:0] in_18;
input   [4:0] in_19;
input   [3:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [2:0] in_24;
input   [2:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [4:0] in_37;
input   [2:0] in_38;
output  [9:0] out_0;
wire  n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_43, n_41, n_39, n_37, n_35, n_34, n_33, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
    n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_1;
wire   [9:0] out_0;
wire   [3:0] in_20;
wire   [1:0] in_29;
wire   [1:0] in_27;
wire   [1:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_19;
wire   [4:0] in_1;
wire   [2:0] in_38;
wire   [2:0] in_36;
wire   [2:0] in_25;
wire   [2:0] in_24;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  ADDFX1 cdnfadd_000_1(.CO(n_115), .S(n_114), .A(in_6[0]), .B(n_17), .CI(n_2));
  ADDFX1 cdnfadd_000_2(.CO(n_113), .S(n_112), .A(in_9[0]), .B(n_6), .CI(in_11[0]));
  ADDFX1 cdnfadd_000_3(.CO(n_111), .S(n_110), .A(n_12), .B(in_27[0]), .CI(
    in_17[0]));
  ADDFX1 cdnfadd_000_4(.CO(n_109), .S(n_108), .A(n_11), .B(n_8), .CI(n_20));
  ADDFX1 cdnfadd_000_5(.CO(n_107), .S(n_106), .A(in_18[0]), .B(in_10[0]), .CI(
    in_29[0]));
  ADDFX1 cdnfadd_000_6(.CO(n_105), .S(n_104), .A(n_15), .B(in_12[0]), .CI(
    in_16[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_103), .S(n_102), .A(in_3[0]), .B(in_7[0]), .CI(
    in_5[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_85), .S(n_116), .A(in_15[0]), .B(n_26), .CI(n_114));
  ADDFX1 cdnfadd_000_9(.CO(n_84), .S(n_123), .A(n_106), .B(n_104), .CI(n_108));
  ADDFX1 cdnfadd_000_10(.CO(n_83), .S(n_117), .A(n_110), .B(n_112), .CI(n_102));
  ADDFX1 cdnfadd_001_0(.CO(n_101), .S(n_100), .A(n_5), .B(n_3), .CI(n_9));
  ADDFX1 cdnfadd_001_2(.CO(n_82), .S(n_81), .A(n_100), .B(n_27), .CI(in_36[1]));
  ADDFX1 cdnfadd_001_3(.CO(n_99), .S(n_98), .A(in_4[1]), .B(n_21), .CI(in_24[1]));
  ADDFX1 cdnfadd_001_4(.CO(n_97), .S(n_96), .A(in_0[1]), .B(in_25[1]), .CI(n_4));
  ADDFX1 cdnfadd_001_5(.CO(n_95), .S(n_94), .A(n_1), .B(n_18), .CI(n_14));
  ADDFX1 cdnfadd_001_6(.CO(n_93), .S(n_92), .A(in_38[1]), .B(in_6[1]), .CI(n_10));
  ADDFX1 cdnfadd_001_7(.CO(n_91), .S(n_90), .A(in_3[1]), .B(in_7[1]), .CI(n_16));
  ADDFX1 cdnfadd_001_8(.CO(n_89), .S(n_88), .A(in_9[1]), .B(in_16[1]), .CI(
    in_12[1]));
  ADDFX1 cdnfadd_001_9(.CO(n_80), .S(n_79), .A(n_24), .B(n_109), .CI(n_111));
  ADDFX1 cdnfadd_001_10(.CO(n_68), .S(n_67), .A(n_81), .B(n_113), .CI(n_105));
  ADDFX1 cdnfadd_001_11(.CO(n_78), .S(n_77), .A(n_107), .B(n_115), .CI(n_92));
  ADDFX1 cdnfadd_001_12(.CO(n_76), .S(n_75), .A(n_98), .B(n_94), .CI(n_96));
  ADDFX1 cdnfadd_001_13(.CO(n_74), .S(n_73), .A(n_103), .B(n_90), .CI(n_88));
  ADDFX1 cdnfadd_001_14(.CO(n_62), .S(n_61), .A(n_79), .B(n_85), .CI(n_77));
  ADDFX1 cdnfadd_001_15(.CO(n_57), .S(n_124), .A(n_67), .B(n_84), .CI(n_75));
  ADDFX1 cdnfadd_001_16(.CO(n_56), .S(n_118), .A(n_83), .B(n_73), .CI(n_61));
  ADDFX1 cdnfadd_002_0(.CO(n_69), .S(n_72), .A(n_101), .B(n_25), .CI(in_20[2]));
  ADDFX1 cdnfadd_002_1(.CO(n_87), .S(n_86), .A(n_7), .B(n_13), .CI(n_19));
  ADDFX1 cdnfadd_002_2(.CO(n_66), .S(n_65), .A(in_6[2]), .B(n_82), .CI(n_99));
  ADDFX1 cdnfadd_002_3(.CO(n_64), .S(n_63), .A(n_97), .B(n_72), .CI(n_95));
  ADDFX1 cdnfadd_002_4(.CO(n_71), .S(n_70), .A(n_93), .B(n_91), .CI(n_86));
  ADDFX1 cdnfadd_002_5(.CO(n_60), .S(n_59), .A(n_89), .B(n_68), .CI(n_80));
  ADDFX1 cdnfadd_002_6(.CO(n_55), .S(n_54), .A(n_76), .B(n_78), .CI(n_65));
  ADDFX1 cdnfadd_002_7(.CO(n_53), .S(n_52), .A(n_63), .B(n_70), .CI(n_74));
  ADDFX1 cdnfadd_002_8(.CO(n_50), .S(n_125), .A(n_62), .B(n_59), .CI(n_57));
  ADDFX1 cdnfadd_002_9(.CO(n_126), .S(n_119), .A(n_54), .B(n_52), .CI(n_56));
  ADDFX1 cdnfadd_003_1(.CO(n_51), .S(n_58), .A(n_87), .B(n_30), .CI(n_66));
  ADDFX1 cdnfadd_003_2(.CO(n_47), .S(n_46), .A(n_64), .B(n_71), .CI(n_60));
  ADDFX1 cdnfadd_003_3(.CO(n_49), .S(n_48), .A(n_55), .B(n_58), .CI(n_53));
  ADDFX1 cdnfadd_003_4(.CO(n_127), .S(n_120), .A(n_46), .B(n_50), .CI(n_48));
  ADDFX1 cdnfadd_004_0(.CO(n_122), .S(n_121), .A(n_34), .B(n_47), .CI(n_49));
  INVX1 g294(.Y(out_0[9]), .A(n_43));
  ADDFX1 g295(.CO(n_43), .S(out_0[5]), .A(n_33), .B(n_122), .CI(n_41));
  ADDFX1 g296(.CO(n_41), .S(out_0[4]), .A(n_127), .B(n_121), .CI(n_39));
  ADDFX1 g297(.CO(n_39), .S(out_0[3]), .A(n_126), .B(n_37), .CI(n_120));
  ADDFX1 g298(.CO(n_37), .S(out_0[2]), .A(n_35), .B(n_125), .CI(n_119));
  ADDFX1 g299(.CO(n_35), .S(out_0[1]), .A(n_31), .B(n_124), .CI(n_118));
  ADDHX1 g300(.CO(n_33), .S(n_34), .A(n_29), .B(n_51));
  ADDFX1 g301(.CO(n_31), .S(out_0[0]), .A(n_116), .B(n_123), .CI(n_117));
  OAI21X1 g302(.Y(n_30), .A0(in_6[3]), .A1(n_28), .B0(n_29));
  NAND2X1 g303(.Y(n_29), .A(in_6[3]), .B(n_28));
  INVX1 g304(.Y(n_28), .A(n_69));
  OAI21X1 g305(.Y(n_27), .A0(in_11[1]), .A1(n_22), .B0(n_25));
  OAI21X1 g306(.Y(n_26), .A0(in_28[0]), .A1(n_23), .B0(n_24));
  NAND2X1 g307(.Y(n_25), .A(in_11[1]), .B(n_22));
  NAND2X1 g308(.Y(n_24), .A(in_28[0]), .B(n_23));
  XNOR2X1 g309(.Y(n_23), .A(in_13[0]), .B(in_2[0]));
  OR2XL g310(.Y(n_22), .A(in_13[0]), .B(in_2[0]));
  INVX1 g311(.Y(n_21), .A(in_35[1]));
  INVX1 g312(.Y(n_20), .A(in_1[0]));
  INVX1 g313(.Y(n_19), .A(in_16[2]));
  INVX1 g314(.Y(n_18), .A(in_19[1]));
  INVX1 g315(.Y(n_17), .A(in_31[0]));
  INVX1 g316(.Y(n_16), .A(in_5[1]));
  INVX1 g317(.Y(n_15), .A(in_32[0]));
  INVX1 g318(.Y(n_14), .A(in_37[1]));
  INVX1 g319(.Y(n_13), .A(in_9[2]));
  INVX1 g320(.Y(n_12), .A(in_23[0]));
  INVX1 g321(.Y(n_11), .A(in_33[0]));
  INVX1 g322(.Y(n_10), .A(in_15[1]));
  INVX1 g323(.Y(n_9), .A(in_10[1]));
  INVX1 g324(.Y(n_8), .A(in_34[0]));
  INVX1 g325(.Y(n_7), .A(in_12[2]));
  INVX1 g326(.Y(n_6), .A(in_22[0]));
  INVX1 g327(.Y(n_5), .A(in_14[1]));
  INVX1 g328(.Y(n_4), .A(in_26[1]));
  INVX1 g329(.Y(n_3), .A(in_8[1]));
  INVX1 g330(.Y(n_2), .A(in_21[0]));
  INVX1 g331(.Y(n_1), .A(in_30[1]));
endmodule

module WALLACE_CSA_DUMMY_OP78_group_359273(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, out_0);
input  in_20, in_21, in_23;
input   [4:0] in_0;
input   [1:0] in_1;
input   [1:0] in_2;
input   [7:0] in_3;
input   [5:0] in_4;
input   [4:0] in_5;
input   [4:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [1:0] in_22;
input   [4:0] in_24;
input   [2:0] in_25;
input   [2:0] in_26;
input   [4:0] in_27;
input   [1:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [2:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
output  [9:0] out_0;
wire  n_92, n_90, n_88, n_87, n_86, n_84, n_83, n_82, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_58, n_57, n_56, n_55, n_54, n_53, n_52, 
    n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_1, in_23, in_21, in_20;
wire   [9:0] out_0;
wire   [2:0] in_31;
wire   [2:0] in_26;
wire   [2:0] in_25;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_4;
wire   [7:0] in_3;
wire   [1:0] in_32;
wire   [1:0] in_28;
wire   [1:0] in_22;
wire   [1:0] in_2;
wire   [1:0] in_1;
wire   [4:0] in_33;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_24;
wire   [4:0] in_6;
wire   [4:0] in_5;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1130(.Y(out_0[9]), .A(n_92));
  ADDFX1 g1131(.CO(n_92), .S(out_0[5]), .A(n_46), .B(n_82), .CI(n_90));
  ADDFX1 g1132(.CO(n_90), .S(out_0[4]), .A(n_83), .B(n_86), .CI(n_88));
  ADDFX1 g1133(.CO(n_88), .S(out_0[3]), .A(n_78), .B(n_87), .CI(n_84));
  ADDFX1 g1134(.CO(n_86), .S(n_87), .A(n_68), .B(n_74), .CI(n_77));
  ADDFX1 g1135(.CO(n_84), .S(out_0[2]), .A(n_75), .B(n_79), .CI(n_80));
  ADDFX1 g1136(.CO(n_82), .S(n_83), .A(n_47), .B(n_70), .CI(n_76));
  ADDFX1 g1137(.CO(n_80), .S(out_0[1]), .A(n_61), .B(n_58), .CI(n_73));
  ADDFX1 g1138(.CO(n_78), .S(n_79), .A(n_52), .B(n_69), .CI(n_72));
  ADDFX1 g1139(.CO(n_76), .S(n_77), .A(n_5), .B(n_71), .CI(n_66));
  ADDFX1 g1140(.CO(n_74), .S(n_75), .A(n_60), .B(n_62), .CI(n_67));
  ADDFX1 g1141(.CO(n_72), .S(n_73), .A(n_37), .B(n_53), .CI(n_63));
  ADDFX1 g1142(.CO(n_70), .S(n_71), .A(n_47), .B(n_56), .CI(n_64));
  ADDFX1 g1143(.CO(n_68), .S(n_69), .A(n_35), .B(n_43), .CI(n_65));
  ADDFX1 g1144(.CO(n_66), .S(n_67), .A(n_50), .B(n_57), .CI(in_3[2]));
  ADDFX1 g1145(.CO(n_64), .S(n_65), .A(n_20), .B(n_12), .CI(n_48));
  ADDFX1 g1146(.CO(n_62), .S(n_63), .A(n_21), .B(n_14), .CI(n_49));
  ADDFX1 g1147(.CO(n_60), .S(n_61), .A(n_44), .B(n_41), .CI(n_51));
  ADDFX1 g1148(.CO(n_58), .S(out_0[0]), .A(n_40), .B(n_42), .CI(n_38));
  INVX1 g1149(.Y(n_57), .A(n_55));
  INVX1 g1150(.Y(n_56), .A(n_54));
  ADDFX1 g1151(.CO(n_54), .S(n_55), .A(in_5[0]), .B(in_30[0]), .CI(n_45));
  ADDFX1 g1152(.CO(n_52), .S(n_53), .A(n_36), .B(n_39), .CI(in_3[1]));
  ADDFX1 g1153(.CO(n_50), .S(n_51), .A(n_16), .B(n_22), .CI(n_33));
  ADDFX1 g1154(.CO(n_48), .S(n_49), .A(in_1[1]), .B(in_22[1]), .CI(n_32));
  INVX1 g1155(.Y(n_46), .A(n_47));
  ADDFX1 g1156(.CO(n_47), .S(n_45), .A(in_9[0]), .B(n_28), .CI(n_31));
  ADDFX1 g1157(.CO(n_43), .S(n_44), .A(n_26), .B(n_18), .CI(n_13));
  ADDFX1 g1158(.CO(n_41), .S(n_42), .A(in_13[0]), .B(n_17), .CI(n_34));
  ADDFX1 g1159(.CO(n_39), .S(n_40), .A(n_23), .B(n_27), .CI(n_19));
  ADDFX1 g1160(.CO(n_37), .S(n_38), .A(n_25), .B(n_15), .CI(in_3[0]));
  ADDFX1 g1161(.CO(n_35), .S(n_36), .A(n_4), .B(n_6), .CI(n_24));
  ADDFX1 g1162(.CO(n_33), .S(n_34), .A(in_19[0]), .B(in_28[0]), .CI(n_11));
  OAI21X1 g1163(.Y(n_32), .A0(n_10), .A1(n_29), .B0(n_30));
  INVX1 g1164(.Y(n_31), .A(n_30));
  NAND2X1 g1165(.Y(n_30), .A(n_10), .B(n_29));
  ADDFX1 g1166(.CO(n_28), .S(n_29), .A(in_7[1]), .B(in_15[1]), .CI(in_16[1]));
  ADDFX1 g1167(.CO(n_26), .S(n_27), .A(in_5[0]), .B(in_4[0]), .CI(n_8));
  ADDFX1 g1168(.CO(n_24), .S(n_25), .A(in_14[0]), .B(in_18[0]), .CI(in_30[0]));
  ADDFX1 g1169(.CO(n_22), .S(n_23), .A(in_2[0]), .B(in_32[0]), .CI(n_9));
  ADDFX1 g1170(.CO(n_20), .S(n_21), .A(in_11[1]), .B(n_2), .CI(in_25[1]));
  ADDFX1 g1171(.CO(n_18), .S(n_19), .A(in_10[0]), .B(in_17[0]), .CI(n_7));
  ADDFX1 g1172(.CO(n_16), .S(n_17), .A(in_21), .B(in_23), .CI(n_3));
  ADDFX1 g1173(.CO(n_14), .S(n_15), .A(n_1), .B(in_20), .CI(in_8[0]));
  ADDFX1 g1174(.CO(n_12), .S(n_13), .A(in_2[0]), .B(in_26[1]), .CI(in_31[1]));
  XNOR2X1 g1175(.Y(n_11), .A(in_12[0]), .B(in_9[0]));
  NAND2BX1 g1176(.Y(n_10), .AN(in_12[0]), .B(in_9[0]));
  INVX1 g1177(.Y(n_9), .A(in_33[0]));
  INVX1 g1178(.Y(n_8), .A(in_29[0]));
  INVX1 g1179(.Y(n_7), .A(in_24[0]));
  INVX1 g1180(.Y(n_6), .A(in_8[1]));
  INVX1 g1181(.Y(n_5), .A(in_3[3]));
  INVX1 g1182(.Y(n_4), .A(in_13[1]));
  INVX1 g1183(.Y(n_3), .A(in_27[0]));
  INVX1 g1184(.Y(n_2), .A(in_6[1]));
  INVX1 g1185(.Y(n_1), .A(in_0[0]));
endmodule

module WALLACE_CSA_DUMMY_OP82_group_359272(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, out_0);
input  in_9, in_10, in_15, in_16;
input   [4:0] in_0;
input   [2:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [2:0] in_6;
input   [2:0] in_7;
input   [4:0] in_8;
input   [4:0] in_11;
input   [2:0] in_12;
input   [4:0] in_13;
input   [1:0] in_14;
input   [2:0] in_17;
input   [2:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
output  [9:0] out_0;
wire  n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_21, n_18, n_16, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
    n_6, n_5, n_4, n_3, n_2, n_1, in_16, in_15, in_10, in_9;
wire   [9:0] out_0;
wire   [1:0] in_14;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [2:0] in_18;
wire   [2:0] in_17;
wire   [2:0] in_12;
wire   [2:0] in_7;
wire   [2:0] in_6;
wire   [2:0] in_1;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_13;
wire   [4:0] in_11;
wire   [4:0] in_8;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  assign out_0[5] = 1'b0;
  ADDFX1 cdnfadd_000_1(.CO(n_51), .S(n_52), .A(in_9), .B(n_6), .CI(in_7[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_50), .S(n_49), .A(in_16), .B(in_14[0]), .CI(n_4));
  ADDFX1 cdnfadd_000_3(.CO(n_48), .S(n_47), .A(in_15), .B(n_2), .CI(in_10));
  ADDFX1 cdnfadd_000_4(.CO(n_46), .S(n_45), .A(n_5), .B(n_9), .CI(in_6[0]));
  ADDFX1 cdnfadd_000_5(.CO(n_44), .S(n_58), .A(in_3[0]), .B(in_5[0]), .CI(n_13));
  ADDFX1 cdnfadd_000_6(.CO(n_37), .S(n_53), .A(n_49), .B(n_45), .CI(n_47));
  ADDFX1 cdnfadd_001_0(.CO(n_43), .S(n_42), .A(in_17[1]), .B(n_7), .CI(n_3));
  ADDFX1 cdnfadd_001_1(.CO(n_41), .S(n_40), .A(in_18[1]), .B(in_12[1]), .CI(
    in_1[1]));
  ADDFX1 cdnfadd_001_2(.CO(n_39), .S(n_38), .A(n_8), .B(in_7[0]), .CI(in_5[1]));
  ADDFX1 cdnfadd_001_3(.CO(n_36), .S(n_35), .A(in_3[1]), .B(n_12), .CI(n_46));
  ADDFX1 cdnfadd_001_4(.CO(n_34), .S(n_33), .A(n_51), .B(n_50), .CI(n_48));
  ADDFX1 cdnfadd_001_5(.CO(n_32), .S(n_31), .A(n_11), .B(n_38), .CI(n_42));
  ADDFX1 cdnfadd_001_6(.CO(n_28), .S(n_59), .A(n_40), .B(n_44), .CI(n_35));
  ADDFX1 cdnfadd_001_7(.CO(n_60), .S(n_54), .A(n_33), .B(n_37), .CI(n_31));
  ADDFX1 cdnfadd_002_0(.CO(n_30), .S(n_29), .A(n_1), .B(n_10), .CI(n_43));
  ADDFX1 cdnfadd_002_1(.CO(n_27), .S(n_26), .A(n_41), .B(n_39), .CI(n_36));
  ADDFX1 cdnfadd_002_2(.CO(n_25), .S(n_24), .A(n_29), .B(n_34), .CI(n_32));
  ADDFX1 cdnfadd_002_3(.CO(n_61), .S(n_55), .A(n_28), .B(n_26), .CI(n_24));
  ADDFX1 cdnfadd_003_0(.CO(n_57), .S(n_56), .A(n_30), .B(n_27), .CI(n_25));
  AO21XL g218(.Y(out_0[4]), .A0(n_57), .A1(n_21), .B0(out_0[9]));
  NOR2X1 g219(.Y(out_0[9]), .A(n_57), .B(n_21));
  ADDFX1 g220(.CO(n_21), .S(out_0[3]), .A(n_56), .B(n_61), .CI(n_18));
  ADDFX1 g221(.CO(n_18), .S(out_0[2]), .A(n_60), .B(n_16), .CI(n_55));
  ADDFX1 g222(.CO(n_16), .S(out_0[1]), .A(n_14), .B(n_59), .CI(n_54));
  ADDFX1 g223(.CO(n_14), .S(out_0[0]), .A(n_52), .B(n_58), .CI(n_53));
  OAI2BB1X1 g224(.Y(n_13), .A0N(in_4[0]), .A1N(in_2[0]), .B0(n_11));
  AOI2BB1X1 g225(.Y(n_12), .A0N(in_6[0]), .A1N(in_4[0]), .B0(n_10));
  OR2X1 g226(.Y(n_11), .A(in_4[0]), .B(in_2[0]));
  AND2X1 g227(.Y(n_10), .A(in_6[0]), .B(in_4[0]));
  INVX1 g228(.Y(n_9), .A(in_8[0]));
  INVX1 g229(.Y(n_8), .A(in_22[1]));
  INVX1 g230(.Y(n_7), .A(in_11[1]));
  INVX1 g231(.Y(n_6), .A(in_0[0]));
  INVX1 g232(.Y(n_5), .A(in_19[0]));
  INVX1 g233(.Y(n_4), .A(in_20[0]));
  INVX1 g234(.Y(n_3), .A(in_21[1]));
  INVX1 g235(.Y(n_2), .A(in_13[0]));
  INVX1 g236(.Y(n_1), .A(in_2[0]));
endmodule

module WALLACE_CSA_DUMMY_OP86_group_109840(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, out_0);
input  in_25, in_26, in_44, in_65, in_69;
input   [4:0] in_0;
input   [2:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [7:0] in_4;
input   [7:0] in_5;
input   [6:0] in_6;
input   [6:0] in_7;
input   [6:0] in_8;
input   [6:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [4:0] in_23;
input   [5:0] in_24;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [1:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
input   [4:0] in_42;
input   [1:0] in_43;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [1:0] in_48;
input   [4:0] in_49;
input   [2:0] in_50;
input   [4:0] in_51;
input   [2:0] in_52;
input   [1:0] in_53;
input   [1:0] in_54;
input   [2:0] in_55;
input   [4:0] in_56;
input   [1:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [3:0] in_62;
input   [2:0] in_63;
input   [4:0] in_64;
input   [1:0] in_66;
input   [4:0] in_67;
input   [1:0] in_68;
input   [4:0] in_70;
input   [2:0] in_71;
output  [9:0] out_0;
wire  n_291, n_289, n_287, n_285, n_283, n_282, n_281, n_279, n_278, n_277, 
    n_276, n_275, n_274, n_273, n_271, n_270, n_269, n_268, n_267, n_266, 
    n_265, n_264, n_263, n_262, n_261, n_259, n_258, n_257, n_256, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, 
    n_244, n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, 
    n_234, n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, 
    n_224, n_223, n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, 
    n_214, n_213, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, 
    n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 
    n_193, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, 
    n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, 
    n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, 
    n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, 
    n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, 
    n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, 
    n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, 
    n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
    n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_69, in_65, in_44, in_26, in_25;
wire   [9:0] out_0;
wire   [3:0] in_62;
wire   [1:0] in_68;
wire   [1:0] in_66;
wire   [1:0] in_61;
wire   [1:0] in_57;
wire   [1:0] in_54;
wire   [1:0] in_53;
wire   [1:0] in_48;
wire   [1:0] in_43;
wire   [1:0] in_41;
wire   [1:0] in_38;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_24;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [6:0] in_9;
wire   [6:0] in_8;
wire   [6:0] in_7;
wire   [6:0] in_6;
wire   [7:0] in_5;
wire   [7:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [2:0] in_71;
wire   [2:0] in_63;
wire   [2:0] in_55;
wire   [2:0] in_52;
wire   [2:0] in_50;
wire   [2:0] in_1;
wire   [4:0] in_70;
wire   [4:0] in_67;
wire   [4:0] in_64;
wire   [4:0] in_60;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_56;
wire   [4:0] in_51;
wire   [4:0] in_49;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_42;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_23;
wire   [4:0] in_0;
  INVX1 g9189(.Y(out_0[9]), .A(n_291));
  ADDFX1 g9190(.CO(n_291), .S(out_0[8]), .A(n_34), .B(n_251), .CI(n_289));
  ADDFX1 g9191(.CO(n_289), .S(out_0[7]), .A(n_252), .B(n_277), .CI(n_287));
  ADDFX1 g9192(.CO(n_287), .S(out_0[6]), .A(n_281), .B(n_278), .CI(n_285));
  ADDFX1 g9193(.CO(n_285), .S(out_0[5]), .A(n_275), .B(n_282), .CI(n_283));
  ADDFX1 g9194(.CO(n_283), .S(out_0[4]), .A(n_273), .B(n_276), .CI(n_279));
  ADDFX1 g9195(.CO(n_281), .S(n_282), .A(n_256), .B(n_267), .CI(n_270));
  ADDFX1 g9196(.CO(n_279), .S(out_0[3]), .A(n_257), .B(n_271), .CI(n_274));
  ADDFX1 g9197(.CO(n_277), .S(n_278), .A(n_255), .B(n_236), .CI(n_269));
  ADDFX1 g9198(.CO(n_275), .S(n_276), .A(n_268), .B(n_266), .CI(n_263));
  ADDFX1 g9199(.CO(n_273), .S(n_274), .A(n_262), .B(n_249), .CI(n_264));
  ADDFX1 g9200(.CO(n_271), .S(out_0[2]), .A(n_259), .B(n_258), .CI(n_250));
  ADDFX1 g9201(.CO(n_269), .S(n_270), .A(n_253), .B(n_232), .CI(n_265));
  ADDFX1 g9202(.CO(n_267), .S(n_268), .A(n_245), .B(n_254), .CI(n_261));
  ADDFX1 g9203(.CO(n_265), .S(n_266), .A(n_208), .B(n_247), .CI(n_242));
  ADDFX1 g9204(.CO(n_263), .S(n_264), .A(n_243), .B(n_246), .CI(n_248));
  ADDFX1 g9205(.CO(n_261), .S(n_262), .A(n_238), .B(n_233), .CI(n_210));
  ADDFX1 g9206(.CO(n_259), .S(out_0[1]), .A(n_211), .B(n_240), .CI(n_226));
  ADDFX1 g9207(.CO(n_257), .S(n_258), .A(n_239), .B(n_225), .CI(n_244));
  ADDFX1 g9208(.CO(n_255), .S(n_256), .A(n_219), .B(n_207), .CI(n_241));
  ADDFX1 g9209(.CO(n_253), .S(n_254), .A(n_221), .B(n_237), .CI(n_209));
  ADDFX1 g9210(.CO(n_251), .S(n_252), .A(n_38), .B(n_37), .CI(n_235));
  ADDFX1 g9211(.CO(n_249), .S(n_250), .A(n_216), .B(n_234), .CI(n_230));
  ADDFX1 g9212(.CO(n_247), .S(n_248), .A(n_217), .B(n_227), .CI(in_2[3]));
  ADDFX1 g9213(.CO(n_245), .S(n_246), .A(n_215), .B(n_222), .CI(n_229));
  ADDFX1 g9214(.CO(n_243), .S(n_244), .A(n_218), .B(n_205), .CI(n_228));
  ADDFX1 g9215(.CO(n_241), .S(n_242), .A(n_223), .B(n_220), .CI(in_2[4]));
  ADDFX1 g9216(.CO(n_239), .S(n_240), .A(n_201), .B(n_214), .CI(n_206));
  ADDFX1 g9217(.CO(n_237), .S(n_238), .A(n_224), .B(n_183), .CI(n_168));
  ADDFX1 g9218(.CO(n_235), .S(n_236), .A(n_203), .B(n_39), .CI(n_231));
  ADDFX1 g9219(.CO(n_233), .S(n_234), .A(n_184), .B(n_213), .CI(n_173));
  ADDFX1 g9220(.CO(n_231), .S(n_232), .A(n_204), .B(in_3[5]), .CI(in_2[5]));
  ADDFX1 g9221(.CO(n_229), .S(n_230), .A(n_166), .B(n_199), .CI(in_2[2]));
  ADDFX1 g9222(.CO(n_227), .S(n_228), .A(n_198), .B(n_193), .CI(in_3[2]));
  ADDFX1 g9223(.CO(n_225), .S(n_226), .A(n_192), .B(n_174), .CI(n_200));
  ADDFX1 g9224(.CO(n_223), .S(n_224), .A(n_197), .B(n_189), .CI(n_177));
  ADDFX1 g9225(.CO(n_221), .S(n_222), .A(n_176), .B(n_165), .CI(n_164));
  ADDFX1 g9226(.CO(n_219), .S(n_220), .A(n_175), .B(n_163), .CI(n_167));
  ADDFX1 g9227(.CO(n_217), .S(n_218), .A(n_195), .B(n_181), .CI(n_190));
  ADDFX1 g9228(.CO(n_215), .S(n_216), .A(n_191), .B(n_178), .CI(n_188));
  ADDFX1 g9229(.CO(n_213), .S(n_214), .A(n_182), .B(n_194), .CI(n_115));
  ADDHX1 g9230(.CO(n_211), .S(out_0[0]), .A(n_170), .B(n_202));
  ADDFX1 g9231(.CO(n_209), .S(n_210), .A(n_187), .B(n_186), .CI(in_3[3]));
  ADDFX1 g9232(.CO(n_207), .S(n_208), .A(n_180), .B(n_185), .CI(in_3[4]));
  ADDFX1 g9233(.CO(n_205), .S(n_206), .A(n_196), .B(n_171), .CI(n_169));
  ADDHX1 g9234(.CO(n_203), .S(n_204), .A(n_161), .B(n_179));
  ADDFX1 g9235(.CO(n_201), .S(n_202), .A(n_160), .B(n_172), .CI(n_116));
  ADDFX1 g9236(.CO(n_199), .S(n_200), .A(n_126), .B(n_159), .CI(in_2[1]));
  ADDFX1 g9237(.CO(n_197), .S(n_198), .A(n_139), .B(n_157), .CI(n_137));
  ADDFX1 g9238(.CO(n_195), .S(n_196), .A(n_150), .B(n_138), .CI(n_158));
  ADDFX1 g9239(.CO(n_193), .S(n_194), .A(n_113), .B(n_151), .CI(n_155));
  ADDFX1 g9240(.CO(n_191), .S(n_192), .A(n_112), .B(n_154), .CI(n_142));
  ADDFX1 g9241(.CO(n_189), .S(n_190), .A(n_149), .B(n_106), .CI(n_135));
  ADDFX1 g9242(.CO(n_187), .S(n_188), .A(n_134), .B(n_153), .CI(n_109));
  ADDFX1 g9243(.CO(n_185), .S(n_186), .A(n_120), .B(n_128), .CI(n_123));
  ADDFX1 g9244(.CO(n_183), .S(n_184), .A(n_132), .B(n_147), .CI(n_130));
  ADDFX1 g9245(.CO(n_181), .S(n_182), .A(n_140), .B(n_143), .CI(n_136));
  ADDFX1 g9246(.CO(n_179), .S(n_180), .A(n_127), .B(n_121), .CI(n_162));
  ADDFX1 g9247(.CO(n_177), .S(n_178), .A(n_146), .B(n_111), .CI(n_141));
  ADDFX1 g9248(.CO(n_175), .S(n_176), .A(n_133), .B(n_145), .CI(in_4[3]));
  ADDFX1 g9249(.CO(n_173), .S(n_174), .A(n_110), .B(n_148), .CI(in_3[1]));
  ADDFX1 g9250(.CO(n_171), .S(n_172), .A(n_114), .B(n_144), .CI(n_53));
  ADDFX1 g9251(.CO(n_169), .S(n_170), .A(n_156), .B(n_152), .CI(in_3[0]));
  ADDFX1 g9252(.CO(n_167), .S(n_168), .A(n_131), .B(n_122), .CI(n_129));
  ADDFX1 g9253(.CO(n_165), .S(n_166), .A(n_125), .B(n_108), .CI(n_124));
  ADDFX1 g9254(.CO(n_163), .S(n_164), .A(n_105), .B(n_107), .CI(n_4));
  ADDFX1 g9255(.CO(n_161), .S(n_162), .A(n_35), .B(n_119), .CI(n_29));
  ADDFX1 g9256(.CO(n_159), .S(n_160), .A(n_96), .B(in_8[0]), .CI(n_61));
  ADDFX1 g9257(.CO(n_157), .S(n_158), .A(n_70), .B(n_91), .CI(n_66));
  ADDFX1 g9258(.CO(n_155), .S(n_156), .A(n_43), .B(n_67), .CI(n_92));
  ADDFX1 g9259(.CO(n_153), .S(n_154), .A(n_104), .B(n_47), .CI(in_8[1]));
  ADDFX1 g9260(.CO(n_151), .S(n_152), .A(n_90), .B(n_45), .CI(n_83));
  ADDFX1 g9261(.CO(n_149), .S(n_150), .A(in_20[1]), .B(n_82), .CI(n_78));
  ADDFX1 g9262(.CO(n_147), .S(n_148), .A(n_98), .B(n_68), .CI(n_52));
  ADDFX1 g9263(.CO(n_145), .S(n_146), .A(n_46), .B(n_80), .CI(n_64));
  ADDFX1 g9264(.CO(n_143), .S(n_144), .A(n_79), .B(n_94), .CI(n_71));
  ADDFX1 g9265(.CO(n_141), .S(n_142), .A(n_81), .B(n_49), .CI(in_9[1]));
  ADDFX1 g9266(.CO(n_139), .S(n_140), .A(n_44), .B(n_95), .CI(n_42));
  ADDFX1 g9267(.CO(n_137), .S(n_138), .A(n_56), .B(n_89), .CI(n_93));
  ADDFX1 g9268(.CO(n_135), .S(n_136), .A(n_87), .B(n_72), .CI(in_7[1]));
  ADDFX1 g9269(.CO(n_133), .S(n_134), .A(n_48), .B(n_101), .CI(n_103));
  ADDFX1 g9270(.CO(n_131), .S(n_132), .A(n_97), .B(n_86), .CI(in_8[2]));
  ADDFX1 g9271(.CO(n_129), .S(n_130), .A(n_40), .B(n_100), .CI(in_4[2]));
  ADDFX1 g9272(.CO(n_127), .S(n_128), .A(n_54), .B(n_6), .CI(n_27));
  ADDFX1 g9273(.CO(n_125), .S(n_126), .A(n_58), .B(n_41), .CI(n_75));
  ADDFX1 g9274(.CO(n_123), .S(n_124), .A(n_55), .B(n_84), .CI(in_5[2]));
  ADDFX1 g9275(.CO(n_121), .S(n_122), .A(n_99), .B(n_85), .CI(n_20));
  INVX1 g9276(.Y(n_120), .A(n_118));
  INVX1 g9277(.Y(n_119), .A(n_117));
  ADDFX1 g9278(.CO(n_117), .S(n_118), .A(in_35[2]), .B(n_50), .CI(n_36));
  ADDFX1 g9279(.CO(n_115), .S(n_116), .A(n_69), .B(n_59), .CI(in_2[0]));
  ADDFX1 g9280(.CO(n_113), .S(n_114), .A(n_88), .B(n_73), .CI(n_57));
  ADDFX1 g9281(.CO(n_111), .S(n_112), .A(n_102), .B(n_77), .CI(n_65));
  ADDFX1 g9282(.CO(n_109), .S(n_110), .A(n_60), .B(in_4[1]), .CI(in_5[1]));
  ADDFX1 g9283(.CO(n_107), .S(n_108), .A(n_74), .B(in_7[2]), .CI(in_9[2]));
  ADDFX1 g9284(.CO(n_105), .S(n_106), .A(in_14[2]), .B(in_11[2]), .CI(n_76));
  ADDFX1 g9285(.CO(n_103), .S(n_104), .A(in_68[1]), .B(n_21), .CI(n_3));
  ADDFX1 g9286(.CO(n_101), .S(n_102), .A(in_50[0]), .B(n_26), .CI(in_52[0]));
  ADDFX1 g9287(.CO(n_99), .S(n_100), .A(in_35[2]), .B(n_10), .CI(n_13));
  ADDFX1 g9288(.CO(n_97), .S(n_98), .A(n_33), .B(in_19[1]), .CI(in_15[1]));
  ADDFX1 g9289(.CO(n_95), .S(n_96), .A(in_57[0]), .B(n_15), .CI(in_69));
  ADDFX1 g9290(.CO(n_93), .S(n_94), .A(in_14[0]), .B(in_31[0]), .CI(n_31));
  ADDFX1 g9291(.CO(n_91), .S(n_92), .A(in_34[0]), .B(n_25), .CI(in_64[0]));
  ADDFX1 g9292(.CO(n_89), .S(n_90), .A(in_25), .B(n_23), .CI(n_16));
  ADDFX1 g9293(.CO(n_87), .S(n_88), .A(n_24), .B(n_14), .CI(in_52[0]));
  INVX1 g9294(.Y(n_86), .A(n_63));
  INVX1 g9295(.Y(n_85), .A(n_62));
  INVX1 g9296(.Y(n_84), .A(n_51));
  ADDFX1 g9297(.CO(n_82), .S(n_83), .A(in_6[0]), .B(in_45[0]), .CI(in_48[0]));
  ADDFX1 g9298(.CO(n_80), .S(n_81), .A(in_55[1]), .B(n_22), .CI(in_63[1]));
  ADDFX1 g9299(.CO(n_78), .S(n_79), .A(in_15[0]), .B(in_21[0]), .CI(in_41[0]));
  ADDFX1 g9300(.CO(n_76), .S(n_77), .A(in_11[1]), .B(n_19), .CI(in_54[1]));
  ADDFX1 g9301(.CO(n_74), .S(n_75), .A(in_22[1]), .B(in_23[1]), .CI(in_29[1]));
  ADDFX1 g9302(.CO(n_72), .S(n_73), .A(in_50[0]), .B(in_28[0]), .CI(in_71[0]));
  ADDFX1 g9303(.CO(n_70), .S(n_71), .A(in_19[0]), .B(in_38[0]), .CI(in_61[0]));
  ADDFX1 g9304(.CO(n_68), .S(n_69), .A(in_29[0]), .B(in_24[0]), .CI(in_9[0]));
  ADDFX1 g9305(.CO(n_66), .S(n_67), .A(in_44), .B(n_7), .CI(in_65));
  ADDFX1 g9306(.CO(n_64), .S(n_65), .A(in_14[0]), .B(in_43[0]), .CI(in_71[0]));
  ADDFX1 g9307(.CO(n_62), .S(n_63), .A(in_45[0]), .B(in_19[2]), .CI(in_15[2]));
  ADDFX1 g9308(.CO(n_60), .S(n_61), .A(in_22[0]), .B(in_17[0]), .CI(in_23[0]));
  ADDFX1 g9309(.CO(n_58), .S(n_59), .A(n_0), .B(in_11[0]), .CI(in_27[0]));
  ADDFX1 g9310(.CO(n_56), .S(n_57), .A(in_20[0]), .B(n_2), .CI(n_32));
  ADDFX1 g9311(.CO(n_54), .S(n_55), .A(in_62[2]), .B(n_18), .CI(n_1));
  ADDFX1 g9312(.CO(n_52), .S(n_53), .A(in_5[0]), .B(in_7[0]), .CI(in_4[0]));
  ADDFX1 g9313(.CO(n_50), .S(n_51), .A(in_13[2]), .B(in_16[2]), .CI(in_70[0]));
  ADDFX1 g9314(.CO(n_48), .S(n_49), .A(in_53[1]), .B(in_1[1]), .CI(n_30));
  ADDFX1 g9315(.CO(n_46), .S(n_47), .A(in_6[1]), .B(n_9), .CI(in_66[1]));
  ADDFX1 g9316(.CO(n_44), .S(n_45), .A(n_8), .B(n_11), .CI(in_70[0]));
  ADDFX1 g9317(.CO(n_42), .S(n_43), .A(n_12), .B(n_5), .CI(in_43[0]));
  ADDFX1 g9318(.CO(n_40), .S(n_41), .A(in_26), .B(n_28), .CI(n_17));
  ADDHX1 g9319(.CO(n_38), .S(n_39), .A(in_3[6]), .B(in_2[6]));
  OAI21X1 g9320(.Y(n_37), .A0(in_3[7]), .A1(in_2[6]), .B0(n_34));
  XNOR2X1 g9321(.Y(n_36), .A(in_11[3]), .B(in_14[3]));
  NOR2X1 g9322(.Y(n_35), .A(in_11[3]), .B(in_14[3]));
  NAND2X1 g9323(.Y(n_34), .A(in_3[7]), .B(in_2[6]));
  INVX1 g9324(.Y(n_33), .A(in_24[1]));
  INVX1 g9325(.Y(n_32), .A(in_56[0]));
  INVX1 g9326(.Y(n_31), .A(in_58[0]));
  INVX1 g9327(.Y(n_30), .A(in_60[1]));
  INVX1 g9328(.Y(n_29), .A(in_4[4]));
  INVX1 g9329(.Y(n_28), .A(in_17[1]));
  INVX1 g9330(.Y(n_27), .A(in_9[3]));
  INVX1 g9331(.Y(n_26), .A(in_0[1]));
  INVX1 g9332(.Y(n_25), .A(in_18[0]));
  INVX1 g9333(.Y(n_24), .A(in_12[0]));
  INVX1 g9334(.Y(n_23), .A(in_47[0]));
  INVX1 g9335(.Y(n_22), .A(in_10[1]));
  INVX1 g9336(.Y(n_21), .A(in_40[1]));
  INVX1 g9337(.Y(n_20), .A(in_8[3]));
  INVX1 g9338(.Y(n_19), .A(in_51[1]));
  INVX1 g9339(.Y(n_18), .A(in_34[0]));
  INVX1 g9340(.Y(n_17), .A(in_27[1]));
  INVX1 g9341(.Y(n_16), .A(in_59[0]));
  INVX1 g9342(.Y(n_15), .A(in_67[0]));
  INVX1 g9343(.Y(n_14), .A(in_37[0]));
  INVX1 g9344(.Y(n_13), .A(in_29[2]));
  INVX1 g9345(.Y(n_12), .A(in_42[0]));
  INVX1 g9346(.Y(n_11), .A(in_39[0]));
  INVX1 g9347(.Y(n_10), .A(in_20[2]));
  INVX1 g9348(.Y(n_9), .A(in_30[1]));
  INVX1 g9349(.Y(n_8), .A(in_36[0]));
  INVX1 g9350(.Y(n_7), .A(in_33[0]));
  INVX1 g9351(.Y(n_6), .A(in_7[3]));
  INVX1 g9352(.Y(n_5), .A(in_32[0]));
  INVX1 g9353(.Y(n_4), .A(in_5[3]));
  INVX1 g9354(.Y(n_3), .A(in_46[1]));
  INVX1 g9355(.Y(n_2), .A(in_49[0]));
  INVX1 g9356(.Y(n_1), .A(in_64[0]));
  INVX1 g9357(.Y(n_0), .A(in_26));
endmodule

module WALLACE_CSA_DUMMY_OP89_group_106209(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, out_0);
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [9:0] in_3;
input   [6:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [2:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [2:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [2:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
input   [4:0] in_41;
input   [1:0] in_42;
output  [9:0] out_0;
wire  n_152, n_150, n_148, n_146, n_144, n_143, n_142, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_0;
wire   [9:0] out_0;
wire   [1:0] in_42;
wire   [1:0] in_40;
wire   [1:0] in_37;
wire   [2:0] in_34;
wire   [2:0] in_31;
wire   [2:0] in_25;
wire   [2:0] in_18;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [6:0] in_4;
wire   [9:0] in_3;
wire   [4:0] in_41;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_17;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  OAI2BB1X1 g1970(.Y(out_0[9]), .A0N(in_3[6]), .A1N(n_67), .B0(n_152));
  ADDFX1 g1971(.CO(n_152), .S(out_0[6]), .A(n_83), .B(n_138), .CI(n_150));
  ADDFX1 g1972(.CO(n_150), .S(out_0[5]), .A(n_142), .B(n_139), .CI(n_148));
  ADDFX1 g1973(.CO(n_148), .S(out_0[4]), .A(n_140), .B(n_143), .CI(n_146));
  ADDFX1 g1974(.CO(n_146), .S(out_0[3]), .A(n_136), .B(n_144), .CI(n_141));
  ADDFX1 g1975(.CO(n_144), .S(out_0[2]), .A(n_129), .B(n_134), .CI(n_137));
  ADDFX1 g1976(.CO(n_142), .S(n_143), .A(n_126), .B(n_132), .CI(n_131));
  ADDFX1 g1977(.CO(n_140), .S(n_141), .A(n_128), .B(n_127), .CI(n_133));
  ADDFX1 g1978(.CO(n_138), .S(n_139), .A(n_120), .B(n_130), .CI(n_68));
  ADDFX1 g1979(.CO(n_136), .S(n_137), .A(n_111), .B(n_122), .CI(n_125));
  ADDFX1 g1980(.CO(n_134), .S(out_0[1]), .A(n_116), .B(n_123), .CI(n_109));
  ADDFX1 g1981(.CO(n_132), .S(n_133), .A(n_110), .B(n_119), .CI(n_124));
  ADDFX1 g1982(.CO(n_130), .S(n_131), .A(n_118), .B(n_121), .CI(in_3[4]));
  ADDFX1 g1983(.CO(n_128), .S(n_129), .A(n_105), .B(n_112), .CI(n_108));
  ADDFX1 g1984(.CO(n_126), .S(n_127), .A(n_115), .B(n_104), .CI(in_3[3]));
  ADDFX1 g1985(.CO(n_124), .S(n_125), .A(n_102), .B(n_107), .CI(in_3[2]));
  ADDFX1 g1986(.CO(n_122), .S(n_123), .A(n_103), .B(n_113), .CI(n_98));
  ADDFX1 g1987(.CO(n_120), .S(n_121), .A(n_24), .B(n_96), .CI(n_114));
  ADDFX1 g1988(.CO(n_118), .S(n_119), .A(n_90), .B(n_75), .CI(n_106));
  ADDFX1 g1989(.CO(n_116), .S(out_0[0]), .A(n_89), .B(n_78), .CI(n_99));
  ADDFX1 g1990(.CO(n_114), .S(n_115), .A(n_48), .B(n_94), .CI(n_97));
  ADDFX1 g1991(.CO(n_112), .S(n_113), .A(n_93), .B(n_74), .CI(n_77));
  ADDFX1 g1992(.CO(n_110), .S(n_111), .A(n_81), .B(n_76), .CI(n_100));
  ADDFX1 g1993(.CO(n_108), .S(n_109), .A(n_82), .B(n_101), .CI(in_3[1]));
  ADDFX1 g1994(.CO(n_106), .S(n_107), .A(n_79), .B(n_92), .CI(n_86));
  ADDFX1 g1995(.CO(n_104), .S(n_105), .A(n_95), .B(n_73), .CI(n_91));
  ADDFX1 g1996(.CO(n_102), .S(n_103), .A(n_80), .B(n_87), .CI(n_84));
  ADDFX1 g1997(.CO(n_100), .S(n_101), .A(n_62), .B(n_41), .CI(n_88));
  ADDFX1 g1998(.CO(n_98), .S(n_99), .A(n_51), .B(n_85), .CI(in_3[0]));
  ADDFX1 g1999(.CO(n_96), .S(n_97), .A(n_60), .B(n_27), .CI(n_71));
  ADDFX1 g2000(.CO(n_94), .S(n_95), .A(n_56), .B(n_34), .CI(n_69));
  ADDFX1 g2001(.CO(n_92), .S(n_93), .A(n_46), .B(n_44), .CI(n_25));
  ADDFX1 g2002(.CO(n_90), .S(n_91), .A(n_36), .B(n_61), .CI(n_72));
  ADDFX1 g2003(.CO(n_88), .S(n_89), .A(n_47), .B(n_43), .CI(n_53));
  ADDFX1 g2004(.CO(n_86), .S(n_87), .A(in_7[1]), .B(n_32), .CI(n_70));
  ADDFX1 g2005(.CO(n_84), .S(n_85), .A(n_33), .B(n_65), .CI(n_26));
  XNOR2X1 g2006(.Y(n_83), .A(in_3[6]), .B(n_67));
  ADDFX1 g2007(.CO(n_81), .S(n_82), .A(n_37), .B(n_39), .CI(n_50));
  ADDFX1 g2008(.CO(n_79), .S(n_80), .A(n_30), .B(n_42), .CI(n_64));
  ADDFX1 g2009(.CO(n_77), .S(n_78), .A(n_45), .B(n_31), .CI(n_63));
  ADDFX1 g2010(.CO(n_75), .S(n_76), .A(n_40), .B(n_38), .CI(n_49));
  ADDFX1 g2011(.CO(n_73), .S(n_74), .A(n_52), .B(n_57), .CI(n_35));
  ADDFX1 g2012(.CO(n_71), .S(n_72), .A(in_9[2]), .B(n_2), .CI(n_23));
  ADDFX1 g2013(.CO(n_69), .S(n_70), .A(in_11[1]), .B(n_5), .CI(n_21));
  NAND2BX1 g2014(.Y(n_68), .AN(n_67), .B(n_66));
  NOR2XL g2015(.Y(n_67), .A(n_0), .B(in_3[5]));
  NAND2XL g2016(.Y(n_66), .A(n_0), .B(in_3[5]));
  ADDFX1 g2017(.CO(n_64), .S(n_65), .A(in_8[0]), .B(n_15), .CI(in_10[0]));
  ADDFX1 g2019(.CO(n_62), .S(n_63), .A(in_4[0]), .B(in_13[0]), .CI(in_7[0]));
  INVX1 g2020(.Y(n_61), .A(n_59));
  INVX1 g2021(.Y(n_60), .A(n_58));
  ADDFX1 g2022(.CO(n_58), .S(n_59), .A(in_32[0]), .B(in_39[0]), .CI(in_20[2]));
  INVX1 g2023(.Y(n_57), .A(n_55));
  INVX1 g2024(.Y(n_56), .A(n_54));
  ADDFX1 g2025(.CO(n_54), .S(n_55), .A(in_1[1]), .B(in_27[1]), .CI(in_35[1]));
  INVX1 g2026(.Y(n_53), .A(n_29));
  INVX1 g2027(.Y(n_52), .A(n_28));
  ADDFX1 g2028(.CO(n_50), .S(n_51), .A(n_18), .B(in_16[0]), .CI(in_6[0]));
  ADDFX1 g2029(.CO(n_48), .S(n_49), .A(in_7[2]), .B(n_7), .CI(in_10[2]));
  ADDFX1 g2030(.CO(n_46), .S(n_47), .A(in_5[0]), .B(n_6), .CI(n_17));
  ADDFX1 g2031(.CO(n_44), .S(n_45), .A(n_3), .B(in_26[0]), .CI(in_39[0]));
  ADDFX1 g2032(.CO(n_42), .S(n_43), .A(in_32[0]), .B(n_11), .CI(in_37[0]));
  ADDFX1 g2033(.CO(n_40), .S(n_41), .A(in_4[1]), .B(n_8), .CI(in_15[1]));
  ADDFX1 g2034(.CO(n_38), .S(n_39), .A(in_25[1]), .B(n_12), .CI(n_4));
  ADDFX1 g2035(.CO(n_36), .S(n_37), .A(in_18[1]), .B(in_31[0]), .CI(in_34[1]));
  ADDFX1 g2036(.CO(n_34), .S(n_35), .A(in_10[1]), .B(n_16), .CI(n_14));
  ADDFX1 g2037(.CO(n_32), .S(n_33), .A(in_15[0]), .B(n_13), .CI(in_40[0]));
  ADDFX1 g2038(.CO(n_30), .S(n_31), .A(n_10), .B(n_9), .CI(in_42[0]));
  ADDFX1 g2039(.CO(n_28), .S(n_29), .A(in_0[0]), .B(in_17[0]), .CI(in_41[0]));
  OAI21X1 g2040(.Y(n_27), .A0(n_20), .A1(in_10[3]), .B0(n_0));
  OAI2BB1X1 g2041(.Y(n_26), .A0N(in_31[0]), .A1N(n_22), .B0(n_25));
  OR2X1 g2042(.Y(n_25), .A(in_31[0]), .B(n_22));
  INVX1 g2043(.Y(n_24), .A(n_0));
  NAND2X1 g2044(.Y(n_0), .A(n_20), .B(in_10[3]));
  OAI21X1 g2045(.Y(n_23), .A0(in_12[0]), .A1(in_11[1]), .B0(n_19));
  XNOR2X1 g2046(.Y(n_22), .A(in_12[0]), .B(in_14[0]));
  NOR2BX1 g2047(.Y(n_21), .AN(in_12[0]), .B(in_14[0]));
  INVX1 g2048(.Y(n_20), .A(n_19));
  NAND2XL g2049(.Y(n_19), .A(in_12[0]), .B(in_11[1]));
  INVX1 g2050(.Y(n_18), .A(in_19[0]));
  INVX1 g2051(.Y(n_17), .A(in_28[0]));
  INVX1 g2052(.Y(n_16), .A(in_29[1]));
  INVX1 g2053(.Y(n_15), .A(in_2[0]));
  INVX1 g2054(.Y(n_14), .A(in_21[1]));
  INVX1 g2055(.Y(n_13), .A(in_24[0]));
  INVX1 g2056(.Y(n_12), .A(in_16[1]));
  INVX1 g2057(.Y(n_11), .A(in_33[0]));
  INVX1 g2058(.Y(n_10), .A(in_38[0]));
  INVX1 g2059(.Y(n_9), .A(in_23[0]));
  INVX1 g2060(.Y(n_8), .A(in_6[1]));
  INVX1 g2061(.Y(n_7), .A(in_15[2]));
  INVX1 g2062(.Y(n_6), .A(in_22[0]));
  INVX1 g2063(.Y(n_5), .A(in_30[1]));
  INVX1 g2064(.Y(n_4), .A(in_13[1]));
  INVX1 g2065(.Y(n_3), .A(in_36[0]));
  INVX1 g2066(.Y(n_2), .A(in_26[0]));
endmodule

module WALLACE_CSA_DUMMY_OP91_group_109814(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, out_0);
input  in_32, in_33, in_37, in_41;
input   [4:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [6:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [5:0] in_21;
input   [4:0] in_22;
input   [2:0] in_23;
input   [1:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [1:0] in_28;
input   [4:0] in_29;
input   [1:0] in_30;
input   [4:0] in_31;
input   [4:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [4:0] in_38;
input   [2:0] in_39;
input   [4:0] in_40;
input   [1:0] in_42;
output  [9:0] out_0;
wire  n_167, n_165, n_163, n_161, n_159, n_158, n_157, n_156, n_155, n_154, 
    n_153, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
    n_142, n_141, n_140, n_139, n_137, n_136, n_135, n_134, n_133, n_132, 
    n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_119, n_118, n_117, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, n_0, in_41, in_37, in_33, in_32;
wire   [9:0] out_0;
wire   [1:0] in_42;
wire   [1:0] in_36;
wire   [1:0] in_30;
wire   [1:0] in_28;
wire   [1:0] in_24;
wire   [2:0] in_39;
wire   [2:0] in_23;
wire   [5:0] in_21;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [6:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  NAND2X1 g2145(.Y(out_0[9]), .A(n_63), .B(n_167));
  ADDFX1 g2146(.CO(n_167), .S(out_0[7]), .A(n_149), .B(n_64), .CI(n_165));
  ADDFX1 g2147(.CO(n_165), .S(out_0[6]), .A(n_157), .B(n_150), .CI(n_163));
  ADDFX1 g2148(.CO(n_163), .S(out_0[5]), .A(n_158), .B(n_155), .CI(n_161));
  ADDFX1 g2149(.CO(n_161), .S(out_0[4]), .A(n_153), .B(n_156), .CI(n_159));
  ADDFX1 g2150(.CO(n_159), .S(out_0[3]), .A(n_139), .B(n_151), .CI(n_154));
  ADDFX1 g2151(.CO(n_157), .S(n_158), .A(n_148), .B(in_2[5]), .CI(n_145));
  ADDFX1 g2152(.CO(n_155), .S(n_156), .A(n_136), .B(n_143), .CI(n_146));
  ADDFX1 g2153(.CO(n_153), .S(n_154), .A(n_134), .B(n_141), .CI(n_144));
  ADDFX1 g2154(.CO(n_151), .S(out_0[2]), .A(n_142), .B(n_137), .CI(n_140));
  ADDFX1 g2155(.CO(n_149), .S(n_150), .A(n_26), .B(n_147), .CI(in_2[6]));
  ADDFX1 g2156(.CO(n_147), .S(n_148), .A(n_119), .B(n_135), .CI(n_22));
  ADDFX1 g2157(.CO(n_145), .S(n_146), .A(n_131), .B(n_133), .CI(in_2[4]));
  ADDFX1 g2158(.CO(n_143), .S(n_144), .A(n_132), .B(n_129), .CI(in_2[3]));
  ADDFX1 g2159(.CO(n_141), .S(n_142), .A(n_126), .B(n_101), .CI(n_121));
  ADDFX1 g2160(.CO(n_139), .S(n_140), .A(n_127), .B(n_130), .CI(in_2[2]));
  ADDFX1 g2161(.CO(n_137), .S(out_0[1]), .A(n_115), .B(n_128), .CI(n_122));
  ADDFX1 g2162(.CO(n_135), .S(n_136), .A(n_120), .B(in_3[4]), .CI(n_123));
  ADDFX1 g2163(.CO(n_133), .S(n_134), .A(n_125), .B(n_117), .CI(n_124));
  ADDFX1 g2164(.CO(n_131), .S(n_132), .A(n_113), .B(n_108), .CI(n_111));
  ADDFX1 g2165(.CO(n_129), .S(n_130), .A(n_112), .B(n_97), .CI(n_118));
  ADDFX1 g2166(.CO(n_127), .S(n_128), .A(n_99), .B(n_98), .CI(n_102));
  ADDFX1 g2167(.CO(n_125), .S(n_126), .A(n_114), .B(n_110), .CI(n_103));
  ADDFX1 g2168(.CO(n_123), .S(n_124), .A(n_79), .B(n_109), .CI(in_3[3]));
  ADDFX1 g2169(.CO(n_121), .S(n_122), .A(n_106), .B(n_104), .CI(in_2[1]));
  ADDFX1 g2170(.CO(n_119), .S(n_120), .A(in_27[0]), .B(n_69), .CI(n_107));
  ADDFX1 g2171(.CO(n_117), .S(n_118), .A(n_85), .B(n_105), .CI(in_3[2]));
  ADDHX1 g2172(.CO(n_115), .S(out_0[0]), .A(n_100), .B(n_96));
  ADDFX1 g2173(.CO(n_113), .S(n_114), .A(n_73), .B(n_91), .CI(n_71));
  ADDFX1 g2174(.CO(n_111), .S(n_112), .A(n_94), .B(n_80), .CI(n_87));
  ADDFX1 g2175(.CO(n_109), .S(n_110), .A(n_42), .B(n_89), .CI(n_66));
  ADDFX1 g2176(.CO(n_107), .S(n_108), .A(n_65), .B(n_93), .CI(n_70));
  ADDFX1 g2177(.CO(n_105), .S(n_106), .A(n_74), .B(n_90), .CI(n_81));
  ADDFX1 g2178(.CO(n_103), .S(n_104), .A(n_83), .B(n_92), .CI(n_77));
  ADDFX1 g2179(.CO(n_101), .S(n_102), .A(n_75), .B(n_88), .CI(n_95));
  ADDFX1 g2180(.CO(n_99), .S(n_100), .A(n_78), .B(n_82), .CI(n_76));
  ADDFX1 g2181(.CO(n_97), .S(n_98), .A(n_72), .B(n_86), .CI(in_3[1]));
  ADDFX1 g2182(.CO(n_95), .S(n_96), .A(n_84), .B(in_3[0]), .CI(in_2[0]));
  ADDFX1 g2183(.CO(n_93), .S(n_94), .A(n_47), .B(n_55), .CI(n_35));
  ADDFX1 g2184(.CO(n_91), .S(n_92), .A(n_37), .B(n_53), .CI(n_33));
  ADDFX1 g2185(.CO(n_89), .S(n_90), .A(n_57), .B(n_49), .CI(n_59));
  ADDFX1 g2186(.CO(n_87), .S(n_88), .A(n_39), .B(n_61), .CI(n_52));
  ADDFX1 g2187(.CO(n_85), .S(n_86), .A(n_31), .B(n_44), .CI(n_68));
  ADDFX1 g2188(.CO(n_83), .S(n_84), .A(in_7[0]), .B(n_50), .CI(n_54));
  ADDFX1 g2189(.CO(n_81), .S(n_82), .A(n_58), .B(n_60), .CI(n_30));
  ADDFX1 g2190(.CO(n_79), .S(n_80), .A(n_51), .B(n_43), .CI(n_67));
  ADDFX1 g2191(.CO(n_77), .S(n_78), .A(n_34), .B(n_28), .CI(n_38));
  ADDFX1 g2192(.CO(n_75), .S(n_76), .A(n_32), .B(n_62), .CI(n_40));
  ADDFX1 g2193(.CO(n_73), .S(n_74), .A(n_19), .B(n_29), .CI(n_27));
  ADDFX1 g2194(.CO(n_71), .S(n_72), .A(n_48), .B(n_56), .CI(n_36));
  ADDFX1 g2195(.CO(n_69), .S(n_70), .A(in_27[0]), .B(n_18), .CI(n_41));
  ADDFX1 g2196(.CO(n_67), .S(n_68), .A(in_21[1]), .B(n_24), .CI(in_18[1]));
  ADDFX1 g2197(.CO(n_65), .S(n_66), .A(n_23), .B(n_4), .CI(n_0));
  XNOR2X1 g2198(.Y(n_64), .A(n_25), .B(n_21));
  NAND3X1 g2199(.Y(n_63), .A(in_3[6]), .B(n_25), .C(n_21));
  ADDFX1 g2200(.CO(n_61), .S(n_62), .A(in_30[0]), .B(n_20), .CI(in_5[0]));
  ADDFX1 g2201(.CO(n_59), .S(n_60), .A(in_15[0]), .B(n_3), .CI(in_28[0]));
  ADDFX1 g2202(.CO(n_57), .S(n_58), .A(in_11[0]), .B(in_18[0]), .CI(n_14));
  ADDFX1 g2203(.CO(n_55), .S(n_56), .A(in_27[0]), .B(n_11), .CI(in_42[0]));
  ADDFX1 g2204(.CO(n_53), .S(n_54), .A(in_24[0]), .B(in_33), .CI(n_6));
  INVX1 g2205(.Y(n_52), .A(n_46));
  INVX1 g2206(.Y(n_51), .A(n_45));
  ADDFX1 g2207(.CO(n_49), .S(n_50), .A(in_13[0]), .B(in_32), .CI(n_8));
  ADDFX1 g2208(.CO(n_47), .S(n_48), .A(in_6[1]), .B(n_16), .CI(in_39[0]));
  ADDFX1 g2209(.CO(n_45), .S(n_46), .A(in_16[1]), .B(in_12[1]), .CI(in_7[1]));
  ADDFX1 g2210(.CO(n_43), .S(n_44), .A(in_17[1]), .B(n_7), .CI(in_5[1]));
  ADDFX1 g2211(.CO(n_41), .S(n_42), .A(n_9), .B(in_5[2]), .CI(n_2));
  ADDFX1 g2212(.CO(n_39), .S(n_40), .A(in_10[0]), .B(in_9[0]), .CI(in_21[0]));
  ADDFX1 g2213(.CO(n_37), .S(n_38), .A(in_34[0]), .B(in_37), .CI(in_41));
  ADDFX1 g2214(.CO(n_35), .S(n_36), .A(n_13), .B(in_36[1]), .CI(n_12));
  ADDFX1 g2215(.CO(n_33), .S(n_34), .A(in_19[0]), .B(n_15), .CI(in_39[0]));
  ADDFX1 g2216(.CO(n_31), .S(n_32), .A(in_16[0]), .B(in_17[0]), .CI(in_12[0]));
  ADDFX1 g2217(.CO(n_29), .S(n_30), .A(in_38[0]), .B(n_10), .CI(in_42[0]));
  ADDFX1 g2218(.CO(n_27), .S(n_28), .A(in_20[0]), .B(n_5), .CI(in_27[0]));
  XNOR2X1 g2219(.Y(n_26), .A(in_3[6]), .B(n_17));
  NAND2BX1 g2220(.Y(n_25), .AN(n_17), .B(in_3[6]));
  ADDHX1 g2221(.CO(n_23), .S(n_24), .A(in_19[0]), .B(in_23[1]));
  AO21XL g2222(.Y(n_22), .A0(n_1), .A1(in_3[5]), .B0(n_17));
  XNOR2X1 g2223(.Y(n_21), .A(in_3[6]), .B(in_2[7]));
  XOR2XL g2225(.Y(n_20), .A(in_31[0]), .B(in_40[0]));
  NOR2X1 g2226(.Y(n_19), .A(in_40[0]), .B(in_31[0]));
  NOR2X1 g2227(.Y(n_18), .A(in_38[0]), .B(in_15[0]));
  NOR2X1 g2228(.Y(n_17), .A(n_1), .B(in_3[5]));
  INVX1 g2229(.Y(n_16), .A(in_1[1]));
  INVX1 g2230(.Y(n_15), .A(in_25[0]));
  INVX1 g2231(.Y(n_14), .A(in_8[0]));
  INVX1 g2232(.Y(n_13), .A(in_29[1]));
  INVX1 g2233(.Y(n_12), .A(in_10[1]));
  INVX1 g2234(.Y(n_11), .A(in_26[1]));
  INVX1 g2235(.Y(n_10), .A(in_4[0]));
  INVX1 g2236(.Y(n_9), .A(in_34[0]));
  INVX1 g2238(.Y(n_8), .A(in_35[0]));
  INVX1 g2239(.Y(n_7), .A(in_9[1]));
  INVX1 g2240(.Y(n_6), .A(in_22[0]));
  INVX1 g2241(.Y(n_5), .A(in_14[0]));
  INVX1 g2242(.Y(n_4), .A(in_18[2]));
  INVX1 g2243(.Y(n_3), .A(in_0[0]));
  INVX1 g2244(.Y(n_2), .A(in_21[2]));
  INVX1 g2246(.Y(n_1), .A(in_27[0]));
  XOR2XL g2(.Y(n_0), .A(in_38[0]), .B(in_15[0]));
endmodule

module WALLACE_CSA_DUMMY_OP93_group_109834(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, out_0);
input  in_14, in_22, in_24, in_26;
input   [9:0] in_0;
input   [9:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [2:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [1:0] in_15;
input   [1:0] in_16;
input   [1:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [1:0] in_21;
input   [2:0] in_23;
input   [1:0] in_25;
input   [1:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [2:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [3:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [3:0] in_40;
input   [4:0] in_41;
input   [2:0] in_42;
input   [4:0] in_43;
output  [9:0] out_0;
wire  n_151, n_149, n_147, n_145, n_143, n_141, n_139, n_138, n_137, n_136, 
    n_135, n_134, n_133, n_131, n_130, n_129, n_128, n_127, n_126, n_125, 
    n_124, n_123, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1, n_0, in_26, in_24, in_22, in_14;
wire   [9:0] out_0;
wire   [3:0] in_40;
wire   [3:0] in_33;
wire   [4:0] in_43;
wire   [4:0] in_41;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_32;
wire   [4:0] in_28;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [1:0] in_36;
wire   [1:0] in_31;
wire   [1:0] in_29;
wire   [1:0] in_27;
wire   [1:0] in_25;
wire   [1:0] in_21;
wire   [1:0] in_17;
wire   [1:0] in_16;
wire   [1:0] in_15;
wire   [2:0] in_42;
wire   [2:0] in_37;
wire   [2:0] in_30;
wire   [2:0] in_23;
wire   [2:0] in_6;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [9:0] in_1;
wire   [9:0] in_0;
  INVX1 g4761(.Y(out_0[8]), .A(n_151));
  ADDFX1 g4762(.CO(out_0[9]), .S(n_151), .A(in_0[8]), .B(n_101), .CI(n_149));
  INVX1 g4763(.Y(n_149), .A(n_147));
  ADDFX1 g4764(.CO(n_147), .S(out_0[7]), .A(n_129), .B(n_112), .CI(n_145));
  ADDFX1 g4765(.CO(n_145), .S(out_0[6]), .A(n_133), .B(n_130), .CI(n_143));
  ADDFX1 g4766(.CO(n_143), .S(out_0[5]), .A(n_137), .B(n_134), .CI(n_141));
  ADDFX1 g4767(.CO(n_141), .S(out_0[4]), .A(n_135), .B(n_138), .CI(n_139));
  ADDFX1 g4768(.CO(n_139), .S(out_0[3]), .A(n_117), .B(n_131), .CI(n_136));
  ADDFX1 g4769(.CO(n_137), .S(n_138), .A(n_125), .B(n_128), .CI(in_0[4]));
  ADDFX1 g4770(.CO(n_135), .S(n_136), .A(n_123), .B(n_126), .CI(in_0[3]));
  ADDFX1 g4771(.CO(n_133), .S(n_134), .A(n_120), .B(n_127), .CI(in_0[5]));
  ADDFX1 g4772(.CO(n_131), .S(out_0[2]), .A(n_124), .B(n_121), .CI(n_118));
  ADDFX1 g4773(.CO(n_129), .S(n_130), .A(n_0), .B(n_119), .CI(in_0[6]));
  ADDFX1 g4774(.CO(n_127), .S(n_128), .A(n_115), .B(n_102), .CI(n_114));
  ADDFX1 g4775(.CO(n_125), .S(n_126), .A(n_116), .B(n_103), .CI(n_108));
  ADDFX1 g4776(.CO(n_123), .S(n_124), .A(n_95), .B(n_111), .CI(n_106));
  ADDFX1 g4777(.CO(n_121), .S(out_0[1]), .A(n_107), .B(n_97), .CI(n_105));
  ADDFX1 g4778(.CO(n_119), .S(n_120), .A(n_80), .B(in_1[5]), .CI(n_113));
  ADDFX1 g4779(.CO(n_117), .S(n_118), .A(n_109), .B(n_104), .CI(in_0[2]));
  ADDFX1 g4780(.CO(n_115), .S(n_116), .A(n_94), .B(n_100), .CI(n_110));
  ADDFX1 g4781(.CO(n_113), .S(n_114), .A(n_87), .B(n_99), .CI(in_1[4]));
  AO21XL g4782(.Y(n_112), .A0(n_96), .A1(in_0[7]), .B0(n_101));
  ADDFX1 g4783(.CO(n_110), .S(n_111), .A(n_89), .B(n_85), .CI(n_92));
  ADDFX1 g4784(.CO(n_108), .S(n_109), .A(n_82), .B(in_1[2]), .CI(n_90));
  ADDFX1 g4785(.CO(n_106), .S(n_107), .A(n_86), .B(n_93), .CI(n_76));
  ADDFX1 g4786(.CO(n_104), .S(n_105), .A(n_83), .B(n_91), .CI(in_0[1]));
  ADDFX1 g4787(.CO(n_102), .S(n_103), .A(n_78), .B(n_88), .CI(in_1[3]));
  NOR2X1 g4788(.Y(n_101), .A(n_96), .B(in_0[7]));
  ADDFX1 g4790(.CO(n_99), .S(n_100), .A(n_49), .B(n_72), .CI(n_81));
  ADDHX1 g4791(.CO(n_97), .S(out_0[0]), .A(n_77), .B(n_84));
  NOR2X1 g4792(.Y(n_96), .A(n_80), .B(in_1[6]));
  ADDFX1 g4794(.CO(n_94), .S(n_95), .A(n_62), .B(n_74), .CI(n_73));
  ADDFX1 g4795(.CO(n_92), .S(n_93), .A(n_54), .B(n_66), .CI(n_69));
  ADDFX1 g4796(.CO(n_90), .S(n_91), .A(n_63), .B(n_75), .CI(in_1[1]));
  ADDFX1 g4797(.CO(n_88), .S(n_89), .A(n_57), .B(n_70), .CI(n_59));
  XNOR2X1 g4798(.Y(n_87), .A(n_48), .B(n_79));
  ADDFX1 g4799(.CO(n_85), .S(n_86), .A(n_65), .B(n_71), .CI(n_60));
  ADDFX1 g4800(.CO(n_83), .S(n_84), .A(n_61), .B(n_67), .CI(in_0[0]));
  ADDFX1 g4801(.CO(n_81), .S(n_82), .A(n_52), .B(n_68), .CI(n_64));
  NAND2BX1 g4802(.Y(n_80), .AN(n_48), .B(n_79));
  ADDFX1 g4803(.CO(n_79), .S(n_78), .A(n_26), .B(n_56), .CI(n_58));
  ADDFX1 g4804(.CO(n_76), .S(n_77), .A(n_33), .B(n_55), .CI(in_1[0]));
  ADDFX1 g4805(.CO(n_74), .S(n_75), .A(n_39), .B(n_37), .CI(n_53));
  ADDFX1 g4806(.CO(n_72), .S(n_73), .A(n_38), .B(n_44), .CI(n_27));
  ADDFX1 g4807(.CO(n_70), .S(n_71), .A(n_18), .B(n_40), .CI(n_22));
  ADDFX1 g4808(.CO(n_68), .S(n_69), .A(n_32), .B(n_20), .CI(n_46));
  ADDFX1 g4809(.CO(n_66), .S(n_67), .A(n_43), .B(n_21), .CI(n_41));
  ADDFX1 g4810(.CO(n_64), .S(n_65), .A(in_10[1]), .B(n_16), .CI(n_42));
  ADDFX1 g4811(.CO(n_62), .S(n_63), .A(n_35), .B(n_25), .CI(n_31));
  ADDFX1 g4812(.CO(n_60), .S(n_61), .A(n_19), .B(n_17), .CI(n_23));
  ADDFX1 g4813(.CO(n_58), .S(n_59), .A(n_30), .B(n_34), .CI(n_24));
  ADDFX1 g4814(.CO(n_56), .S(n_57), .A(in_43[0]), .B(n_14), .CI(n_36));
  ADDFX1 g4815(.CO(n_54), .S(n_55), .A(in_2[0]), .B(in_12[0]), .CI(n_47));
  INVX1 g4816(.Y(n_53), .A(n_51));
  INVX1 g4817(.Y(n_52), .A(n_50));
  ADDFX1 g4818(.CO(n_50), .S(n_51), .A(in_12[1]), .B(n_15), .CI(in_2[1]));
  AO21X1 g4819(.Y(n_49), .A0(n_10), .A1(n_45), .B0(n_48));
  NOR2X1 g4820(.Y(n_48), .A(n_10), .B(n_45));
  ADDFX1 g4821(.CO(n_46), .S(n_47), .A(in_5[0]), .B(in_13[0]), .CI(in_33[0]));
  ADDFX1 g4822(.CO(n_45), .S(n_44), .A(n_12), .B(n_1), .CI(in_40[0]));
  ADDFX1 g4823(.CO(n_42), .S(n_43), .A(in_6[0]), .B(in_26), .CI(in_28[0]));
  ADDFX1 g4824(.CO(n_40), .S(n_41), .A(in_8[0]), .B(n_5), .CI(in_21[0]));
  ADDFX1 g4825(.CO(n_38), .S(n_39), .A(in_6[0]), .B(n_6), .CI(in_25[1]));
  ADDFX1 g4826(.CO(n_36), .S(n_37), .A(in_9[1]), .B(in_42[1]), .CI(n_11));
  ADDFX1 g4827(.CO(n_34), .S(n_35), .A(in_16[1]), .B(in_15[1]), .CI(in_37[1]));
  ADDFX1 g4828(.CO(n_32), .S(n_33), .A(in_10[0]), .B(in_14), .CI(n_8));
  INVX1 g4829(.Y(n_31), .A(n_29));
  INVX1 g4830(.Y(n_30), .A(n_28));
  ADDFX1 g4831(.CO(n_28), .S(n_29), .A(in_32[1]), .B(in_35[1]), .CI(in_38[1]));
  ADDFX1 g4832(.CO(n_26), .S(n_27), .A(in_23[2]), .B(in_33[0]), .CI(n_7));
  ADDFX1 g4833(.CO(n_24), .S(n_25), .A(in_5[1]), .B(in_27[1]), .CI(n_3));
  ADDFX1 g4834(.CO(n_22), .S(n_23), .A(in_24), .B(in_29[0]), .CI(in_40[0]));
  ADDFX1 g4835(.CO(n_20), .S(n_21), .A(in_22), .B(in_36[0]), .CI(n_9));
  ADDFX1 g4836(.CO(n_18), .S(n_19), .A(n_13), .B(in_31[0]), .CI(n_2));
  ADDFX1 g4837(.CO(n_16), .S(n_17), .A(in_17[0]), .B(n_4), .CI(in_43[0]));
  XNOR2X1 g4838(.Y(n_15), .A(in_30[1]), .B(in_17[0]));
  AND2XL g4839(.Y(n_14), .A(in_30[1]), .B(in_17[0]));
  INVX1 g4840(.Y(n_13), .A(in_4[0]));
  INVX1 g4841(.Y(n_12), .A(in_19[2]));
  INVX1 g4842(.Y(n_11), .A(in_20[1]));
  INVX1 g4843(.Y(n_10), .A(in_43[0]));
  INVX1 g4844(.Y(n_9), .A(in_39[0]));
  INVX1 g4845(.Y(n_8), .A(in_41[0]));
  INVX1 g4846(.Y(n_7), .A(in_10[2]));
  INVX1 g4847(.Y(n_6), .A(in_3[1]));
  INVX1 g4848(.Y(n_5), .A(in_11[0]));
  INVX1 g4849(.Y(n_4), .A(in_34[0]));
  INVX1 g4850(.Y(n_3), .A(in_18[1]));
  INVX1 g4851(.Y(n_2), .A(in_7[0]));
  INVX1 g4852(.Y(n_1), .A(in_28[0]));
  CLKXOR2X1 g2(.Y(n_0), .A(n_80), .B(in_1[6]));
endmodule

module WALLACE_CSA_DUMMY_OP95_group_109821(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, out_0);
input  in_22, in_32, in_33;
input   [4:0] in_0;
input   [4:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [4:0] in_19;
input   [1:0] in_20;
input   [1:0] in_21;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [1:0] in_27;
input   [1:0] in_28;
input   [4:0] in_29;
input   [1:0] in_30;
input   [4:0] in_31;
input   [4:0] in_34;
input   [1:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
output  [9:0] out_0;
wire  n_119, n_117, n_115, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, 
    n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, 
    n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, 
    n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
    n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
    n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, 
    n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
    n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
    n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_33, in_32, in_22;
wire   [9:0] out_0;
wire   [1:0] in_35;
wire   [1:0] in_30;
wire   [1:0] in_28;
wire   [1:0] in_27;
wire   [1:0] in_26;
wire   [1:0] in_21;
wire   [1:0] in_20;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_34;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_19;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3657(.Y(out_0[9]), .A(n_119));
  ADDFX1 g3658(.CO(n_119), .S(out_0[5]), .A(n_77), .B(n_109), .CI(n_117));
  ADDFX1 g3659(.CO(n_117), .S(out_0[4]), .A(n_110), .B(n_111), .CI(n_115));
  ADDFX1 g3660(.CO(n_115), .S(out_0[3]), .A(n_107), .B(n_112), .CI(n_113));
  ADDFX1 g3661(.CO(n_113), .S(out_0[2]), .A(n_99), .B(n_105), .CI(n_108));
  ADDFX1 g3662(.CO(n_111), .S(n_112), .A(n_96), .B(n_101), .CI(n_104));
  ADDFX1 g3663(.CO(n_109), .S(n_110), .A(n_78), .B(n_95), .CI(n_103));
  ADDFX1 g3664(.CO(n_107), .S(n_108), .A(n_91), .B(n_98), .CI(n_102));
  ADDFX1 g3665(.CO(n_105), .S(out_0[1]), .A(n_93), .B(n_92), .CI(n_100));
  ADDFX1 g3666(.CO(n_103), .S(n_104), .A(n_87), .B(n_89), .CI(n_97));
  ADDFX1 g3667(.CO(n_101), .S(n_102), .A(n_85), .B(n_83), .CI(n_90));
  ADDFX1 g3668(.CO(n_99), .S(n_100), .A(n_79), .B(n_86), .CI(n_84));
  ADDFX1 g3669(.CO(n_97), .S(n_98), .A(n_74), .B(n_82), .CI(n_88));
  ADDFX1 g3670(.CO(n_95), .S(n_96), .A(n_72), .B(n_76), .CI(n_81));
  ADDFX1 g3671(.CO(n_93), .S(out_0[0]), .A(n_71), .B(n_69), .CI(n_80));
  ADDFX1 g3672(.CO(n_91), .S(n_92), .A(n_68), .B(n_63), .CI(n_75));
  ADDFX1 g3673(.CO(n_89), .S(n_90), .A(n_57), .B(n_73), .CI(n_62));
  ADDFX1 g3674(.CO(n_87), .S(n_88), .A(n_54), .B(n_66), .CI(n_64));
  ADDFX1 g3675(.CO(n_85), .S(n_86), .A(n_70), .B(n_61), .CI(n_58));
  ADDFX1 g3676(.CO(n_83), .S(n_84), .A(n_55), .B(n_67), .CI(n_65));
  ADDFX1 g3677(.CO(n_81), .S(n_82), .A(n_50), .B(n_31), .CI(n_60));
  ADDFX1 g3678(.CO(n_79), .S(n_80), .A(n_47), .B(n_33), .CI(n_59));
  INVX1 g3679(.Y(n_78), .A(n_77));
  ADDFX1 g3680(.CO(n_77), .S(n_76), .A(n_7), .B(n_30), .CI(n_56));
  ADDFX1 g3681(.CO(n_74), .S(n_75), .A(n_39), .B(n_51), .CI(n_32));
  ADDFX1 g3682(.CO(n_72), .S(n_73), .A(n_34), .B(n_38), .CI(n_44));
  ADDFX1 g3683(.CO(n_70), .S(n_71), .A(in_16[0]), .B(n_41), .CI(n_37));
  ADDFX1 g3684(.CO(n_68), .S(n_69), .A(n_20), .B(n_43), .CI(n_53));
  ADDFX1 g3685(.CO(n_66), .S(n_67), .A(n_18), .B(n_40), .CI(n_36));
  ADDFX1 g3686(.CO(n_64), .S(n_65), .A(n_21), .B(n_46), .CI(n_24));
  ADDFX1 g3687(.CO(n_62), .S(n_63), .A(n_23), .B(n_35), .CI(n_45));
  ADDFX1 g3688(.CO(n_60), .S(n_61), .A(n_52), .B(n_48), .CI(n_26));
  ADDFX1 g3689(.CO(n_58), .S(n_59), .A(n_27), .B(n_49), .CI(n_25));
  ADDFX1 g3690(.CO(n_56), .S(n_57), .A(in_36[2]), .B(n_19), .CI(n_22));
  ADDFX1 g3691(.CO(n_54), .S(n_55), .A(in_17[1]), .B(in_2[1]), .CI(n_42));
  ADDFX1 g3692(.CO(n_52), .S(n_53), .A(in_15[0]), .B(n_2), .CI(n_14));
  ADDFX1 g3693(.CO(n_50), .S(n_51), .A(in_15[0]), .B(n_9), .CI(n_13));
  ADDFX1 g3694(.CO(n_48), .S(n_49), .A(in_4[0]), .B(in_35[0]), .CI(n_3));
  ADDFX1 g3695(.CO(n_46), .S(n_47), .A(in_6[0]), .B(in_33), .CI(in_9[0]));
  ADDFX1 g3696(.CO(n_44), .S(n_45), .A(in_7[1]), .B(n_11), .CI(n_6));
  ADDFX1 g3697(.CO(n_42), .S(n_43), .A(in_10[0]), .B(in_12[0]), .CI(in_13[0]));
  ADDFX1 g3698(.CO(n_40), .S(n_41), .A(in_2[0]), .B(n_4), .CI(in_30[0]));
  ADDFX1 g3699(.CO(n_38), .S(n_39), .A(in_6[1]), .B(in_12[0]), .CI(n_17));
  ADDFX1 g3700(.CO(n_36), .S(n_37), .A(in_26[0]), .B(in_22), .CI(in_27[0]));
  ADDFX1 g3701(.CO(n_34), .S(n_35), .A(in_4[0]), .B(n_8), .CI(n_15));
  ADDFX1 g3702(.CO(n_32), .S(n_33), .A(in_8[0]), .B(n_5), .CI(in_11[0]));
  INVX1 g3703(.Y(n_31), .A(n_29));
  INVX1 g3704(.Y(n_30), .A(n_28));
  ADDFX1 g3705(.CO(n_28), .S(n_29), .A(in_9[0]), .B(in_17[2]), .CI(in_2[2]));
  ADDFX1 g3706(.CO(n_26), .S(n_27), .A(in_5[0]), .B(n_10), .CI(in_28[0]));
  ADDFX1 g3707(.CO(n_24), .S(n_25), .A(in_32), .B(in_20[0]), .CI(n_12));
  ADDFX1 g3708(.CO(n_22), .S(n_23), .A(n_1), .B(in_5[1]), .CI(n_16));
  OAI2BB1X1 g3709(.Y(n_21), .A0N(in_21[1]), .A1N(in_18[1]), .B0(n_19));
  OAI2BB1X1 g3710(.Y(n_20), .A0N(in_18[0]), .A1N(in_17[0]), .B0(n_18));
  OR2X1 g3711(.Y(n_19), .A(in_21[1]), .B(in_18[1]));
  OR2X1 g3712(.Y(n_18), .A(in_18[0]), .B(in_17[0]));
  INVX1 g3713(.Y(n_17), .A(in_31[1]));
  INVX1 g3714(.Y(n_16), .A(in_29[1]));
  INVX1 g3715(.Y(n_15), .A(in_19[1]));
  INVX1 g3716(.Y(n_14), .A(in_24[0]));
  INVX1 g3717(.Y(n_13), .A(in_16[1]));
  INVX1 g3718(.Y(n_12), .A(in_34[0]));
  INVX1 g3719(.Y(n_11), .A(in_8[1]));
  INVX1 g3720(.Y(n_10), .A(in_14[0]));
  INVX1 g3721(.Y(n_9), .A(in_11[1]));
  INVX1 g3722(.Y(n_8), .A(in_0[1]));
  INVX1 g3723(.Y(n_7), .A(in_36[2]));
  INVX1 g3724(.Y(n_6), .A(in_37[1]));
  INVX1 g3725(.Y(n_5), .A(in_38[0]));
  INVX1 g3726(.Y(n_4), .A(in_3[0]));
  INVX1 g3727(.Y(n_3), .A(in_1[0]));
  INVX1 g3728(.Y(n_2), .A(in_23[0]));
  INVX1 g3729(.Y(n_1), .A(in_25[1]));
endmodule

module WALLACE_CSA_DUMMY_OP98_group_359290(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, out_0);
input  in_30, in_31, in_37, in_39, in_40, in_42, in_62;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [9:0] in_3;
input   [9:0] in_4;
input   [8:0] in_5;
input   [7:0] in_6;
input   [6:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [4:0] in_10;
input   [4:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [4:0] in_32;
input   [2:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_38;
input   [1:0] in_41;
input   [4:0] in_43;
input   [2:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [1:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [1:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [1:0] in_58;
input   [2:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [1:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [4:0] in_67;
input   [2:0] in_68;
input   [1:0] in_69;
input   [1:0] in_70;
input   [4:0] in_71;
input   [2:0] in_72;
input   [4:0] in_73;
input   [2:0] in_74;
output  [9:0] out_0;
wire  n_247, n_245, n_243, n_241, n_239, n_238, n_237, n_236, n_235, n_234, 
    n_233, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
    n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, 
    n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, 
    n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, 
    n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
    n_181, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, 
    n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, 
    n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, 
    n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, 
    n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
    n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, n_0, in_62, in_42, in_40, in_39, in_37, in_31, in_30;
wire   [9:0] out_0;
wire   [2:0] in_74;
wire   [2:0] in_72;
wire   [2:0] in_68;
wire   [2:0] in_59;
wire   [2:0] in_44;
wire   [2:0] in_33;
wire   [1:0] in_70;
wire   [1:0] in_69;
wire   [1:0] in_63;
wire   [1:0] in_61;
wire   [1:0] in_58;
wire   [1:0] in_55;
wire   [1:0] in_51;
wire   [1:0] in_50;
wire   [1:0] in_41;
wire   [1:0] in_38;
wire   [1:0] in_34;
wire   [1:0] in_25;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_7;
wire   [7:0] in_6;
wire   [8:0] in_5;
wire   [9:0] in_4;
wire   [9:0] in_3;
wire   [4:0] in_73;
wire   [4:0] in_71;
wire   [4:0] in_67;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_60;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_43;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_26;
wire   [4:0] in_11;
wire   [4:0] in_10;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g7954(.Y(out_0[9]), .A(n_247));
  ADDFX1 g7955(.CO(n_247), .S(out_0[7]), .A(n_102), .B(n_229), .CI(n_245));
  ADDFX1 g7956(.CO(n_245), .S(out_0[6]), .A(n_230), .B(n_235), .CI(n_243));
  ADDFX1 g7957(.CO(n_243), .S(out_0[5]), .A(n_237), .B(n_236), .CI(n_241));
  ADDFX1 g7958(.CO(n_241), .S(out_0[4]), .A(n_233), .B(n_238), .CI(n_239));
  ADDFX1 g7959(.CO(n_239), .S(out_0[3]), .A(n_223), .B(n_231), .CI(n_234));
  ADDFX1 g7960(.CO(n_237), .S(n_238), .A(n_218), .B(n_227), .CI(n_226));
  ADDFX1 g7961(.CO(n_235), .S(n_236), .A(n_217), .B(n_225), .CI(n_220));
  ADDFX1 g7962(.CO(n_233), .S(n_234), .A(n_212), .B(n_216), .CI(n_228));
  ADDFX1 g7963(.CO(n_231), .S(out_0[2]), .A(n_221), .B(n_210), .CI(n_224));
  ADDFX1 g7964(.CO(n_229), .S(n_230), .A(n_201), .B(n_99), .CI(n_219));
  ADDFX1 g7965(.CO(n_227), .S(n_228), .A(n_213), .B(n_208), .CI(n_209));
  ADDFX1 g7966(.CO(n_225), .S(n_226), .A(n_211), .B(n_206), .CI(n_215));
  ADDFX1 g7967(.CO(n_223), .S(n_224), .A(n_214), .B(n_203), .CI(n_196));
  ADDFX1 g7968(.CO(n_221), .S(out_0[1]), .A(n_179), .B(n_184), .CI(n_204));
  ADDFX1 g7969(.CO(n_219), .S(n_220), .A(n_205), .B(n_100), .CI(n_202));
  ADDFX1 g7970(.CO(n_217), .S(n_218), .A(n_193), .B(n_101), .CI(n_207));
  ADDFX1 g7971(.CO(n_215), .S(n_216), .A(n_194), .B(n_182), .CI(n_195));
  ADDFX1 g7972(.CO(n_213), .S(n_214), .A(n_199), .B(n_198), .CI(n_177));
  ADDFX1 g7973(.CO(n_211), .S(n_212), .A(n_186), .B(n_189), .CI(n_191));
  ADDFX1 g7974(.CO(n_209), .S(n_210), .A(n_190), .B(n_183), .CI(n_192));
  ADDFX1 g7975(.CO(n_207), .S(n_208), .A(n_197), .B(n_175), .CI(in_3[3]));
  ADDFX1 g7976(.CO(n_205), .S(n_206), .A(n_185), .B(n_188), .CI(n_181));
  ADDFX1 g7977(.CO(n_203), .S(n_204), .A(n_200), .B(n_178), .CI(n_170));
  ADDFX1 g7978(.CO(n_201), .S(n_202), .A(n_187), .B(n_34), .CI(in_3[5]));
  ADDFX1 g7979(.CO(n_199), .S(n_200), .A(n_150), .B(n_174), .CI(n_167));
  ADDFX1 g7980(.CO(n_197), .S(n_198), .A(n_159), .B(n_173), .CI(n_145));
  ADDFX1 g7981(.CO(n_195), .S(n_196), .A(n_166), .B(n_169), .CI(n_176));
  ADDFX1 g7982(.CO(n_193), .S(n_194), .A(n_163), .B(n_161), .CI(n_152));
  ADDFX1 g7983(.CO(n_191), .S(n_192), .A(n_164), .B(n_162), .CI(in_3[2]));
  ADDFX1 g7984(.CO(n_189), .S(n_190), .A(n_149), .B(n_148), .CI(n_171));
  ADDFX1 g7985(.CO(n_187), .S(n_188), .A(n_119), .B(n_157), .CI(n_151));
  ADDFX1 g7986(.CO(n_185), .S(n_186), .A(n_107), .B(n_155), .CI(n_147));
  ADDFX1 g7987(.CO(n_183), .S(n_184), .A(n_160), .B(n_153), .CI(n_172));
  ADDFX1 g7988(.CO(n_181), .S(n_182), .A(n_158), .B(n_165), .CI(in_4[3]));
  ADDFX1 g7989(.CO(n_179), .S(out_0[0]), .A(n_168), .B(n_144), .CI(n_154));
  ADDFX1 g7990(.CO(n_177), .S(n_178), .A(n_128), .B(n_143), .CI(n_146));
  ADDFX1 g7991(.CO(n_175), .S(n_176), .A(n_127), .B(n_156), .CI(in_4[2]));
  ADDFX1 g7992(.CO(n_173), .S(n_174), .A(n_140), .B(n_138), .CI(n_115));
  ADDFX1 g7993(.CO(n_171), .S(n_172), .A(n_122), .B(n_135), .CI(in_4[1]));
  ADDFX1 g7994(.CO(n_169), .S(n_170), .A(n_142), .B(n_130), .CI(in_3[1]));
  ADDFX1 g7995(.CO(n_167), .S(n_168), .A(n_116), .B(n_132), .CI(n_136));
  ADDFX1 g7996(.CO(n_165), .S(n_166), .A(n_141), .B(n_129), .CI(in_6[2]));
  ADDFX1 g7997(.CO(n_163), .S(n_164), .A(n_137), .B(n_110), .CI(n_112));
  ADDFX1 g7998(.CO(n_161), .S(n_162), .A(n_118), .B(n_121), .CI(n_108));
  ADDFX1 g7999(.CO(n_159), .S(n_160), .A(n_114), .B(n_134), .CI(n_103));
  ADDFX1 g8000(.CO(n_157), .S(n_158), .A(n_109), .B(n_111), .CI(n_117));
  ADDFX1 g8001(.CO(n_155), .S(n_156), .A(n_139), .B(n_113), .CI(n_105));
  ADDFX1 g8002(.CO(n_153), .S(n_154), .A(n_124), .B(n_126), .CI(in_3[0]));
  ADDFX1 g8003(.CO(n_151), .S(n_152), .A(n_120), .B(n_6), .CI(in_5[3]));
  ADDFX1 g8004(.CO(n_149), .S(n_150), .A(n_106), .B(n_123), .CI(n_125));
  ADDFX1 g8005(.CO(n_147), .S(n_148), .A(n_84), .B(n_133), .CI(in_5[2]));
  ADDFX1 g8006(.CO(n_145), .S(n_146), .A(n_131), .B(in_6[1]), .CI(in_5[1]));
  ADDFX1 g8007(.CO(n_143), .S(n_144), .A(n_72), .B(n_104), .CI(in_4[0]));
  ADDFX1 g8008(.CO(n_141), .S(n_142), .A(n_81), .B(n_98), .CI(n_56));
  ADDFX1 g8009(.CO(n_139), .S(n_140), .A(n_65), .B(n_91), .CI(n_63));
  ADDFX1 g8010(.CO(n_137), .S(n_138), .A(n_85), .B(n_37), .CI(n_35));
  ADDFX1 g8011(.CO(n_135), .S(n_136), .A(n_54), .B(n_82), .CI(in_6[0]));
  ADDFX1 g8012(.CO(n_133), .S(n_134), .A(n_89), .B(n_53), .CI(n_69));
  ADDFX1 g8013(.CO(n_131), .S(n_132), .A(n_70), .B(n_38), .CI(n_36));
  ADDFX1 g8014(.CO(n_129), .S(n_130), .A(n_96), .B(n_44), .CI(n_68));
  ADDFX1 g8015(.CO(n_127), .S(n_128), .A(n_88), .B(n_71), .CI(n_52));
  ADDFX1 g8016(.CO(n_125), .S(n_126), .A(n_50), .B(in_5[0]), .CI(n_86));
  ADDFX1 g8017(.CO(n_123), .S(n_124), .A(n_90), .B(n_74), .CI(n_92));
  ADDFX1 g8018(.CO(n_121), .S(n_122), .A(n_40), .B(n_80), .CI(n_48));
  ADDFX1 g8019(.CO(n_119), .S(n_120), .A(in_16[1]), .B(n_75), .CI(n_83));
  ADDFX1 g8020(.CO(n_117), .S(n_118), .A(n_97), .B(n_87), .CI(n_47));
  ADDFX1 g8021(.CO(n_115), .S(n_116), .A(n_94), .B(n_62), .CI(n_64));
  ADDFX1 g8022(.CO(n_113), .S(n_114), .A(n_73), .B(n_49), .CI(n_45));
  ADDFX1 g8023(.CO(n_111), .S(n_112), .A(n_43), .B(n_55), .CI(n_39));
  ADDFX1 g8024(.CO(n_109), .S(n_110), .A(n_16), .B(n_95), .CI(n_79));
  ADDFX1 g8025(.CO(n_107), .S(n_108), .A(n_76), .B(n_67), .CI(n_51));
  ADDFX1 g8026(.CO(n_105), .S(n_106), .A(n_61), .B(n_77), .CI(n_93));
  ADDFX1 g8027(.CO(n_103), .S(n_104), .A(n_78), .B(n_66), .CI(n_46));
  OAI22X1 g8028(.Y(n_102), .A0(n_33), .A1(n_31), .B0(in_4[6]), .B1(in_3[6]));
  ADDFX1 g8029(.CO(n_100), .S(n_101), .A(n_32), .B(in_4[4]), .CI(in_3[4]));
  XOR2XL g8030(.Y(n_99), .A(n_33), .B(n_31));
  ADDFX1 g8031(.CO(n_97), .S(n_98), .A(n_0), .B(in_74[1]), .CI(n_3));
  ADDFX1 g8032(.CO(n_95), .S(n_96), .A(in_41[1]), .B(in_44[1]), .CI(n_13));
  ADDFX1 g8033(.CO(n_93), .S(n_94), .A(in_28[0]), .B(in_29[0]), .CI(n_4));
  ADDFX1 g8034(.CO(n_91), .S(n_92), .A(in_24[0]), .B(in_17[0]), .CI(in_58[0]));
  ADDFX1 g8035(.CO(n_89), .S(n_90), .A(in_37), .B(n_18), .CI(in_48[0]));
  ADDFX1 g8036(.CO(n_87), .S(n_88), .A(in_9[1]), .B(in_68[0]), .CI(in_59[0]));
  ADDFX1 g8037(.CO(n_85), .S(n_86), .A(in_26[0]), .B(n_17), .CI(in_62));
  ADDFX1 g8038(.CO(n_83), .S(n_84), .A(n_15), .B(n_26), .CI(in_16[2]));
  ADDFX1 g8039(.CO(n_81), .S(n_82), .A(in_40), .B(in_51[0]), .CI(in_59[0]));
  INVX1 g8040(.Y(n_80), .A(n_60));
  INVX1 g8041(.Y(n_79), .A(n_59));
  INVX1 g8042(.Y(n_78), .A(n_58));
  INVX1 g8043(.Y(n_77), .A(n_57));
  INVX1 g8044(.Y(n_76), .A(n_42));
  INVX1 g8045(.Y(n_75), .A(n_41));
  ADDFX1 g8046(.CO(n_73), .S(n_74), .A(in_55[0]), .B(n_5), .CI(n_12));
  ADDFX1 g8047(.CO(n_71), .S(n_72), .A(in_33[0]), .B(in_27[0]), .CI(in_16[0]));
  ADDFX1 g8048(.CO(n_69), .S(n_70), .A(in_46[0]), .B(n_8), .CI(n_23));
  ADDFX1 g8049(.CO(n_67), .S(n_68), .A(n_25), .B(n_7), .CI(in_16[1]));
  ADDFX1 g8050(.CO(n_65), .S(n_66), .A(in_12[0]), .B(n_19), .CI(in_61[0]));
  ADDFX1 g8051(.CO(n_63), .S(n_64), .A(in_21[0]), .B(in_34[0]), .CI(n_10));
  ADDFX1 g8052(.CO(n_61), .S(n_62), .A(in_25[0]), .B(in_30), .CI(n_27));
  ADDFX1 g8053(.CO(n_59), .S(n_60), .A(in_7[1]), .B(in_12[1]), .CI(in_71[1]));
  ADDFX1 g8054(.CO(n_57), .S(n_58), .A(in_14[0]), .B(in_18[0]), .CI(in_19[0]));
  ADDFX1 g8055(.CO(n_55), .S(n_56), .A(in_38[1]), .B(n_21), .CI(n_28));
  ADDFX1 g8056(.CO(n_53), .S(n_54), .A(in_69[0]), .B(in_39), .CI(n_11));
  ADDFX1 g8057(.CO(n_51), .S(n_52), .A(n_1), .B(in_21[1]), .CI(in_28[1]));
  ADDFX1 g8058(.CO(n_49), .S(n_50), .A(in_22[0]), .B(in_50[0]), .CI(n_22));
  ADDFX1 g8059(.CO(n_47), .S(n_48), .A(in_63[1]), .B(n_2), .CI(n_14));
  ADDFX1 g8060(.CO(n_45), .S(n_46), .A(in_15[0]), .B(in_31), .CI(in_20[0]));
  ADDFX1 g8061(.CO(n_43), .S(n_44), .A(in_33[0]), .B(n_20), .CI(n_29));
  ADDFX1 g8062(.CO(n_41), .S(n_42), .A(in_46[0]), .B(in_35[2]), .CI(in_48[0]));
  ADDFX1 g8063(.CO(n_39), .S(n_40), .A(in_17[0]), .B(n_24), .CI(in_72[1]));
  ADDFX1 g8064(.CO(n_37), .S(n_38), .A(in_23[0]), .B(in_42), .CI(n_9));
  ADDFX1 g8065(.CO(n_35), .S(n_36), .A(in_13[0]), .B(in_68[0]), .CI(in_70[0]));
  XOR2XL g8066(.Y(n_34), .A(n_30), .B(in_4[5]));
  NAND2X1 g8067(.Y(n_33), .A(n_30), .B(in_4[5]));
  OAI21X1 g8068(.Y(n_32), .A0(in_16[1]), .A1(in_5[4]), .B0(n_30));
  XNOR2X1 g8069(.Y(n_31), .A(in_4[6]), .B(in_3[6]));
  NAND2X1 g8070(.Y(n_30), .A(in_16[1]), .B(in_5[4]));
  INVX1 g8071(.Y(n_29), .A(in_49[1]));
  INVX1 g8072(.Y(n_28), .A(in_57[1]));
  INVX1 g8073(.Y(n_27), .A(in_52[0]));
  INVX1 g8074(.Y(n_26), .A(in_28[2]));
  INVX1 g8075(.Y(n_25), .A(in_15[1]));
  INVX1 g8076(.Y(n_24), .A(in_67[1]));
  INVX1 g8077(.Y(n_23), .A(in_10[0]));
  INVX1 g8078(.Y(n_22), .A(in_11[0]));
  INVX1 g8079(.Y(n_21), .A(in_1[1]));
  INVX1 g8080(.Y(n_20), .A(in_32[1]));
  INVX1 g8081(.Y(n_19), .A(in_54[0]));
  INVX1 g8082(.Y(n_18), .A(in_2[0]));
  INVX1 g8083(.Y(n_17), .A(in_43[0]));
  INVX1 g8084(.Y(n_16), .A(in_21[2]));
  INVX1 g8085(.Y(n_15), .A(in_26[0]));
  INVX1 g8086(.Y(n_14), .A(in_65[1]));
  INVX1 g8087(.Y(n_13), .A(in_56[1]));
  INVX1 g8088(.Y(n_12), .A(in_66[0]));
  INVX1 g8089(.Y(n_11), .A(in_73[0]));
  INVX1 g8090(.Y(n_10), .A(in_47[0]));
  INVX1 g8091(.Y(n_9), .A(in_45[0]));
  INVX1 g8092(.Y(n_8), .A(in_64[0]));
  INVX1 g8093(.Y(n_7), .A(in_24[1]));
  INVX1 g8094(.Y(n_6), .A(in_6[3]));
  INVX1 g8095(.Y(n_5), .A(in_36[0]));
  INVX1 g8096(.Y(n_4), .A(in_0[0]));
  INVX1 g8097(.Y(n_3), .A(in_8[1]));
  INVX1 g8098(.Y(n_2), .A(in_53[1]));
  INVX1 g8099(.Y(n_1), .A(in_27[1]));
  INVX1 g8100(.Y(n_0), .A(in_60[1]));
endmodule

module WALLACE_CSA_DUMMY_OP99_group_106220(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88, in_89, in_90
    , in_91, in_92, out_0);
input  in_78, in_79, in_80, in_81, in_92;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [9:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [1:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [4:0] in_45;
input   [1:0] in_46;
input   [4:0] in_47;
input   [2:0] in_48;
input   [1:0] in_49;
input   [4:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [1:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [4:0] in_60;
input   [4:0] in_61;
input   [4:0] in_62;
input   [2:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [4:0] in_67;
input   [4:0] in_68;
input   [2:0] in_69;
input   [1:0] in_70;
input   [1:0] in_71;
input   [1:0] in_72;
input   [4:0] in_73;
input   [4:0] in_74;
input   [4:0] in_75;
input   [1:0] in_76;
input   [4:0] in_77;
input   [4:0] in_82;
input   [4:0] in_83;
input   [2:0] in_84;
input   [4:0] in_85;
input   [4:0] in_86;
input   [1:0] in_87;
input   [4:0] in_88;
input   [2:0] in_89;
input   [4:0] in_90;
input   [1:0] in_91;
output  [9:0] out_0;
wire  n_301, n_298, n_296, n_294, n_293, n_292, n_290, n_289, n_288, n_287, 
    n_286, n_285, n_284, n_283, n_282, n_280, n_279, n_278, n_277, n_276, 
    n_275, n_274, n_273, n_272, n_270, n_269, n_268, n_267, n_266, n_265, 
    n_264, n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, 
    n_244, n_243, n_242, n_240, n_239, n_238, n_237, n_236, n_235, n_234, 
    n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, 
    n_223, n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, 
    n_213, n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, 
    n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 
    n_193, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, 
    n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, 
    n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, 
    n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, 
    n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, 
    n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, 
    n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, 
    n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
    n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_92, in_81, in_80, in_79, in_78;
wire   [9:0] out_0;
wire   [1:0] in_91;
wire   [1:0] in_87;
wire   [1:0] in_76;
wire   [1:0] in_72;
wire   [1:0] in_71;
wire   [1:0] in_70;
wire   [1:0] in_56;
wire   [1:0] in_51;
wire   [1:0] in_49;
wire   [1:0] in_46;
wire   [1:0] in_39;
wire   [1:0] in_37;
wire   [1:0] in_36;
wire   [1:0] in_34;
wire   [1:0] in_33;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [9:0] in_3;
wire   [4:0] in_90;
wire   [4:0] in_88;
wire   [4:0] in_86;
wire   [4:0] in_85;
wire   [4:0] in_83;
wire   [4:0] in_82;
wire   [4:0] in_77;
wire   [4:0] in_75;
wire   [4:0] in_74;
wire   [4:0] in_73;
wire   [4:0] in_68;
wire   [4:0] in_67;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_62;
wire   [4:0] in_61;
wire   [4:0] in_60;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_50;
wire   [4:0] in_47;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_89;
wire   [2:0] in_84;
wire   [2:0] in_69;
wire   [2:0] in_63;
wire   [2:0] in_48;
wire   [2:0] in_0;
  OAI21XL g9260(.Y(out_0[9]), .A0(n_217), .A1(n_301), .B0(n_224));
  XNOR2X1 g9261(.Y(out_0[8]), .A(n_225), .B(n_301));
  ADDFX1 g9262(.CO(n_301), .S(out_0[7]), .A(n_216), .B(n_286), .CI(n_298));
  ADDFX1 g9263(.CO(n_298), .S(out_0[6]), .A(n_292), .B(n_287), .CI(n_296));
  ADDFX1 g9264(.CO(n_296), .S(out_0[5]), .A(n_288), .B(n_293), .CI(n_294));
  ADDFX1 g9265(.CO(n_294), .S(out_0[4]), .A(n_282), .B(n_289), .CI(n_290));
  ADDFX1 g9266(.CO(n_292), .S(n_293), .A(n_255), .B(n_284), .CI(n_279));
  ADDFX1 g9267(.CO(n_290), .S(out_0[3]), .A(n_272), .B(n_280), .CI(n_283));
  ADDFX1 g9268(.CO(n_288), .S(n_289), .A(n_274), .B(n_268), .CI(n_285));
  ADDFX1 g9269(.CO(n_286), .S(n_287), .A(n_254), .B(n_278), .CI(n_187));
  ADDFX1 g9270(.CO(n_284), .S(n_285), .A(n_262), .B(n_267), .CI(n_277));
  ADDFX1 g9271(.CO(n_282), .S(n_283), .A(n_275), .B(n_258), .CI(n_269));
  ADDFX1 g9272(.CO(n_280), .S(out_0[2]), .A(n_273), .B(n_270), .CI(n_259));
  ADDFX1 g9273(.CO(n_278), .S(n_279), .A(n_266), .B(in_3[5]), .CI(n_276));
  ADDFX1 g9274(.CO(n_276), .S(n_277), .A(n_249), .B(n_264), .CI(in_3[4]));
  ADDFX1 g9275(.CO(n_274), .S(n_275), .A(n_265), .B(n_260), .CI(n_263));
  ADDFX1 g9276(.CO(n_272), .S(n_273), .A(n_256), .B(n_261), .CI(n_253));
  ADDFX1 g9277(.CO(n_270), .S(out_0[1]), .A(n_257), .B(n_240), .CI(n_239));
  ADDFX1 g9278(.CO(n_268), .S(n_269), .A(n_242), .B(n_252), .CI(in_3[3]));
  ADDFX1 g9279(.CO(n_266), .S(n_267), .A(n_231), .B(n_246), .CI(n_236));
  ADDFX1 g9280(.CO(n_264), .S(n_265), .A(n_227), .B(n_234), .CI(n_250));
  ADDFX1 g9281(.CO(n_262), .S(n_263), .A(n_247), .B(n_232), .CI(n_237));
  ADDFX1 g9282(.CO(n_260), .S(n_261), .A(n_212), .B(n_251), .CI(n_228));
  ADDFX1 g9283(.CO(n_258), .S(n_259), .A(n_243), .B(n_238), .CI(in_3[2]));
  ADDFX1 g9284(.CO(n_256), .S(n_257), .A(n_210), .B(n_229), .CI(n_245));
  ADDFX1 g9285(.CO(n_254), .S(n_255), .A(n_181), .B(n_230), .CI(n_248));
  ADDFX1 g9286(.CO(n_252), .S(n_253), .A(n_235), .B(n_233), .CI(n_244));
  ADDFX1 g9287(.CO(n_250), .S(n_251), .A(n_153), .B(n_219), .CI(n_222));
  ADDFX1 g9288(.CO(n_248), .S(n_249), .A(n_190), .B(n_188), .CI(n_226));
  ADDFX1 g9289(.CO(n_246), .S(n_247), .A(n_218), .B(n_191), .CI(n_199));
  ADDFX1 g9290(.CO(n_244), .S(n_245), .A(n_223), .B(n_203), .CI(n_220));
  ADDFX1 g9291(.CO(n_242), .S(n_243), .A(n_194), .B(n_215), .CI(n_205));
  ADDFX1 g9292(.CO(n_240), .S(out_0[0]), .A(n_221), .B(n_211), .CI(in_3[0]));
  ADDFX1 g9293(.CO(n_238), .S(n_239), .A(n_195), .B(n_213), .CI(in_3[1]));
  ADDFX1 g9294(.CO(n_236), .S(n_237), .A(n_208), .B(n_204), .CI(n_189));
  ADDFX1 g9295(.CO(n_234), .S(n_235), .A(n_207), .B(n_202), .CI(n_200));
  ADDFX1 g9296(.CO(n_232), .S(n_233), .A(n_193), .B(n_196), .CI(n_209));
  ADDFX1 g9297(.CO(n_230), .S(n_231), .A(n_141), .B(n_176), .CI(n_198));
  ADDFX1 g9298(.CO(n_228), .S(n_229), .A(n_185), .B(n_201), .CI(n_197));
  ADDFX1 g9299(.CO(n_226), .S(n_227), .A(n_206), .B(n_192), .CI(n_214));
  NAND2BX1 g9300(.Y(n_225), .AN(n_217), .B(n_224));
  OAI2BB1X1 g9301(.Y(n_224), .A0N(n_1), .A1N(in_3[7]), .B0(in_3[8]));
  ADDFX1 g9302(.CO(n_222), .S(n_223), .A(n_125), .B(n_178), .CI(n_179));
  ADDFX1 g9303(.CO(n_220), .S(n_221), .A(n_140), .B(n_180), .CI(n_157));
  ADDFX1 g9304(.CO(n_218), .S(n_219), .A(n_177), .B(n_158), .CI(n_150));
  NOR3BX1 g9305(.Y(n_217), .AN(in_3[7]), .B(n_184), .C(in_3[8]));
  MX2XL g9306(.Y(n_216), .A(n_1), .B(n_184), .S0(in_3[7]));
  ADDFX1 g9307(.CO(n_214), .S(n_215), .A(n_144), .B(n_167), .CI(n_172));
  ADDFX1 g9308(.CO(n_212), .S(n_213), .A(n_146), .B(n_151), .CI(n_183));
  ADDFX1 g9309(.CO(n_210), .S(n_211), .A(n_171), .B(n_136), .CI(n_186));
  ADDFX1 g9311(.CO(n_208), .S(n_209), .A(n_165), .B(n_155), .CI(n_174));
  ADDFX1 g9312(.CO(n_206), .S(n_207), .A(n_147), .B(n_89), .CI(n_160));
  ADDFX1 g9313(.CO(n_204), .S(n_205), .A(n_134), .B(n_145), .CI(n_182));
  ADDFX1 g9314(.CO(n_202), .S(n_203), .A(n_148), .B(n_135), .CI(n_163));
  ADDFX1 g9315(.CO(n_200), .S(n_201), .A(n_139), .B(n_138), .CI(n_156));
  ADDFX1 g9316(.CO(n_198), .S(n_199), .A(n_143), .B(n_166), .CI(n_43));
  ADDFX1 g9317(.CO(n_196), .S(n_197), .A(n_170), .B(n_159), .CI(n_168));
  ADDFX1 g9318(.CO(n_194), .S(n_195), .A(n_161), .B(n_175), .CI(n_173));
  ADDFX1 g9319(.CO(n_192), .S(n_193), .A(n_124), .B(n_137), .CI(n_162));
  ADDFX1 g9320(.CO(n_190), .S(n_191), .A(n_154), .B(n_164), .CI(n_130));
  ADDFX1 g9321(.CO(n_188), .S(n_189), .A(n_133), .B(n_152), .CI(n_142));
  OAI2BB1X1 g9322(.Y(n_187), .A0N(n_149), .A1N(in_3[6]), .B0(n_1));
  ADDFX1 g9323(.CO(n_185), .S(n_186), .A(n_85), .B(n_127), .CI(n_169));
  INVX1 g9324(.Y(n_1), .A(n_184));
  NOR2X1 g9325(.Y(n_184), .A(n_149), .B(in_3[6]));
  ADDFX1 g9326(.CO(n_182), .S(n_183), .A(n_49), .B(n_109), .CI(n_126));
  INVX1 g9327(.Y(n_181), .A(n_149));
  ADDFX1 g9328(.CO(n_179), .S(n_180), .A(n_69), .B(n_103), .CI(n_47));
  ADDFX1 g9329(.CO(n_177), .S(n_178), .A(n_68), .B(n_112), .CI(n_100));
  OAI21X1 g9330(.Y(n_176), .A0(n_129), .A1(n_97), .B0(n_149));
  ADDFX1 g9331(.CO(n_174), .S(n_175), .A(n_99), .B(n_81), .CI(n_121));
  ADDFX1 g9332(.CO(n_172), .S(n_173), .A(n_123), .B(n_79), .CI(n_111));
  ADDFX1 g9333(.CO(n_170), .S(n_171), .A(n_67), .B(n_71), .CI(n_101));
  ADDFX1 g9334(.CO(n_168), .S(n_169), .A(n_91), .B(n_105), .CI(n_59));
  ADDFX1 g9335(.CO(n_166), .S(n_167), .A(n_74), .B(n_92), .CI(n_110));
  ADDFX1 g9336(.CO(n_164), .S(n_165), .A(n_44), .B(n_120), .CI(n_80));
  ADDFX1 g9337(.CO(n_162), .S(n_163), .A(n_46), .B(n_104), .CI(n_95));
  ADDFX1 g9338(.CO(n_160), .S(n_161), .A(n_50), .B(n_58), .CI(n_66));
  ADDFX1 g9339(.CO(n_158), .S(n_159), .A(n_102), .B(n_106), .CI(in_16[1]));
  ADDFX1 g9340(.CO(n_156), .S(n_157), .A(n_113), .B(n_53), .CI(n_96));
  ADDFX1 g9341(.CO(n_154), .S(n_155), .A(n_122), .B(n_114), .CI(n_98));
  ADDFX1 g9342(.CO(n_152), .S(n_153), .A(n_48), .B(n_108), .CI(n_73));
  ADDFX1 g9343(.CO(n_150), .S(n_151), .A(n_45), .B(n_93), .CI(n_115));
  NAND2X1 g9344(.Y(n_149), .A(n_129), .B(n_97));
  ADDFX1 g9345(.CO(n_147), .S(n_148), .A(n_52), .B(n_90), .CI(n_76));
  ADDFX1 g9346(.CO(n_145), .S(n_146), .A(n_55), .B(n_75), .CI(n_84));
  ADDFX1 g9347(.CO(n_143), .S(n_144), .A(n_41), .B(n_78), .CI(n_54));
  ADDFX1 g9348(.CO(n_141), .S(n_142), .A(n_94), .B(n_72), .CI(n_88));
  ADDFX1 g9349(.CO(n_139), .S(n_140), .A(in_28[0]), .B(n_107), .CI(n_61));
  ADDFX1 g9350(.CO(n_137), .S(n_138), .A(n_62), .B(n_60), .CI(n_70));
  ADDFX1 g9351(.CO(n_135), .S(n_136), .A(n_51), .B(n_77), .CI(n_63));
  INVX1 g9352(.Y(n_134), .A(n_132));
  INVX1 g9353(.Y(n_133), .A(n_131));
  ADDFX1 g9354(.CO(n_131), .S(n_132), .A(n_65), .B(n_87), .CI(n_57));
  INVX1 g9355(.Y(n_130), .A(n_128));
  ADDFX1 g9356(.CO(n_129), .S(n_128), .A(in_60[0]), .B(n_86), .CI(n_64));
  ADDFX1 g9357(.CO(n_126), .S(n_127), .A(n_39), .B(in_7[0]), .CI(in_15[0]));
  ADDFX1 g9358(.CO(n_124), .S(n_125), .A(n_0), .B(n_42), .CI(in_13[1]));
  INVX1 g9359(.Y(n_123), .A(n_119));
  INVX1 g9360(.Y(n_122), .A(n_118));
  INVX1 g9361(.Y(n_121), .A(n_117));
  INVX1 g9362(.Y(n_120), .A(n_116));
  ADDFX1 g9363(.CO(n_118), .S(n_119), .A(in_44[1]), .B(in_86[1]), .CI(in_64[1]));
  ADDFX1 g9364(.CO(n_116), .S(n_117), .A(in_40[1]), .B(in_55[1]), .CI(in_88[1]));
  ADDFX1 g9365(.CO(n_114), .S(n_115), .A(in_48[1]), .B(n_28), .CI(n_21));
  ADDFX1 g9366(.CO(n_112), .S(n_113), .A(in_9[0]), .B(in_74[0]), .CI(in_91[0]));
  ADDFX1 g9367(.CO(n_110), .S(n_111), .A(in_18[1]), .B(in_21[1]), .CI(n_20));
  ADDFX1 g9368(.CO(n_108), .S(n_109), .A(in_28[1]), .B(in_7[1]), .CI(in_17[1]));
  ADDFX1 g9369(.CO(n_106), .S(n_107), .A(in_34[0]), .B(in_72[0]), .CI(in_92));
  ADDFX1 g9370(.CO(n_104), .S(n_105), .A(in_56[0]), .B(in_81), .CI(n_27));
  ADDFX1 g9371(.CO(n_102), .S(n_103), .A(in_63[0]), .B(n_37), .CI(n_29));
  ADDFX1 g9372(.CO(n_100), .S(n_101), .A(in_75[0]), .B(in_80), .CI(n_10));
  ADDFX1 g9373(.CO(n_98), .S(n_99), .A(n_5), .B(n_14), .CI(in_91[0]));
  OAI2BB1X1 g9374(.Y(n_97), .A0N(in_45[0]), .A1N(n_38), .B0(n_40));
  INVX1 g9375(.Y(n_96), .A(n_83));
  INVX1 g9376(.Y(n_95), .A(n_82));
  INVX1 g9377(.Y(n_94), .A(n_56));
  ADDFX1 g9378(.CO(n_92), .S(n_93), .A(in_14[1]), .B(n_9), .CI(in_89[1]));
  ADDFX1 g9379(.CO(n_90), .S(n_91), .A(in_12[0]), .B(in_70[0]), .CI(n_17));
  ADDFX1 g9380(.CO(n_88), .S(n_89), .A(in_60[0]), .B(n_34), .CI(in_14[2]));
  ADDFX1 g9381(.CO(n_86), .S(n_87), .A(in_50[0]), .B(in_58[2]), .CI(in_74[0]));
  ADDFX1 g9382(.CO(n_84), .S(n_85), .A(in_29[0]), .B(in_17[0]), .CI(in_23[0]));
  ADDFX1 g9383(.CO(n_82), .S(n_83), .A(in_52[0]), .B(in_57[0]), .CI(in_67[0]));
  ADDFX1 g9384(.CO(n_80), .S(n_81), .A(n_6), .B(in_27[1]), .CI(n_36));
  ADDFX1 g9385(.CO(n_78), .S(n_79), .A(n_16), .B(n_33), .CI(in_70[0]));
  ADDFX1 g9386(.CO(n_76), .S(n_77), .A(in_62[0]), .B(in_76[0]), .CI(n_7));
  ADDFX1 g9387(.CO(n_74), .S(n_75), .A(in_45[0]), .B(n_12), .CI(in_63[0]));
  ADDFX1 g9388(.CO(n_72), .S(n_73), .A(n_23), .B(n_35), .CI(in_7[2]));
  ADDFX1 g9389(.CO(n_70), .S(n_71), .A(in_5[0]), .B(in_37[0]), .CI(in_87[0]));
  ADDFX1 g9390(.CO(n_68), .S(n_69), .A(in_22[0]), .B(n_11), .CI(in_51[0]));
  ADDFX1 g9391(.CO(n_66), .S(n_67), .A(in_16[0]), .B(n_2), .CI(in_79));
  ADDFX1 g9392(.CO(n_64), .S(n_65), .A(in_12[0]), .B(in_17[2]), .CI(in_22[0]));
  ADDFX1 g9393(.CO(n_62), .S(n_63), .A(n_32), .B(n_13), .CI(in_45[0]));
  ADDFX1 g9394(.CO(n_60), .S(n_61), .A(in_6[0]), .B(in_46[0]), .CI(in_50[0]));
  ADDFX1 g9395(.CO(n_58), .S(n_59), .A(in_33[0]), .B(in_36[0]), .CI(in_49[0]));
  ADDFX1 g9396(.CO(n_56), .S(n_57), .A(in_9[0]), .B(in_59[2]), .CI(in_75[0]));
  ADDFX1 g9397(.CO(n_54), .S(n_55), .A(in_0[1]), .B(n_26), .CI(in_71[1]));
  ADDFX1 g9398(.CO(n_52), .S(n_53), .A(n_15), .B(in_39[0]), .CI(n_25));
  ADDFX1 g9399(.CO(n_50), .S(n_51), .A(in_78), .B(n_31), .CI(n_3));
  ADDFX1 g9400(.CO(n_48), .S(n_49), .A(n_19), .B(in_15[1]), .CI(n_30));
  ADDFX1 g9401(.CO(n_46), .S(n_47), .A(in_14[0]), .B(n_24), .CI(n_18));
  ADDFX1 g9402(.CO(n_44), .S(n_45), .A(n_8), .B(n_4), .CI(in_69[1]));
  OAI2BB1X1 g9403(.Y(n_43), .A0N(n_22), .A1N(n_38), .B0(n_40));
  ADDHX1 g9404(.CO(n_41), .S(n_42), .A(in_24[1]), .B(in_84[1]));
  OR2X1 g9405(.Y(n_40), .A(n_22), .B(n_38));
  XNOR2X1 g9406(.Y(n_39), .A(in_90[0]), .B(in_60[0]));
  XNOR2X1 g9407(.Y(n_38), .A(in_45[0]), .B(in_7[2]));
  INVX1 g9409(.Y(n_37), .A(in_77[0]));
  INVX1 g9410(.Y(n_36), .A(in_35[1]));
  INVX1 g9411(.Y(n_35), .A(in_13[2]));
  INVX1 g9412(.Y(n_34), .A(in_16[2]));
  INVX1 g9413(.Y(n_33), .A(in_53[1]));
  INVX1 g9414(.Y(n_32), .A(in_42[0]));
  INVX1 g9415(.Y(n_31), .A(in_41[0]));
  INVX1 g9416(.Y(n_30), .A(in_23[1]));
  INVX1 g9417(.Y(n_29), .A(in_61[0]));
  INVX1 g9418(.Y(n_28), .A(in_1[1]));
  INVX1 g9419(.Y(n_27), .A(in_4[0]));
  INVX1 g9420(.Y(n_26), .A(in_65[1]));
  INVX1 g9421(.Y(n_25), .A(in_10[0]));
  INVX1 g9422(.Y(n_24), .A(in_26[0]));
  INVX1 g9423(.Y(n_23), .A(in_62[0]));
  INVX1 g9424(.Y(n_22), .A(in_14[3]));
  INVX1 g9425(.Y(n_21), .A(in_85[1]));
  INVX1 g9426(.Y(n_20), .A(in_47[1]));
  INVX1 g9427(.Y(n_19), .A(in_82[1]));
  INVX1 g9428(.Y(n_18), .A(in_73[0]));
  INVX1 g9429(.Y(n_17), .A(in_83[0]));
  INVX1 g9430(.Y(n_16), .A(in_68[1]));
  INVX1 g9431(.Y(n_15), .A(in_2[0]));
  INVX1 g9432(.Y(n_14), .A(in_5[1]));
  INVX1 g9433(.Y(n_13), .A(in_8[0]));
  INVX1 g9434(.Y(n_12), .A(in_54[1]));
  INVX1 g9435(.Y(n_11), .A(in_31[0]));
  INVX1 g9436(.Y(n_10), .A(in_25[0]));
  INVX1 g9437(.Y(n_9), .A(in_43[1]));
  INVX1 g9438(.Y(n_8), .A(in_32[1]));
  INVX1 g9439(.Y(n_7), .A(in_66[0]));
  INVX1 g9440(.Y(n_6), .A(in_11[1]));
  INVX1 g9441(.Y(n_5), .A(in_30[1]));
  INVX1 g9442(.Y(n_4), .A(in_38[1]));
  INVX1 g9443(.Y(n_3), .A(in_19[0]));
  INVX1 g9444(.Y(n_2), .A(in_20[0]));
  NOR2BX1 g2(.Y(n_0), .AN(in_60[0]), .B(in_90[0]));
endmodule

module WALLACE_CSA_DUMMY_OP102_group_106219(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, in_85, in_86, in_87, out_0);
input  in_38, in_45, in_46, in_51, in_58, in_59, in_60, in_67, in_73, in_74, 
    in_75;
input   [4:0] in_0;
input   [9:0] in_1;
input   [9:0] in_2;
input   [6:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [1:0] in_34;
input   [1:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [1:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
input   [1:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [1:0] in_50;
input   [4:0] in_52;
input   [4:0] in_53;
input   [1:0] in_54;
input   [2:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [1:0] in_61;
input   [4:0] in_62;
input   [1:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [1:0] in_68;
input   [1:0] in_69;
input   [4:0] in_70;
input   [4:0] in_71;
input   [1:0] in_72;
input   [4:0] in_76;
input   [1:0] in_77;
input   [4:0] in_78;
input   [4:0] in_79;
input   [1:0] in_80;
input   [4:0] in_81;
input   [4:0] in_82;
input   [3:0] in_83;
input   [4:0] in_84;
input   [4:0] in_85;
input   [1:0] in_86;
input   [4:0] in_87;
output  [9:0] out_0;
wire  n_262, n_260, n_258, n_256, n_254, n_253, n_252, n_250, n_249, n_248, 
    n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_238, n_237, 
    n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, n_227, 
    n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, n_218, n_217, 
    n_216, n_215, n_214, n_213, n_212, n_210, n_209, n_208, n_207, n_206, 
    n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, 
    n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, n_187, n_186, 
    n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, 
    n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, 
    n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156, 
    n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, 
    n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, 
    n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, 
    n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, 
    n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, 
    n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, 
    n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, 
    n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, 
    n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, 
    n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, 
    n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, 
    n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, 
    n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_75, in_74, 
    in_73, in_67, in_60, in_59, in_58, in_51, in_46, in_45, in_38;
wire   [9:0] out_0;
wire   [3:0] in_83;
wire   [2:0] in_55;
wire   [1:0] in_86;
wire   [1:0] in_80;
wire   [1:0] in_77;
wire   [1:0] in_72;
wire   [1:0] in_69;
wire   [1:0] in_68;
wire   [1:0] in_63;
wire   [1:0] in_61;
wire   [1:0] in_54;
wire   [1:0] in_50;
wire   [1:0] in_42;
wire   [1:0] in_41;
wire   [1:0] in_39;
wire   [1:0] in_37;
wire   [1:0] in_35;
wire   [1:0] in_34;
wire   [1:0] in_31;
wire   [1:0] in_29;
wire   [1:0] in_27;
wire   [1:0] in_25;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [6:0] in_3;
wire   [9:0] in_2;
wire   [9:0] in_1;
wire   [4:0] in_87;
wire   [4:0] in_85;
wire   [4:0] in_84;
wire   [4:0] in_82;
wire   [4:0] in_81;
wire   [4:0] in_79;
wire   [4:0] in_78;
wire   [4:0] in_76;
wire   [4:0] in_71;
wire   [4:0] in_70;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_62;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_40;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g8637(.Y(out_0[9]), .A(n_262));
  ADDFX1 g8638(.CO(n_262), .S(out_0[7]), .A(n_190), .B(n_244), .CI(n_260));
  ADDFX1 g8639(.CO(n_260), .S(out_0[6]), .A(n_245), .B(n_252), .CI(n_258));
  ADDFX1 g8640(.CO(n_258), .S(out_0[5]), .A(n_253), .B(n_248), .CI(n_256));
  ADDFX1 g8641(.CO(n_256), .S(out_0[4]), .A(n_246), .B(n_249), .CI(n_254));
  ADDFX1 g8642(.CO(n_254), .S(out_0[3]), .A(n_236), .B(n_250), .CI(n_247));
  ADDFX1 g8643(.CO(n_252), .S(n_253), .A(n_230), .B(n_241), .CI(n_242));
  ADDFX1 g8644(.CO(n_250), .S(out_0[2]), .A(n_229), .B(n_238), .CI(n_237));
  ADDFX1 g8645(.CO(n_248), .S(n_249), .A(n_232), .B(n_234), .CI(n_243));
  ADDFX1 g8646(.CO(n_246), .S(n_247), .A(n_228), .B(n_233), .CI(n_235));
  ADDFX1 g8647(.CO(n_244), .S(n_245), .A(n_184), .B(n_191), .CI(n_240));
  ADDFX1 g8648(.CO(n_242), .S(n_243), .A(n_218), .B(n_220), .CI(n_231));
  ADDFX1 g8649(.CO(n_240), .S(n_241), .A(n_224), .B(n_196), .CI(n_185));
  ADDFX1 g8650(.CO(n_238), .S(out_0[1]), .A(n_210), .B(n_223), .CI(n_199));
  ADDFX1 g8651(.CO(n_236), .S(n_237), .A(n_222), .B(n_227), .CI(n_217));
  ADDFX1 g8652(.CO(n_234), .S(n_235), .A(n_216), .B(n_221), .CI(n_219));
  ADDFX1 g8653(.CO(n_232), .S(n_233), .A(n_214), .B(n_226), .CI(n_193));
  ADDFX1 g8654(.CO(n_230), .S(n_231), .A(n_192), .B(n_225), .CI(n_197));
  ADDFX1 g8655(.CO(n_228), .S(n_229), .A(n_203), .B(n_215), .CI(n_198));
  ADDFX1 g8656(.CO(n_226), .S(n_227), .A(n_194), .B(n_212), .CI(n_209));
  ADDFX1 g8657(.CO(n_224), .S(n_225), .A(n_0), .B(n_206), .CI(n_200));
  ADDFX1 g8658(.CO(n_222), .S(n_223), .A(n_195), .B(n_186), .CI(n_213));
  ADDFX1 g8659(.CO(n_220), .S(n_221), .A(n_202), .B(n_201), .CI(n_204));
  ADDFX1 g8660(.CO(n_218), .S(n_219), .A(n_162), .B(n_207), .CI(n_208));
  ADDFX1 g8661(.CO(n_216), .S(n_217), .A(n_163), .B(n_156), .CI(n_205));
  ADDFX1 g8662(.CO(n_214), .S(n_215), .A(n_171), .B(n_176), .CI(n_164));
  ADDFX1 g8663(.CO(n_212), .S(n_213), .A(n_174), .B(n_177), .CI(n_154));
  ADDFX1 g8664(.CO(n_210), .S(out_0[0]), .A(n_175), .B(n_187), .CI(n_155));
  ADDFX1 g8665(.CO(n_208), .S(n_209), .A(n_179), .B(n_168), .CI(in_1[2]));
  ADDFX1 g8666(.CO(n_206), .S(n_207), .A(n_137), .B(n_178), .CI(n_172));
  ADDFX1 g8667(.CO(n_204), .S(n_205), .A(n_182), .B(n_173), .CI(in_2[2]));
  ADDFX1 g8668(.CO(n_202), .S(n_203), .A(n_160), .B(n_166), .CI(n_159));
  ADDFX1 g8669(.CO(n_200), .S(n_201), .A(n_131), .B(n_181), .CI(in_2[3]));
  ADDFX1 g8670(.CO(n_198), .S(n_199), .A(n_167), .B(n_157), .CI(n_165));
  ADDFX1 g8671(.CO(n_196), .S(n_197), .A(n_180), .B(in_2[4]), .CI(in_1[4]));
  ADDFX1 g8672(.CO(n_194), .S(n_195), .A(n_161), .B(n_183), .CI(n_169));
  ADDFX1 g8673(.CO(n_192), .S(n_193), .A(n_158), .B(n_170), .CI(in_1[3]));
  INVX1 g8674(.Y(n_191), .A(n_189));
  INVX1 g8675(.Y(n_190), .A(n_188));
  ADDFX1 g8676(.CO(n_188), .S(n_189), .A(n_147), .B(in_2[6]), .CI(in_1[6]));
  ADDFX1 g8677(.CO(n_186), .S(n_187), .A(n_122), .B(n_149), .CI(n_120));
  ADDFX1 g8678(.CO(n_184), .S(n_185), .A(n_147), .B(in_2[5]), .CI(in_1[5]));
  ADDFX1 g8679(.CO(n_182), .S(n_183), .A(n_153), .B(n_124), .CI(n_148));
  ADDFX1 g8680(.CO(n_180), .S(n_181), .A(n_142), .B(n_129), .CI(n_117));
  ADDFX1 g8681(.CO(n_178), .S(n_179), .A(n_123), .B(n_109), .CI(n_152));
  ADDFX1 g8682(.CO(n_176), .S(n_177), .A(n_150), .B(n_135), .CI(n_128));
  ADDFX1 g8683(.CO(n_174), .S(n_175), .A(n_141), .B(n_136), .CI(n_151));
  ADDFX1 g8684(.CO(n_172), .S(n_173), .A(n_133), .B(n_113), .CI(n_104));
  ADDFX1 g8685(.CO(n_170), .S(n_171), .A(n_115), .B(n_127), .CI(n_111));
  ADDFX1 g8686(.CO(n_168), .S(n_169), .A(n_106), .B(n_134), .CI(n_140));
  ADDFX1 g8687(.CO(n_166), .S(n_167), .A(n_114), .B(n_110), .CI(n_138));
  ADDFX1 g8688(.CO(n_164), .S(n_165), .A(n_145), .B(n_119), .CI(in_2[1]));
  ADDFX1 g8689(.CO(n_162), .S(n_163), .A(n_118), .B(n_144), .CI(n_132));
  ADDFX1 g8690(.CO(n_160), .S(n_161), .A(n_107), .B(n_126), .CI(n_121));
  ADDFX1 g8691(.CO(n_158), .S(n_159), .A(n_125), .B(n_130), .CI(n_143));
  ADDFX1 g8692(.CO(n_156), .S(n_157), .A(n_112), .B(n_116), .CI(in_1[1]));
  ADDFX1 g8693(.CO(n_154), .S(n_155), .A(n_108), .B(n_139), .CI(in_1[0]));
  ADDFX1 g8695(.CO(n_152), .S(n_153), .A(n_89), .B(n_63), .CI(n_99));
  ADDFX1 g8696(.CO(n_150), .S(n_151), .A(n_92), .B(n_46), .CI(n_64));
  ADDFX1 g8697(.CO(n_148), .S(n_149), .A(n_98), .B(n_40), .CI(n_90));
  NOR2X1 g8699(.Y(n_147), .A(n_28), .B(n_146));
  ADDFX1 g8700(.CO(n_144), .S(n_145), .A(n_37), .B(n_60), .CI(n_31));
  ADDFX1 g8701(.CO(n_142), .S(n_143), .A(n_83), .B(n_55), .CI(n_87));
  ADDFX1 g8702(.CO(n_140), .S(n_141), .A(n_76), .B(n_52), .CI(n_96));
  ADDFX1 g8703(.CO(n_138), .S(n_139), .A(n_70), .B(n_50), .CI(n_94));
  ADDFX1 g8704(.CO(n_146), .S(n_137), .A(n_30), .B(n_57), .CI(n_103));
  ADDFX1 g8705(.CO(n_135), .S(n_136), .A(n_74), .B(n_36), .CI(n_100));
  ADDFX1 g8706(.CO(n_133), .S(n_134), .A(n_97), .B(n_93), .CI(n_91));
  ADDFX1 g8707(.CO(n_131), .S(n_132), .A(n_53), .B(n_105), .CI(n_67));
  ADDFX1 g8708(.CO(n_129), .S(n_130), .A(n_77), .B(n_43), .CI(n_85));
  ADDFX1 g8709(.CO(n_127), .S(n_128), .A(n_78), .B(n_84), .CI(n_88));
  ADDFX1 g8710(.CO(n_125), .S(n_126), .A(n_95), .B(n_71), .CI(n_81));
  ADDFX1 g8711(.CO(n_123), .S(n_124), .A(n_49), .B(n_47), .CI(n_73));
  ADDFX1 g8712(.CO(n_121), .S(n_122), .A(n_82), .B(n_48), .CI(n_42));
  ADDFX1 g8713(.CO(n_119), .S(n_120), .A(n_38), .B(n_32), .CI(in_2[0]));
  ADDFX1 g8714(.CO(n_117), .S(n_118), .A(n_79), .B(n_58), .CI(n_59));
  ADDFX1 g8715(.CO(n_115), .S(n_116), .A(n_86), .B(n_44), .CI(n_56));
  ADDFX1 g8716(.CO(n_113), .S(n_114), .A(n_75), .B(n_41), .CI(n_51));
  ADDFX1 g8717(.CO(n_111), .S(n_112), .A(n_80), .B(n_54), .CI(n_68));
  ADDFX1 g8718(.CO(n_109), .S(n_110), .A(n_39), .B(n_35), .CI(n_69));
  ADDFX1 g8719(.CO(n_107), .S(n_108), .A(in_18[0]), .B(in_23[0]), .CI(n_72));
  ADDFX1 g8720(.CO(n_105), .S(n_106), .A(in_79[1]), .B(n_18), .CI(n_45));
  INVX1 g8721(.Y(n_104), .A(n_102));
  INVX1 g8722(.Y(n_103), .A(n_101));
  ADDFX1 g8723(.CO(n_101), .S(n_102), .A(in_79[1]), .B(in_3[2]), .CI(n_29));
  ADDFX1 g8724(.CO(n_99), .S(n_100), .A(in_35[0]), .B(in_54[0]), .CI(in_61[0]));
  ADDFX1 g8725(.CO(n_97), .S(n_98), .A(in_60), .B(in_74), .CI(n_5));
  ADDFX1 g8726(.CO(n_95), .S(n_96), .A(in_37[0]), .B(in_69[0]), .CI(in_72[0]));
  ADDFX1 g8727(.CO(n_93), .S(n_94), .A(in_67), .B(in_11[0]), .CI(in_68[0]));
  ADDFX1 g8728(.CO(n_91), .S(n_92), .A(in_46), .B(n_8), .CI(in_55[0]));
  ADDFX1 g8729(.CO(n_89), .S(n_90), .A(in_25[0]), .B(n_3), .CI(n_11));
  ADDFX1 g8730(.CO(n_87), .S(n_88), .A(in_50[0]), .B(in_72[0]), .CI(in_14[1]));
  ADDFX1 g8731(.CO(n_85), .S(n_86), .A(in_61[0]), .B(n_27), .CI(n_17));
  INVX1 g8732(.Y(n_84), .A(n_66));
  INVX1 g8733(.Y(n_83), .A(n_65));
  INVX1 g8734(.Y(n_82), .A(n_62));
  INVX1 g8735(.Y(n_81), .A(n_61));
  INVX1 g8736(.Y(n_80), .A(n_34));
  INVX1 g8737(.Y(n_79), .A(n_33));
  ADDFX1 g8738(.CO(n_77), .S(n_78), .A(in_15[1]), .B(n_15), .CI(n_25));
  ADDFX1 g8739(.CO(n_75), .S(n_76), .A(in_10[0]), .B(in_20[0]), .CI(n_13));
  ADDFX1 g8740(.CO(n_73), .S(n_74), .A(in_34[0]), .B(n_10), .CI(in_75));
  ADDFX1 g8741(.CO(n_71), .S(n_72), .A(in_40[0]), .B(n_20), .CI(n_26));
  ADDFX1 g8742(.CO(n_69), .S(n_70), .A(in_5[0]), .B(in_31[0]), .CI(in_45));
  ADDFX1 g8743(.CO(n_67), .S(n_68), .A(in_18[1]), .B(in_21[1]), .CI(in_3[1]));
  ADDFX1 g8744(.CO(n_65), .S(n_66), .A(in_47[1]), .B(in_13[1]), .CI(in_48[1]));
  ADDFX1 g8745(.CO(n_63), .S(n_64), .A(in_27[0]), .B(n_16), .CI(in_58));
  ADDFX1 g8746(.CO(n_61), .S(n_62), .A(in_16[0]), .B(in_52[0]), .CI(in_65[0]));
  ADDFX1 g8747(.CO(n_59), .S(n_60), .A(in_9[1]), .B(in_22[1]), .CI(in_12[1]));
  ADDFX1 g8748(.CO(n_57), .S(n_58), .A(n_1), .B(in_83[2]), .CI(n_14));
  ADDFX1 g8749(.CO(n_55), .S(n_56), .A(in_42[1]), .B(n_9), .CI(in_68[0]));
  ADDFX1 g8750(.CO(n_53), .S(n_54), .A(in_19[1]), .B(n_24), .CI(n_22));
  ADDFX1 g8751(.CO(n_51), .S(n_52), .A(in_29[0]), .B(in_50[0]), .CI(in_77[0]));
  ADDFX1 g8752(.CO(n_49), .S(n_50), .A(n_21), .B(in_59), .CI(n_4));
  ADDFX1 g8753(.CO(n_47), .S(n_48), .A(in_3[0]), .B(in_62[0]), .CI(n_23));
  ADDFX1 g8754(.CO(n_45), .S(n_46), .A(n_6), .B(n_7), .CI(in_63[0]));
  ADDFX1 g8755(.CO(n_43), .S(n_44), .A(in_39[1]), .B(in_41[1]), .CI(in_55[0]));
  ADDFX1 g8756(.CO(n_41), .S(n_42), .A(in_38), .B(in_80[0]), .CI(n_12));
  ADDFX1 g8757(.CO(n_39), .S(n_40), .A(in_51), .B(n_2), .CI(in_86[0]));
  ADDFX1 g8758(.CO(n_37), .S(n_38), .A(in_17[0]), .B(in_21[0]), .CI(in_6[0]));
  ADDFX1 g8759(.CO(n_35), .S(n_36), .A(in_4[0]), .B(n_19), .CI(in_73));
  ADDFX1 g8760(.CO(n_33), .S(n_34), .A(in_36[1]), .B(in_49[1]), .CI(in_76[1]));
  ADDFX1 g8761(.CO(n_31), .S(n_32), .A(in_22[0]), .B(in_9[0]), .CI(in_12[0]));
  INVX1 g8762(.Y(n_30), .A(n_28));
  XNOR2X1 g8763(.Y(n_29), .A(in_70[2]), .B(in_62[0]));
  NOR2X1 g8764(.Y(n_28), .A(in_70[2]), .B(in_62[0]));
  INVX1 g8765(.Y(n_27), .A(in_84[1]));
  INVX1 g8766(.Y(n_26), .A(in_81[0]));
  INVX1 g8767(.Y(n_25), .A(in_64[1]));
  INVX1 g8768(.Y(n_24), .A(in_78[1]));
  INVX1 g8769(.Y(n_23), .A(in_66[0]));
  INVX1 g8770(.Y(n_22), .A(in_23[1]));
  INVX1 g8771(.Y(n_21), .A(in_8[0]));
  INVX1 g8772(.Y(n_20), .A(in_26[0]));
  INVX1 g8773(.Y(n_19), .A(in_56[0]));
  INVX1 g8774(.Y(n_18), .A(in_6[1]));
  INVX1 g8775(.Y(n_17), .A(in_53[1]));
  INVX1 g8776(.Y(n_16), .A(in_28[0]));
  INVX1 g8777(.Y(n_15), .A(in_43[1]));
  INVX1 g8778(.Y(n_14), .A(in_11[0]));
  INVX1 g8779(.Y(n_13), .A(in_44[0]));
  INVX1 g8780(.Y(n_12), .A(in_85[0]));
  INVX1 g8781(.Y(n_11), .A(in_87[0]));
  INVX1 g8782(.Y(n_10), .A(in_24[0]));
  INVX1 g8783(.Y(n_9), .A(in_57[1]));
  INVX1 g8784(.Y(n_8), .A(in_30[0]));
  INVX1 g8785(.Y(n_7), .A(in_33[0]));
  INVX1 g8786(.Y(n_6), .A(in_32[0]));
  INVX1 g8787(.Y(n_5), .A(in_71[0]));
  INVX1 g8788(.Y(n_4), .A(in_7[0]));
  INVX1 g8789(.Y(n_3), .A(in_0[0]));
  INVX1 g8790(.Y(n_2), .A(in_82[0]));
  INVX1 g8791(.Y(n_1), .A(in_40[0]));
  AO21X1 g2(.Y(n_0), .A0(n_28), .A1(n_146), .B0(n_147));
endmodule

module WALLACE_CSA_DUMMY_OP106_group_109836_6302(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, out_0);
input  in_23, in_24, in_35, in_36, in_37;
input   [4:0] in_0;
input   [2:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [4:0] in_4;
input   [4:0] in_5;
input   [9:0] in_6;
input   [6:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [2:0] in_20;
input   [2:0] in_21;
input   [4:0] in_22;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [1:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [1:0] in_44;
input   [4:0] in_45;
output  [9:0] out_0;
wire  n_144, n_142, n_140, n_138, n_136, n_135, n_134, n_133, n_132, n_130, 
    n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, 
    n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_37, 
    in_36, in_35, in_24, in_23;
wire   [9:0] out_0;
wire   [1:0] in_44;
wire   [1:0] in_41;
wire   [1:0] in_38;
wire   [1:0] in_32;
wire   [1:0] in_31;
wire   [1:0] in_27;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_7;
wire   [9:0] in_6;
wire   [2:0] in_21;
wire   [2:0] in_20;
wire   [2:0] in_1;
wire   [4:0] in_45;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_22;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_5;
wire   [4:0] in_4;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  INVX1 g1701(.Y(out_0[9]), .A(n_144));
  ADDFX1 g1702(.CO(n_144), .S(out_0[6]), .A(n_20), .B(n_124), .CI(n_142));
  ADDFX1 g1703(.CO(n_142), .S(out_0[5]), .A(n_125), .B(n_132), .CI(n_140));
  ADDFX1 g1704(.CO(n_140), .S(out_0[4]), .A(n_134), .B(n_133), .CI(n_138));
  ADDFX1 g1705(.CO(n_138), .S(out_0[3]), .A(n_128), .B(n_135), .CI(n_136));
  ADDFX1 g1706(.CO(n_136), .S(out_0[2]), .A(n_123), .B(n_130), .CI(n_129));
  ADDFX1 g1707(.CO(n_134), .S(n_135), .A(n_122), .B(n_115), .CI(n_127));
  ADDFX1 g1708(.CO(n_132), .S(n_133), .A(n_114), .B(n_126), .CI(n_117));
  ADDFX1 g1709(.CO(n_130), .S(out_0[1]), .A(n_121), .B(n_110), .CI(n_109));
  ADDFX1 g1710(.CO(n_128), .S(n_129), .A(n_120), .B(n_108), .CI(n_119));
  ADDFX1 g1711(.CO(n_126), .S(n_127), .A(n_99), .B(n_112), .CI(n_118));
  ADDFX1 g1712(.CO(n_124), .S(n_125), .A(n_100), .B(in_6[5]), .CI(n_116));
  ADDFX1 g1713(.CO(n_122), .S(n_123), .A(n_97), .B(n_106), .CI(n_113));
  ADDFX1 g1714(.CO(n_120), .S(n_121), .A(n_95), .B(n_105), .CI(n_107));
  ADDFX1 g1715(.CO(n_118), .S(n_119), .A(n_104), .B(n_94), .CI(in_6[2]));
  ADDFX1 g1716(.CO(n_116), .S(n_117), .A(n_101), .B(n_98), .CI(in_6[4]));
  ADDFX1 g1717(.CO(n_114), .S(n_115), .A(n_102), .B(n_96), .CI(in_6[3]));
  ADDFX1 g1718(.CO(n_112), .S(n_113), .A(n_78), .B(n_81), .CI(n_103));
  ADDFX1 g1719(.CO(n_110), .S(out_0[0]), .A(n_85), .B(n_83), .CI(n_93));
  ADDFX1 g1720(.CO(n_108), .S(n_109), .A(n_82), .B(n_92), .CI(in_6[1]));
  ADDFX1 g1721(.CO(n_106), .S(n_107), .A(n_87), .B(n_73), .CI(n_79));
  ADDFX1 g1722(.CO(n_104), .S(n_105), .A(n_66), .B(n_84), .CI(n_89));
  ADDFX1 g1723(.CO(n_102), .S(n_103), .A(n_88), .B(n_86), .CI(n_68));
  ADDHX1 g1724(.CO(n_100), .S(n_101), .A(n_48), .B(n_90));
  ADDFX1 g1725(.CO(n_98), .S(n_99), .A(n_74), .B(n_80), .CI(n_91));
  ADDFX1 g1726(.CO(n_96), .S(n_97), .A(n_71), .B(n_72), .CI(n_75));
  ADDFX1 g1727(.CO(n_94), .S(n_95), .A(n_60), .B(n_76), .CI(n_69));
  ADDFX1 g1728(.CO(n_92), .S(n_93), .A(n_67), .B(n_77), .CI(in_6[0]));
  ADDFX1 g1729(.CO(n_90), .S(n_91), .A(n_44), .B(n_63), .CI(n_70));
  ADDFX1 g1730(.CO(n_88), .S(n_89), .A(n_49), .B(n_61), .CI(n_53));
  ADDFX1 g1731(.CO(n_86), .S(n_87), .A(n_31), .B(n_51), .CI(n_57));
  ADDFX1 g1732(.CO(n_84), .S(n_85), .A(n_34), .B(n_58), .CI(n_28));
  ADDFX1 g1733(.CO(n_82), .S(n_83), .A(n_32), .B(n_54), .CI(n_65));
  ADDFX1 g1734(.CO(n_80), .S(n_81), .A(n_24), .B(n_45), .CI(n_59));
  ADDFX1 g1735(.CO(n_78), .S(n_79), .A(n_47), .B(n_30), .CI(n_64));
  ADDFX1 g1736(.CO(n_76), .S(n_77), .A(n_62), .B(n_56), .CI(n_52));
  ADDFX1 g1737(.CO(n_74), .S(n_75), .A(n_25), .B(n_39), .CI(n_29));
  ADDFX1 g1738(.CO(n_72), .S(n_73), .A(n_41), .B(n_26), .CI(n_36));
  ADDFX1 g1739(.CO(n_70), .S(n_71), .A(n_46), .B(n_35), .CI(n_40));
  ADDFX1 g1740(.CO(n_68), .S(n_69), .A(n_55), .B(n_33), .CI(n_27));
  ADDFX1 g1741(.CO(n_66), .S(n_67), .A(in_12[0]), .B(in_9[0]), .CI(n_50));
  ADDFX1 g1742(.CO(n_64), .S(n_65), .A(in_41[0]), .B(n_23), .CI(in_11[0]));
  XNOR2X1 g1743(.Y(n_63), .A(n_21), .B(n_38));
  ADDFX1 g1744(.CO(n_61), .S(n_62), .A(in_18[0]), .B(in_44[0]), .CI(in_28[0]));
  ADDFX1 g1745(.CO(n_59), .S(n_60), .A(n_22), .B(n_7), .CI(in_16[1]));
  ADDFX1 g1746(.CO(n_57), .S(n_58), .A(in_31[0]), .B(n_11), .CI(in_37));
  ADDFX1 g1747(.CO(n_55), .S(n_56), .A(n_3), .B(in_35), .CI(in_10[0]));
  ADDFX1 g1748(.CO(n_53), .S(n_54), .A(in_23), .B(in_24), .CI(n_4));
  ADDFX1 g1749(.CO(n_51), .S(n_52), .A(in_21[0]), .B(n_2), .CI(n_19));
  ADDFX1 g1750(.CO(n_49), .S(n_50), .A(n_14), .B(n_1), .CI(in_25[0]));
  NOR2BX1 g1751(.Y(n_48), .AN(n_21), .B(n_38));
  ADDFX1 g1752(.CO(n_46), .S(n_47), .A(in_7[1]), .B(in_1[1]), .CI(n_16));
  INVX1 g1753(.Y(n_45), .A(n_43));
  INVX1 g1754(.Y(n_44), .A(n_42));
  ADDFX1 g1755(.CO(n_42), .S(n_43), .A(in_43[0]), .B(in_16[2]), .CI(in_12[2]));
  ADDFX1 g1756(.CO(n_40), .S(n_41), .A(in_20[1]), .B(n_5), .CI(in_38[1]));
  INVX1 g1757(.Y(n_39), .A(n_37));
  ADDFX1 g1758(.CO(n_38), .S(n_37), .A(in_18[0]), .B(in_10[0]), .CI(in_25[0]));
  ADDFX1 g1759(.CO(n_35), .S(n_36), .A(in_14[1]), .B(n_18), .CI(n_13));
  ADDFX1 g1760(.CO(n_33), .S(n_34), .A(in_7[0]), .B(in_27[0]), .CI(in_36));
  ADDFX1 g1761(.CO(n_31), .S(n_32), .A(n_12), .B(n_8), .CI(in_43[0]));
  ADDFX1 g1762(.CO(n_29), .S(n_30), .A(n_17), .B(in_9[1]), .CI(in_12[1]));
  ADDFX1 g1763(.CO(n_27), .S(n_28), .A(in_30[0]), .B(n_6), .CI(n_15));
  ADDFX1 g1764(.CO(n_25), .S(n_26), .A(n_10), .B(n_9), .CI(in_21[0]));
  OAI21X1 g1765(.Y(n_24), .A0(in_28[0]), .A1(in_30[0]), .B0(n_21));
  XNOR2X1 g1766(.Y(n_23), .A(in_0[0]), .B(in_32[0]));
  NOR2BX1 g1767(.Y(n_22), .AN(in_32[0]), .B(in_0[0]));
  NAND2X1 g1768(.Y(n_21), .A(in_30[0]), .B(in_28[0]));
  INVX1 g1769(.Y(n_20), .A(in_6[6]));
  INVX1 g1770(.Y(n_19), .A(in_39[0]));
  INVX1 g1771(.Y(n_18), .A(in_40[1]));
  INVX1 g1772(.Y(n_17), .A(in_33[1]));
  INVX1 g1773(.Y(n_16), .A(in_26[1]));
  INVX1 g1774(.Y(n_15), .A(in_45[0]));
  INVX1 g1775(.Y(n_14), .A(in_4[0]));
  INVX1 g1776(.Y(n_13), .A(in_34[1]));
  INVX1 g1777(.Y(n_12), .A(in_3[0]));
  INVX1 g1778(.Y(n_11), .A(in_22[0]));
  INVX1 g1779(.Y(n_10), .A(in_15[1]));
  INVX1 g1780(.Y(n_9), .A(in_19[1]));
  INVX1 g1781(.Y(n_8), .A(in_42[0]));
  INVX1 g1782(.Y(n_7), .A(in_11[1]));
  INVX1 g1783(.Y(n_6), .A(in_8[0]));
  INVX1 g1784(.Y(n_5), .A(in_2[1]));
  INVX1 g1785(.Y(n_4), .A(in_5[0]));
  INVX1 g1786(.Y(n_3), .A(in_13[0]));
  INVX1 g1787(.Y(n_2), .A(in_29[0]));
  INVX1 g1788(.Y(n_1), .A(in_17[0]));
endmodule

module WALLACE_CSA_DUMMY_OP106_group_109836(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, out_0);
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [4:0] in_5;
input   [6:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [4:0] in_12;
input   [1:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [2:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [1:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
output  [9:0] out_0;
wire  n_127, n_125, n_123, n_121, n_120, n_119, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_105, n_104, n_103, 
    n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_0;
wire   [9:0] out_0;
wire   [1:0] in_30;
wire   [1:0] in_29;
wire   [1:0] in_22;
wire   [1:0] in_13;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [6:0] in_6;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_12;
wire   [4:0] in_5;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_24;
wire   [2:0] in_3;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3867(.Y(out_0[9]), .A(n_127));
  ADDFX1 g3868(.CO(n_127), .S(out_0[5]), .A(n_91), .B(n_113), .CI(n_125));
  ADDFX1 g3869(.CO(n_125), .S(out_0[4]), .A(n_114), .B(n_119), .CI(n_123));
  ADDFX1 g3870(.CO(n_123), .S(out_0[3]), .A(n_115), .B(n_120), .CI(n_121));
  ADDFX1 g3871(.CO(n_121), .S(out_0[2]), .A(n_109), .B(n_116), .CI(n_117));
  ADDFX1 g3872(.CO(n_119), .S(n_120), .A(n_103), .B(n_108), .CI(n_111));
  ADDFX1 g3873(.CO(n_117), .S(out_0[1]), .A(n_102), .B(n_105), .CI(n_110));
  ADDFX1 g3874(.CO(n_115), .S(n_116), .A(n_101), .B(n_104), .CI(n_112));
  ADDFX1 g3875(.CO(n_113), .S(n_114), .A(n_92), .B(n_95), .CI(n_107));
  ADDFX1 g3876(.CO(n_111), .S(n_112), .A(n_93), .B(n_99), .CI(n_98));
  ADDFX1 g3877(.CO(n_109), .S(n_110), .A(n_87), .B(n_94), .CI(n_100));
  ADDFX1 g3878(.CO(n_107), .S(n_108), .A(n_89), .B(n_97), .CI(n_96));
  ADDFX1 g3879(.CO(n_105), .S(out_0[0]), .A(n_68), .B(n_76), .CI(n_88));
  ADDFX1 g3880(.CO(n_103), .S(n_104), .A(n_69), .B(n_82), .CI(n_90));
  ADDFX1 g3881(.CO(n_101), .S(n_102), .A(n_75), .B(n_84), .CI(n_70));
  ADDFX1 g3882(.CO(n_99), .S(n_100), .A(n_80), .B(n_67), .CI(n_77));
  ADDFX1 g3883(.CO(n_97), .S(n_98), .A(n_71), .B(n_66), .CI(n_83));
  ADDFX1 g3884(.CO(n_95), .S(n_96), .A(n_63), .B(n_81), .CI(n_86));
  ADDFX1 g3885(.CO(n_93), .S(n_94), .A(n_62), .B(n_74), .CI(n_72));
  ADDHX1 g3886(.CO(n_91), .S(n_92), .A(n_16), .B(n_85));
  ADDFX1 g3887(.CO(n_89), .S(n_90), .A(n_64), .B(n_79), .CI(n_73));
  ADDFX1 g3888(.CO(n_87), .S(n_88), .A(n_28), .B(n_40), .CI(n_78));
  ADDFX1 g3889(.CO(n_85), .S(n_86), .A(n_0), .B(n_22), .CI(n_65));
  ADDFX1 g3890(.CO(n_83), .S(n_84), .A(n_26), .B(n_50), .CI(n_54));
  ADDFX1 g3891(.CO(n_81), .S(n_82), .A(n_23), .B(n_43), .CI(n_61));
  ADDFX1 g3892(.CO(n_79), .S(n_80), .A(n_59), .B(n_29), .CI(n_31));
  ADDFX1 g3893(.CO(n_77), .S(n_78), .A(n_30), .B(n_48), .CI(n_60));
  ADDFX1 g3894(.CO(n_75), .S(n_76), .A(n_46), .B(n_58), .CI(n_32));
  ADDFX1 g3895(.CO(n_73), .S(n_74), .A(n_27), .B(n_21), .CI(n_57));
  ADDFX1 g3896(.CO(n_71), .S(n_72), .A(n_45), .B(n_37), .CI(n_47));
  ADDFX1 g3897(.CO(n_69), .S(n_70), .A(n_34), .B(n_39), .CI(n_44));
  ADDFX1 g3898(.CO(n_67), .S(n_68), .A(in_16[0]), .B(n_38), .CI(n_24));
  ADDFX1 g3899(.CO(n_65), .S(n_66), .A(n_49), .B(n_33), .CI(n_25));
  ADDFX1 g3900(.CO(n_63), .S(n_64), .A(in_38[0]), .B(n_15), .CI(n_53));
  ADDFX1 g3901(.CO(n_61), .S(n_62), .A(n_3), .B(n_19), .CI(in_10[1]));
  ADDFX1 g3902(.CO(n_59), .S(n_60), .A(in_11[0]), .B(n_10), .CI(in_30[0]));
  INVX1 g3903(.Y(n_58), .A(n_56));
  INVX1 g3904(.Y(n_57), .A(n_55));
  ADDFX1 g3905(.CO(n_55), .S(n_56), .A(in_1[0]), .B(in_2[0]), .CI(in_14[0]));
  INVX1 g3906(.Y(n_54), .A(n_52));
  INVX1 g3907(.Y(n_53), .A(n_51));
  ADDFX1 g3908(.CO(n_51), .S(n_52), .A(in_26[1]), .B(in_20[1]), .CI(in_36[1]));
  ADDFX1 g3909(.CO(n_49), .S(n_50), .A(in_29[1]), .B(in_7[1]), .CI(in_30[0]));
  ADDFX1 g3910(.CO(n_47), .S(n_48), .A(in_22[0]), .B(n_5), .CI(n_2));
  ADDFX1 g3911(.CO(n_45), .S(n_46), .A(in_38[0]), .B(n_14), .CI(n_8));
  INVX1 g3912(.Y(n_44), .A(n_42));
  INVX1 g3913(.Y(n_43), .A(n_41));
  ADDFX1 g3914(.CO(n_41), .S(n_42), .A(in_16[1]), .B(in_6[1]), .CI(in_17[1]));
  ADDFX1 g3915(.CO(n_39), .S(n_40), .A(in_19[0]), .B(in_17[0]), .CI(in_6[0]));
  INVX1 g3916(.Y(n_38), .A(n_36));
  INVX1 g3917(.Y(n_37), .A(n_35));
  ADDFX1 g3918(.CO(n_35), .S(n_36), .A(in_31[0]), .B(in_32[0]), .CI(in_34[0]));
  ADDFX1 g3919(.CO(n_33), .S(n_34), .A(in_0[1]), .B(in_9[1]), .CI(n_7));
  ADDFX1 g3920(.CO(n_31), .S(n_32), .A(in_27[0]), .B(n_11), .CI(n_6));
  ADDFX1 g3921(.CO(n_29), .S(n_30), .A(in_15[0]), .B(n_9), .CI(n_13));
  ADDFX1 g3922(.CO(n_27), .S(n_28), .A(in_7[0]), .B(in_13[0]), .CI(n_12));
  ADDFX1 g3923(.CO(n_25), .S(n_26), .A(in_24[1]), .B(n_4), .CI(in_27[0]));
  XNOR2X1 g3924(.Y(n_24), .A(in_10[0]), .B(n_18));
  XOR2XL g3925(.Y(n_23), .A(in_10[2]), .B(n_18));
  OAI22X1 g3926(.Y(n_22), .A0(in_37[0]), .A1(n_17), .B0(in_25[0]), .B1(in_10[2]));
  OAI2BB1X1 g3927(.Y(n_21), .A0N(in_10[0]), .A1N(in_25[0]), .B0(n_20));
  OAI21XL g3928(.Y(n_20), .A0(in_10[0]), .A1(in_25[0]), .B0(in_37[0]));
  XNOR2X1 g3929(.Y(n_19), .A(in_33[1]), .B(in_3[1]));
  XNOR2X1 g3930(.Y(n_18), .A(in_37[0]), .B(in_25[0]));
  AND2XL g3932(.Y(n_17), .A(in_25[0]), .B(in_10[2]));
  NOR2XL g3933(.Y(n_16), .A(in_27[0]), .B(in_38[0]));
  NOR2BX1 g3934(.Y(n_15), .AN(in_3[1]), .B(in_33[1]));
  INVX1 g3935(.Y(n_14), .A(in_39[0]));
  INVX1 g3936(.Y(n_13), .A(in_18[0]));
  INVX1 g3937(.Y(n_12), .A(in_21[0]));
  INVX1 g3938(.Y(n_11), .A(in_23[0]));
  INVX1 g3939(.Y(n_10), .A(in_4[0]));
  INVX1 g3940(.Y(n_9), .A(in_12[0]));
  INVX1 g3941(.Y(n_8), .A(in_5[0]));
  INVX1 g3943(.Y(n_7), .A(in_28[1]));
  INVX1 g3944(.Y(n_6), .A(in_35[0]));
  INVX1 g3945(.Y(n_5), .A(in_41[0]));
  INVX1 g3946(.Y(n_4), .A(in_8[1]));
  INVX1 g3947(.Y(n_3), .A(in_19[1]));
  INVX1 g3948(.Y(n_2), .A(in_40[0]));
  CLKXOR2X1 g2(.Y(n_0), .A(in_27[0]), .B(in_38[0]));
endmodule

module WALLACE_CSA_DUMMY_OP109_group_109822_6312(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, out_0);
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [2:0] in_5;
input   [6:0] in_6;
input   [4:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [2:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [2:0] in_38;
output  [9:0] out_0;
wire  n_104, n_101, n_99, n_98, n_97, n_96, n_95, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_81, n_80, n_79, n_78, n_77, n_76, 
    n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, 
    n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, 
    n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_1;
wire   [9:0] out_0;
wire   [1:0] in_37;
wire   [1:0] in_33;
wire   [1:0] in_27;
wire   [1:0] in_25;
wire   [1:0] in_22;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_6;
wire   [2:0] in_38;
wire   [2:0] in_24;
wire   [2:0] in_5;
wire   [2:0] in_3;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_7;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  OA21X1 g2993(.Y(out_0[5]), .A0(n_89), .A1(n_104), .B0(out_0[9]));
  NAND2X1 g2994(.Y(out_0[9]), .A(n_89), .B(n_104));
  ADDFX1 g2995(.CO(n_104), .S(out_0[4]), .A(n_90), .B(n_97), .CI(n_101));
  ADDFX1 g2996(.CO(n_101), .S(out_0[3]), .A(n_98), .B(n_95), .CI(n_99));
  ADDFX1 g2997(.CO(n_99), .S(out_0[2]), .A(n_85), .B(n_93), .CI(n_96));
  ADDFX1 g2998(.CO(n_97), .S(n_98), .A(n_77), .B(n_87), .CI(n_91));
  ADDFX1 g2999(.CO(n_95), .S(n_96), .A(n_79), .B(n_78), .CI(n_92));
  ADDFX1 g3000(.CO(n_93), .S(out_0[1]), .A(n_81), .B(n_80), .CI(n_86));
  ADDFX1 g3001(.CO(n_91), .S(n_92), .A(n_61), .B(n_75), .CI(n_84));
  OAI2BB1X1 g3002(.Y(n_90), .A0N(n_73), .A1N(n_88), .B0(n_89));
  OR2X1 g3003(.Y(n_89), .A(n_73), .B(n_88));
  ADDFX1 g3004(.CO(n_88), .S(n_87), .A(n_74), .B(n_57), .CI(n_83));
  ADDFX1 g3005(.CO(n_85), .S(n_86), .A(n_71), .B(n_62), .CI(n_76));
  ADDFX1 g3006(.CO(n_83), .S(n_84), .A(n_55), .B(n_65), .CI(n_67));
  ADDFX1 g3007(.CO(n_81), .S(out_0[0]), .A(n_60), .B(n_54), .CI(n_72));
  ADDFX1 g3008(.CO(n_79), .S(n_80), .A(n_56), .B(n_68), .CI(n_64));
  ADDFX1 g3009(.CO(n_77), .S(n_78), .A(n_69), .B(n_63), .CI(n_58));
  ADDFX1 g3010(.CO(n_75), .S(n_76), .A(n_59), .B(n_66), .CI(n_53));
  OAI2BB1X1 g3011(.Y(n_74), .A0N(n_52), .A1N(n_70), .B0(n_73));
  OR2X1 g3012(.Y(n_73), .A(n_52), .B(n_70));
  ADDFX1 g3013(.CO(n_71), .S(n_72), .A(n_38), .B(n_26), .CI(n_46));
  ADDFX1 g3014(.CO(n_70), .S(n_69), .A(n_21), .B(n_41), .CI(n_47));
  ADDFX1 g3015(.CO(n_67), .S(n_68), .A(n_17), .B(n_49), .CI(n_19));
  ADDFX1 g3016(.CO(n_65), .S(n_66), .A(n_29), .B(n_33), .CI(n_22));
  ADDFX1 g3017(.CO(n_63), .S(n_64), .A(n_36), .B(n_42), .CI(n_48));
  ADDFX1 g3018(.CO(n_61), .S(n_62), .A(n_25), .B(n_45), .CI(n_44));
  ADDFX1 g3019(.CO(n_59), .S(n_60), .A(n_20), .B(n_34), .CI(n_50));
  ADDFX1 g3020(.CO(n_57), .S(n_58), .A(n_35), .B(n_43), .CI(n_51));
  ADDFX1 g3021(.CO(n_55), .S(n_56), .A(n_37), .B(n_31), .CI(n_23));
  ADDFX1 g3022(.CO(n_53), .S(n_54), .A(n_24), .B(n_32), .CI(n_30));
  ADDFX1 g3023(.CO(n_52), .S(n_51), .A(n_2), .B(n_1), .CI(n_18));
  ADDFX1 g3024(.CO(n_49), .S(n_50), .A(in_19[0]), .B(in_22[0]), .CI(n_15));
  ADDFX1 g3025(.CO(n_47), .S(n_48), .A(in_9[1]), .B(in_24[1]), .CI(n_6));
  ADDFX1 g3026(.CO(n_45), .S(n_46), .A(in_6[0]), .B(in_8[0]), .CI(in_15[0]));
  ADDFX1 g3027(.CO(n_43), .S(n_44), .A(n_4), .B(in_14[1]), .CI(n_13));
  INVX1 g3028(.Y(n_42), .A(n_40));
  INVX1 g3029(.Y(n_41), .A(n_39));
  ADDFX1 g3030(.CO(n_39), .S(n_40), .A(in_4[1]), .B(in_1[1]), .CI(in_35[1]));
  ADDFX1 g3031(.CO(n_37), .S(n_38), .A(in_27[0]), .B(n_7), .CI(n_16));
  ADDFX1 g3032(.CO(n_35), .S(n_36), .A(in_16[1]), .B(n_5), .CI(in_38[1]));
  ADDFX1 g3033(.CO(n_33), .S(n_34), .A(in_23[0]), .B(n_3), .CI(n_8));
  ADDFX1 g3034(.CO(n_31), .S(n_32), .A(in_25[0]), .B(n_10), .CI(in_33[0]));
  INVX1 g3035(.Y(n_30), .A(n_28));
  INVX1 g3036(.Y(n_29), .A(n_27));
  ADDFX1 g3037(.CO(n_27), .S(n_28), .A(in_2[0]), .B(in_7[0]), .CI(in_36[0]));
  ADDFX1 g3038(.CO(n_25), .S(n_26), .A(n_12), .B(n_14), .CI(in_14[0]));
  ADDFX1 g3039(.CO(n_23), .S(n_24), .A(in_11[0]), .B(n_11), .CI(in_37[0]));
  ADDFX1 g3040(.CO(n_21), .S(n_22), .A(in_3[1]), .B(in_5[1]), .CI(in_10[1]));
  OAI2BB1X1 g3041(.Y(n_20), .A0N(in_20[0]), .A1N(n_9), .B0(n_17));
  XOR2XL g3042(.Y(n_19), .A(in_30[1]), .B(in_6[1]));
  NOR2X1 g3043(.Y(n_18), .A(in_30[1]), .B(in_6[1]));
  OR2X1 g3044(.Y(n_17), .A(in_20[0]), .B(n_9));
  INVX1 g3045(.Y(n_16), .A(in_34[0]));
  INVX1 g3046(.Y(n_15), .A(in_32[0]));
  INVX1 g3047(.Y(n_14), .A(in_28[0]));
  INVX1 g3048(.Y(n_13), .A(in_15[1]));
  INVX1 g3049(.Y(n_12), .A(in_17[0]));
  INVX1 g3050(.Y(n_11), .A(in_13[0]));
  INVX1 g3051(.Y(n_10), .A(in_31[0]));
  INVX1 g3052(.Y(n_9), .A(in_21[0]));
  INVX1 g3053(.Y(n_8), .A(in_29[0]));
  INVX1 g3054(.Y(n_7), .A(in_0[0]));
  INVX1 g3055(.Y(n_6), .A(in_12[1]));
  INVX1 g3056(.Y(n_5), .A(in_18[1]));
  INVX1 g3057(.Y(n_4), .A(in_8[1]));
  INVX1 g3058(.Y(n_3), .A(in_26[0]));
  INVX1 g3059(.Y(n_2), .A(in_19[0]));
  INVX1 g3060(.Y(n_1), .A(in_23[0]));
endmodule

module WALLACE_CSA_DUMMY_OP109_group_109822(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, out_0);
input  in_39, in_40, in_43, in_44, in_53, in_58, in_60;
input   [4:0] in_0;
input   [2:0] in_1;
input   [4:0] in_2;
input   [1:0] in_3;
input   [1:0] in_4;
input   [9:0] in_5;
input   [7:0] in_6;
input   [6:0] in_7;
input   [6:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [4:0] in_24;
input   [2:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [5:0] in_34;
input   [5:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [2:0] in_38;
input   [2:0] in_41;
input   [1:0] in_42;
input   [1:0] in_45;
input   [1:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [1:0] in_49;
input   [4:0] in_50;
input   [4:0] in_51;
input   [1:0] in_52;
input   [1:0] in_54;
input   [1:0] in_55;
input   [1:0] in_56;
input   [1:0] in_57;
input   [1:0] in_59;
input   [1:0] in_61;
input   [1:0] in_62;
input   [4:0] in_63;
input   [1:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [2:0] in_67;
input   [1:0] in_68;
input   [1:0] in_69;
input   [4:0] in_70;
input   [4:0] in_71;
input   [2:0] in_72;
input   [1:0] in_73;
input   [1:0] in_74;
input   [4:0] in_75;
input   [3:0] in_76;
input   [1:0] in_77;
input   [1:0] in_78;
output  [9:0] out_0;
wire  n_220, n_218, n_216, n_214, n_212, n_210, n_208, n_207, n_206, n_204, 
    n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 
    n_193, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
    n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, 
    n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
    n_162, n_161, n_160, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
    n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, 
    n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, 
    n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, 
    n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
    n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, 
    n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, 
    n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
    n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_1, n_0, in_60, in_58, in_53, in_44, in_43, in_40, in_39;
wire   [9:0] out_0;
wire   [3:0] in_76;
wire   [5:0] in_35;
wire   [5:0] in_34;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [6:0] in_8;
wire   [6:0] in_7;
wire   [7:0] in_6;
wire   [9:0] in_5;
wire   [1:0] in_78;
wire   [1:0] in_77;
wire   [1:0] in_74;
wire   [1:0] in_73;
wire   [1:0] in_69;
wire   [1:0] in_68;
wire   [1:0] in_64;
wire   [1:0] in_62;
wire   [1:0] in_61;
wire   [1:0] in_59;
wire   [1:0] in_57;
wire   [1:0] in_56;
wire   [1:0] in_55;
wire   [1:0] in_54;
wire   [1:0] in_52;
wire   [1:0] in_49;
wire   [1:0] in_46;
wire   [1:0] in_45;
wire   [1:0] in_42;
wire   [1:0] in_37;
wire   [1:0] in_4;
wire   [1:0] in_3;
wire   [2:0] in_72;
wire   [2:0] in_67;
wire   [2:0] in_41;
wire   [2:0] in_38;
wire   [2:0] in_25;
wire   [2:0] in_1;
wire   [4:0] in_75;
wire   [4:0] in_71;
wire   [4:0] in_70;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_63;
wire   [4:0] in_51;
wire   [4:0] in_50;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_36;
wire   [4:0] in_24;
wire   [4:0] in_2;
wire   [4:0] in_0;
  INVX1 g2744(.Y(out_0[8]), .A(n_220));
  ADDFX1 g2745(.CO(out_0[9]), .S(n_220), .A(in_5[8]), .B(n_0), .CI(n_218));
  INVX1 g2746(.Y(n_218), .A(n_216));
  ADDFX1 g2747(.CO(n_216), .S(out_0[7]), .A(n_0), .B(n_190), .CI(n_214));
  ADDFX1 g2748(.CO(n_214), .S(out_0[6]), .A(n_206), .B(n_193), .CI(n_212));
  ADDFX1 g2749(.CO(n_212), .S(out_0[5]), .A(n_202), .B(n_207), .CI(n_210));
  ADDFX1 g2750(.CO(n_210), .S(out_0[4]), .A(n_200), .B(n_208), .CI(n_203));
  ADDFX1 g2751(.CO(n_208), .S(out_0[3]), .A(n_201), .B(n_195), .CI(n_204));
  ADDFX1 g2752(.CO(n_206), .S(n_207), .A(n_180), .B(n_198), .CI(n_188));
  ADDFX1 g2753(.CO(n_204), .S(out_0[2]), .A(n_176), .B(n_191), .CI(n_197));
  ADDFX1 g2754(.CO(n_202), .S(n_203), .A(n_181), .B(n_194), .CI(n_199));
  ADDFX1 g2755(.CO(n_200), .S(n_201), .A(n_182), .B(n_185), .CI(n_196));
  ADDFX1 g2756(.CO(n_198), .S(n_199), .A(n_186), .B(n_184), .CI(in_5[4]));
  ADDFX1 g2757(.CO(n_196), .S(n_197), .A(n_179), .B(n_183), .CI(in_5[2]));
  ADDFX1 g2758(.CO(n_194), .S(n_195), .A(n_178), .B(n_187), .CI(in_5[3]));
  OAI2BB1X1 g2759(.Y(n_193), .A0N(in_5[6]), .A1N(n_189), .B0(n_190));
  ADDFX1 g2760(.CO(n_191), .S(out_0[1]), .A(n_147), .B(n_158), .CI(n_177));
  OR2X1 g2761(.Y(n_190), .A(in_5[6]), .B(n_189));
  ADDFX1 g2762(.CO(n_189), .S(n_188), .A(n_156), .B(n_174), .CI(in_5[5]));
  ADDFX1 g2763(.CO(n_186), .S(n_187), .A(n_172), .B(n_168), .CI(n_161));
  ADDFX1 g2764(.CO(n_184), .S(n_185), .A(n_162), .B(n_165), .CI(n_167));
  ADDFX1 g2765(.CO(n_182), .S(n_183), .A(n_173), .B(n_163), .CI(n_169));
  ADDFX1 g2766(.CO(n_180), .S(n_181), .A(n_166), .B(n_164), .CI(n_175));
  ADDFX1 g2767(.CO(n_178), .S(n_179), .A(n_146), .B(n_143), .CI(n_170));
  ADDFX1 g2768(.CO(n_176), .S(n_177), .A(n_141), .B(n_171), .CI(in_5[1]));
  ADDFX1 g2769(.CO(n_174), .S(n_175), .A(n_150), .B(n_160), .CI(n_157));
  ADDFX1 g2770(.CO(n_172), .S(n_173), .A(n_116), .B(n_152), .CI(n_144));
  ADDFX1 g2771(.CO(n_170), .S(n_171), .A(n_135), .B(n_153), .CI(n_145));
  ADDFX1 g2772(.CO(n_168), .S(n_169), .A(n_123), .B(n_134), .CI(n_155));
  ADDFX1 g2773(.CO(n_166), .S(n_167), .A(n_122), .B(n_137), .CI(n_151));
  ADDFX1 g2774(.CO(n_164), .S(n_165), .A(n_132), .B(n_148), .CI(n_142));
  ADDFX1 g2775(.CO(n_162), .S(n_163), .A(n_133), .B(n_140), .CI(n_149));
  ADDFX1 g2776(.CO(n_160), .S(n_161), .A(n_131), .B(n_154), .CI(n_82));
  ADDFX1 g2777(.CO(n_158), .S(out_0[0]), .A(n_119), .B(n_139), .CI(in_5[0]));
  ADDFX1 g2778(.CO(n_156), .S(n_157), .A(n_130), .B(n_136), .CI(n_14));
  ADDFX1 g2779(.CO(n_154), .S(n_155), .A(n_108), .B(n_128), .CI(n_126));
  ADDFX1 g2780(.CO(n_152), .S(n_153), .A(n_86), .B(n_120), .CI(n_129));
  ADDFX1 g2781(.CO(n_150), .S(n_151), .A(n_114), .B(n_124), .CI(in_6[3]));
  ADDFX1 g2782(.CO(n_148), .S(n_149), .A(n_115), .B(n_90), .CI(n_125));
  ADDFX1 g2783(.CO(n_146), .S(n_147), .A(n_118), .B(n_117), .CI(n_138));
  ADDFX1 g2784(.CO(n_144), .S(n_145), .A(n_109), .B(n_99), .CI(n_127));
  ADDFX1 g2785(.CO(n_142), .S(n_143), .A(n_85), .B(n_110), .CI(n_83));
  ADDFX1 g2786(.CO(n_140), .S(n_141), .A(n_111), .B(n_113), .CI(n_91));
  ADDFX1 g2787(.CO(n_138), .S(n_139), .A(n_87), .B(n_101), .CI(n_121));
  ADDFX1 g2788(.CO(n_136), .S(n_137), .A(n_104), .B(n_94), .CI(n_84));
  ADDFX1 g2789(.CO(n_134), .S(n_135), .A(n_88), .B(n_100), .CI(n_93));
  ADDFX1 g2790(.CO(n_132), .S(n_133), .A(n_95), .B(n_92), .CI(n_112));
  ADDFX1 g2791(.CO(n_130), .S(n_131), .A(n_19), .B(n_24), .CI(n_102));
  ADDFX1 g2792(.CO(n_128), .S(n_129), .A(n_48), .B(n_64), .CI(n_106));
  ADDFX1 g2793(.CO(n_126), .S(n_127), .A(n_72), .B(n_44), .CI(n_97));
  ADDFX1 g2794(.CO(n_124), .S(n_125), .A(n_54), .B(n_96), .CI(n_103));
  ADDFX1 g2795(.CO(n_122), .S(n_123), .A(n_80), .B(n_98), .CI(n_105));
  ADDFX1 g2796(.CO(n_120), .S(n_121), .A(n_73), .B(in_6[0]), .CI(n_107));
  ADDFX1 g2797(.CO(n_118), .S(n_119), .A(n_35), .B(n_63), .CI(n_89));
  ADDFX1 g2798(.CO(n_116), .S(n_117), .A(n_67), .B(n_29), .CI(n_81));
  ADDFX1 g2799(.CO(n_114), .S(n_115), .A(n_11), .B(n_66), .CI(n_68));
  ADDFX1 g2800(.CO(n_112), .S(n_113), .A(n_61), .B(n_43), .CI(n_23));
  ADDFX1 g2801(.CO(n_110), .S(n_111), .A(n_69), .B(n_31), .CI(n_55));
  ADDFX1 g2802(.CO(n_108), .S(n_109), .A(n_58), .B(n_76), .CI(n_26));
  ADDFX1 g2803(.CO(n_106), .S(n_107), .A(in_30[0]), .B(n_5), .CI(n_57));
  ADDFX1 g2804(.CO(n_104), .S(n_105), .A(n_42), .B(n_50), .CI(n_60));
  ADDFX1 g2805(.CO(n_102), .S(n_103), .A(in_76[0]), .B(n_20), .CI(n_78));
  ADDFX1 g2806(.CO(n_100), .S(n_101), .A(n_77), .B(n_65), .CI(n_45));
  ADDFX1 g2807(.CO(n_98), .S(n_99), .A(n_32), .B(n_34), .CI(n_62));
  ADDFX1 g2808(.CO(n_96), .S(n_97), .A(in_20[1]), .B(n_79), .CI(n_56));
  ADDFX1 g2809(.CO(n_94), .S(n_95), .A(n_74), .B(n_52), .CI(n_36));
  ADDFX1 g2810(.CO(n_92), .S(n_93), .A(n_75), .B(n_37), .CI(n_41));
  ADDFX1 g2811(.CO(n_90), .S(n_91), .A(n_53), .B(n_51), .CI(in_6[1]));
  ADDFX1 g2812(.CO(n_88), .S(n_89), .A(n_59), .B(n_27), .CI(n_49));
  ADDFX1 g2813(.CO(n_86), .S(n_87), .A(in_32[0]), .B(n_33), .CI(n_39));
  ADDFX1 g2814(.CO(n_84), .S(n_85), .A(n_22), .B(n_40), .CI(n_30));
  ADDFX1 g2815(.CO(n_82), .S(n_83), .A(n_25), .B(n_28), .CI(in_6[2]));
  ADDFX1 g2816(.CO(n_80), .S(n_81), .A(n_16), .B(in_34[1]), .CI(n_38));
  INVX1 g2817(.Y(n_79), .A(n_71));
  INVX1 g2818(.Y(n_78), .A(n_70));
  ADDFX1 g2819(.CO(n_76), .S(n_77), .A(in_27[0]), .B(in_53), .CI(in_64[0]));
  ADDFX1 g2820(.CO(n_74), .S(n_75), .A(n_9), .B(n_1), .CI(in_62[1]));
  ADDFX1 g2821(.CO(n_72), .S(n_73), .A(in_12[0]), .B(in_34[0]), .CI(in_76[0]));
  ADDFX1 g2822(.CO(n_70), .S(n_71), .A(in_16[1]), .B(in_22[1]), .CI(n_18));
  ADDFX1 g2823(.CO(n_68), .S(n_69), .A(in_1[1]), .B(in_56[1]), .CI(in_9[0]));
  ADDFX1 g2824(.CO(n_66), .S(n_67), .A(in_10[1]), .B(in_73[1]), .CI(in_78[0]));
  ADDFX1 g2825(.CO(n_64), .S(n_65), .A(in_31[0]), .B(n_15), .CI(in_54[0]));
  ADDFX1 g2826(.CO(n_62), .S(n_63), .A(in_39), .B(in_57[0]), .CI(n_6));
  ADDFX1 g2827(.CO(n_60), .S(n_61), .A(in_74[1]), .B(n_12), .CI(in_77[1]));
  ADDFX1 g2828(.CO(n_58), .S(n_59), .A(in_11[0]), .B(in_58), .CI(in_9[0]));
  ADDFX1 g2829(.CO(n_56), .S(n_57), .A(n_4), .B(n_3), .CI(n_21));
  INVX1 g2830(.Y(n_55), .A(n_47));
  INVX1 g2831(.Y(n_54), .A(n_46));
  ADDFX1 g2832(.CO(n_52), .S(n_53), .A(in_25[1]), .B(in_38[1]), .CI(in_69[1]));
  ADDFX1 g2833(.CO(n_50), .S(n_51), .A(in_46[1]), .B(in_52[1]), .CI(in_61[1]));
  ADDFX1 g2834(.CO(n_48), .S(n_49), .A(in_60), .B(in_19[0]), .CI(n_7));
  ADDFX1 g2835(.CO(n_46), .S(n_47), .A(in_48[1]), .B(in_47[1]), .CI(in_50[1]));
  ADDFX1 g2836(.CO(n_44), .S(n_45), .A(in_17[0]), .B(in_40), .CI(in_44));
  ADDFX1 g2837(.CO(n_42), .S(n_43), .A(in_17[0]), .B(in_68[1]), .CI(in_55[0]));
  ADDFX1 g2838(.CO(n_40), .S(n_41), .A(in_57[0]), .B(n_10), .CI(n_17));
  ADDFX1 g2839(.CO(n_38), .S(n_39), .A(in_13[0]), .B(n_2), .CI(in_55[0]));
  ADDFX1 g2840(.CO(n_36), .S(n_37), .A(in_23[1]), .B(n_13), .CI(in_72[1]));
  ADDFX1 g2841(.CO(n_34), .S(n_35), .A(in_10[0]), .B(in_33[0]), .CI(in_78[0]));
  ADDFX1 g2842(.CO(n_32), .S(n_33), .A(in_37[0]), .B(in_26[0]), .CI(in_49[0]));
  ADDFX1 g2843(.CO(n_30), .S(n_31), .A(in_45[1]), .B(in_59[1]), .CI(in_67[1]));
  ADDFX1 g2844(.CO(n_28), .S(n_29), .A(in_41[1]), .B(in_7[1]), .CI(in_18[1]));
  ADDFX1 g2845(.CO(n_26), .S(n_27), .A(in_15[0]), .B(in_42[0]), .CI(in_43));
  ADDFX1 g2846(.CO(n_24), .S(n_25), .A(in_28[2]), .B(in_35[2]), .CI(n_8));
  ADDFX1 g2847(.CO(n_22), .S(n_23), .A(in_4[1]), .B(in_3[1]), .CI(in_19[0]));
  XNOR2X1 g2848(.Y(n_21), .A(in_29[0]), .B(in_14[0]));
  XOR2XL g2849(.Y(n_20), .A(in_14[0]), .B(in_7[2]));
  NOR2X1 g2850(.Y(n_19), .A(in_14[0]), .B(in_7[2]));
  NAND2BX1 g2851(.Y(n_18), .AN(in_29[0]), .B(in_14[0]));
  INVX1 g2852(.Y(n_17), .A(in_75[1]));
  INVX1 g2853(.Y(n_16), .A(in_32[1]));
  INVX1 g2854(.Y(n_15), .A(in_0[0]));
  INVX1 g2855(.Y(n_14), .A(in_6[4]));
  INVX1 g2856(.Y(n_13), .A(in_70[1]));
  INVX1 g2857(.Y(n_12), .A(in_66[1]));
  INVX1 g2858(.Y(n_11), .A(in_18[2]));
  INVX1 g2859(.Y(n_10), .A(in_71[1]));
  INVX1 g2860(.Y(n_9), .A(in_2[1]));
  INVX1 g2861(.Y(n_8), .A(in_34[2]));
  INVX1 g2862(.Y(n_7), .A(in_65[0]));
  INVX1 g2863(.Y(n_6), .A(in_63[0]));
  INVX1 g2864(.Y(n_5), .A(in_24[0]));
  INVX1 g2865(.Y(n_4), .A(in_8[0]));
  INVX1 g2866(.Y(n_3), .A(in_21[0]));
  INVX1 g2867(.Y(n_2), .A(in_51[0]));
  INVX1 g2868(.Y(n_1), .A(in_36[1]));
  INVX1 g2869(.Y(n_0), .A(in_5[7]));
endmodule

module WALLACE_CSA_DUMMY_OP125_group_106193(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, out_0);
input  in_4;
input   [2:0] in_0;
input   [4:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [1:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [4:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [1:0] in_18;
input   [1:0] in_19;
input   [4:0] in_20;
input   [2:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [1:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [2:0] in_40;
input   [2:0] in_41;
output  [9:0] out_0;
wire  n_124, n_122, n_120, n_118, n_117, n_116, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_92, n_91, n_90, n_89, n_88, 
    n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, 
    n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, 
    n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, 
    n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_0, in_4;
wire   [9:0] out_0;
wire   [1:0] in_28;
wire   [1:0] in_19;
wire   [1:0] in_18;
wire   [1:0] in_5;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_15;
wire   [4:0] in_1;
wire   [2:0] in_41;
wire   [2:0] in_40;
wire   [2:0] in_37;
wire   [2:0] in_21;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3682(.Y(out_0[9]), .A(n_124));
  ADDFX1 g3683(.CO(n_124), .S(out_0[5]), .A(n_98), .B(n_110), .CI(n_122));
  ADDFX1 g3684(.CO(n_122), .S(out_0[4]), .A(n_111), .B(n_116), .CI(n_120));
  ADDFX1 g3685(.CO(n_120), .S(out_0[3]), .A(n_112), .B(n_117), .CI(n_118));
  ADDFX1 g3686(.CO(n_118), .S(out_0[2]), .A(n_107), .B(n_114), .CI(n_113));
  ADDFX1 g3687(.CO(n_116), .S(n_117), .A(n_101), .B(n_109), .CI(n_106));
  ADDFX1 g3688(.CO(n_114), .S(out_0[1]), .A(n_92), .B(n_89), .CI(n_105));
  ADDFX1 g3689(.CO(n_112), .S(n_113), .A(n_103), .B(n_87), .CI(n_104));
  ADDFX1 g3690(.CO(n_110), .S(n_111), .A(n_99), .B(n_100), .CI(n_108));
  ADDFX1 g3691(.CO(n_108), .S(n_109), .A(n_85), .B(n_86), .CI(n_102));
  ADDFX1 g3692(.CO(n_106), .S(n_107), .A(n_94), .B(n_97), .CI(n_88));
  ADDFX1 g3693(.CO(n_104), .S(n_105), .A(n_76), .B(n_91), .CI(n_95));
  ADDFX1 g3694(.CO(n_102), .S(n_103), .A(n_67), .B(n_83), .CI(n_90));
  ADDFX1 g3695(.CO(n_100), .S(n_101), .A(n_82), .B(n_66), .CI(n_96));
  ADDHX1 g3696(.CO(n_98), .S(n_99), .A(n_49), .B(n_84));
  ADDFX1 g3697(.CO(n_96), .S(n_97), .A(n_64), .B(n_78), .CI(n_75));
  ADDFX1 g3698(.CO(n_94), .S(n_95), .A(n_57), .B(n_73), .CI(n_80));
  ADDFX1 g3699(.CO(n_92), .S(out_0[0]), .A(n_71), .B(n_81), .CI(n_77));
  ADDFX1 g3700(.CO(n_90), .S(n_91), .A(n_58), .B(n_79), .CI(n_70));
  ADDFX1 g3701(.CO(n_88), .S(n_89), .A(n_65), .B(n_63), .CI(n_69));
  ADDFX1 g3702(.CO(n_86), .S(n_87), .A(n_72), .B(n_62), .CI(n_68));
  ADDFX1 g3703(.CO(n_84), .S(n_85), .A(n_60), .B(n_74), .CI(n_0));
  ADDFX1 g3704(.CO(n_82), .S(n_83), .A(n_35), .B(n_61), .CI(n_56));
  ADDFX1 g3705(.CO(n_80), .S(n_81), .A(n_33), .B(n_53), .CI(n_40));
  ADDFX1 g3706(.CO(n_78), .S(n_79), .A(n_22), .B(n_39), .CI(n_52));
  ADDFX1 g3707(.CO(n_76), .S(n_77), .A(n_23), .B(in_2[0]), .CI(n_59));
  ADDFX1 g3708(.CO(n_74), .S(n_75), .A(n_45), .B(n_28), .CI(n_26));
  ADDFX1 g3709(.CO(n_72), .S(n_73), .A(n_50), .B(n_37), .CI(n_31));
  ADDFX1 g3710(.CO(n_70), .S(n_71), .A(n_55), .B(n_42), .CI(n_51));
  ADDFX1 g3711(.CO(n_68), .S(n_69), .A(n_44), .B(n_27), .CI(in_2[1]));
  ADDFX1 g3712(.CO(n_66), .S(n_67), .A(n_43), .B(n_48), .CI(n_17));
  ADDFX1 g3713(.CO(n_64), .S(n_65), .A(n_54), .B(n_41), .CI(n_32));
  ADDFX1 g3714(.CO(n_62), .S(n_63), .A(n_46), .B(n_29), .CI(n_36));
  ADDFX1 g3715(.CO(n_60), .S(n_61), .A(in_35[2]), .B(n_10), .CI(n_30));
  ADDFX1 g3716(.CO(n_58), .S(n_59), .A(in_10[0]), .B(in_3[0]), .CI(n_38));
  ADDFX1 g3718(.CO(n_56), .S(n_57), .A(n_3), .B(in_7[1]), .CI(in_14[1]));
  ADDFX1 g3719(.CO(n_54), .S(n_55), .A(in_7[0]), .B(n_18), .CI(n_7));
  ADDFX1 g3720(.CO(n_52), .S(n_53), .A(n_15), .B(in_8[0]), .CI(n_6));
  ADDFX1 g3721(.CO(n_50), .S(n_51), .A(in_9[0]), .B(n_19), .CI(in_37[0]));
  NOR2X1 g3722(.Y(n_49), .A(in_35[2]), .B(n_47));
  INVX1 g3723(.Y(n_48), .A(n_34));
  INVX1 g3724(.Y(n_46), .A(n_25));
  INVX1 g3725(.Y(n_45), .A(n_24));
  ADDFX1 g3726(.CO(n_43), .S(n_44), .A(in_12[0]), .B(n_11), .CI(in_37[0]));
  ADDFX1 g3727(.CO(n_41), .S(n_42), .A(in_4), .B(n_2), .CI(in_19[0]));
  ADDFX1 g3728(.CO(n_39), .S(n_40), .A(n_12), .B(in_12[0]), .CI(n_8));
  ADDFX1 g3729(.CO(n_37), .S(n_38), .A(in_6[0]), .B(in_14[0]), .CI(n_21));
  ADDFX1 g3730(.CO(n_35), .S(n_36), .A(n_13), .B(in_40[1]), .CI(n_14));
  ADDFX1 g3731(.CO(n_47), .S(n_34), .A(in_9[0]), .B(in_34[0]), .CI(in_14[2]));
  ADDFX1 g3732(.CO(n_32), .S(n_33), .A(in_28[0]), .B(in_18[0]), .CI(in_34[0]));
  ADDFX1 g3733(.CO(n_30), .S(n_31), .A(in_0[1]), .B(n_5), .CI(in_41[1]));
  ADDFX1 g3734(.CO(n_28), .S(n_29), .A(in_5[1]), .B(n_4), .CI(n_9));
  ADDFX1 g3735(.CO(n_26), .S(n_27), .A(in_21[1]), .B(n_16), .CI(n_20));
  ADDFX1 g3736(.CO(n_24), .S(n_25), .A(in_16[1]), .B(in_26[1]), .CI(in_27[1]));
  OAI21X1 g3737(.Y(n_23), .A0(in_20[0]), .A1(in_15[0]), .B0(n_22));
  NAND2X1 g3738(.Y(n_22), .A(in_20[0]), .B(in_15[0]));
  INVX1 g3739(.Y(n_21), .A(in_39[0]));
  INVX1 g3740(.Y(n_20), .A(in_32[1]));
  INVX1 g3741(.Y(n_19), .A(in_25[0]));
  INVX1 g3742(.Y(n_18), .A(in_17[0]));
  INVX1 g3743(.Y(n_17), .A(in_2[2]));
  INVX1 g3744(.Y(n_16), .A(in_22[1]));
  INVX1 g3745(.Y(n_15), .A(in_11[0]));
  INVX1 g3746(.Y(n_14), .A(in_3[1]));
  INVX1 g3747(.Y(n_13), .A(in_36[1]));
  INVX1 g3748(.Y(n_12), .A(in_13[0]));
  INVX1 g3749(.Y(n_11), .A(in_24[1]));
  INVX1 g3750(.Y(n_10), .A(in_7[2]));
  INVX1 g3752(.Y(n_9), .A(in_30[1]));
  INVX1 g3753(.Y(n_8), .A(in_33[0]));
  INVX1 g3754(.Y(n_7), .A(in_29[0]));
  INVX1 g3755(.Y(n_6), .A(in_31[0]));
  INVX1 g3756(.Y(n_5), .A(in_38[1]));
  INVX1 g3757(.Y(n_4), .A(in_23[1]));
  INVX1 g3758(.Y(n_3), .A(in_10[1]));
  INVX1 g3759(.Y(n_2), .A(in_1[0]));
  XOR2XL g2(.Y(n_0), .A(in_35[2]), .B(n_47));
endmodule

module WALLACE_CSA_DUMMY_OP127_group_109819(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    out_0);
input  in_23;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [6:0] in_4;
input   [4:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [1:0] in_19;
input   [2:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [1:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [4:0] in_37;
output  [9:0] out_0;
wire  n_112, n_110, n_108, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_23;
wire   [9:0] out_0;
wire   [1:0] in_32;
wire   [1:0] in_29;
wire   [1:0] in_28;
wire   [1:0] in_22;
wire   [1:0] in_19;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_4;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_21;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_5;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_36;
wire   [2:0] in_20;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3192(.Y(out_0[9]), .A(n_112));
  ADDFX1 g3193(.CO(n_112), .S(out_0[5]), .A(n_55), .B(n_102), .CI(n_110));
  ADDFX1 g3194(.CO(n_110), .S(out_0[4]), .A(n_103), .B(n_104), .CI(n_108));
  ADDFX1 g3195(.CO(n_108), .S(out_0[3]), .A(n_100), .B(n_105), .CI(n_106));
  ADDFX1 g3196(.CO(n_106), .S(out_0[2]), .A(n_92), .B(n_98), .CI(n_101));
  ADDFX1 g3197(.CO(n_104), .S(n_105), .A(n_85), .B(n_97), .CI(n_94));
  ADDFX1 g3198(.CO(n_102), .S(n_103), .A(n_57), .B(n_84), .CI(n_96));
  ADDFX1 g3199(.CO(n_100), .S(n_101), .A(n_88), .B(n_83), .CI(n_95));
  ADDFX1 g3200(.CO(n_98), .S(out_0[1]), .A(n_90), .B(n_89), .CI(n_93));
  ADDFX1 g3201(.CO(n_96), .S(n_97), .A(n_78), .B(n_86), .CI(n_82));
  ADDFX1 g3202(.CO(n_94), .S(n_95), .A(n_79), .B(n_80), .CI(n_87));
  ADDFX1 g3203(.CO(n_92), .S(n_93), .A(n_76), .B(n_71), .CI(n_81));
  ADDFX1 g3204(.CO(n_90), .S(out_0[0]), .A(n_63), .B(n_65), .CI(n_77));
  ADDFX1 g3205(.CO(n_88), .S(n_89), .A(n_67), .B(n_75), .CI(n_73));
  ADDFX1 g3206(.CO(n_86), .S(n_87), .A(n_66), .B(n_61), .CI(n_74));
  ADDFX1 g3207(.CO(n_84), .S(n_85), .A(n_56), .B(n_60), .CI(n_68));
  ADDFX1 g3208(.CO(n_82), .S(n_83), .A(n_72), .B(n_69), .CI(n_70));
  ADDFX1 g3209(.CO(n_80), .S(n_81), .A(n_64), .B(n_59), .CI(n_62));
  ADDFX1 g3210(.CO(n_78), .S(n_79), .A(n_50), .B(n_44), .CI(n_58));
  ADDFX1 g3211(.CO(n_76), .S(n_77), .A(n_54), .B(n_31), .CI(n_41));
  ADDFX1 g3212(.CO(n_74), .S(n_75), .A(n_46), .B(n_25), .CI(n_29));
  ADDFX1 g3213(.CO(n_72), .S(n_73), .A(n_21), .B(n_39), .CI(n_40));
  ADDFX1 g3214(.CO(n_70), .S(n_71), .A(n_19), .B(n_30), .CI(n_45));
  ADDFX1 g3215(.CO(n_68), .S(n_69), .A(n_15), .B(n_38), .CI(n_18));
  ADDFX1 g3216(.CO(n_66), .S(n_67), .A(n_53), .B(n_34), .CI(n_3));
  ADDFX1 g3217(.CO(n_64), .S(n_65), .A(in_9[0]), .B(n_33), .CI(n_47));
  ADDFX1 g3218(.CO(n_62), .S(n_63), .A(n_23), .B(n_17), .CI(n_35));
  ADDFX1 g3219(.CO(n_60), .S(n_61), .A(n_24), .B(n_28), .CI(n_20));
  ADDFX1 g3220(.CO(n_58), .S(n_59), .A(n_16), .B(n_22), .CI(n_32));
  INVX1 g3221(.Y(n_57), .A(n_55));
  XNOR2X1 g3222(.Y(n_56), .A(n_13), .B(n_49));
  NOR2BX1 g3223(.Y(n_55), .AN(n_13), .B(n_49));
  INVX1 g3224(.Y(n_54), .A(n_52));
  INVX1 g3225(.Y(n_53), .A(n_51));
  ADDFX1 g3226(.CO(n_51), .S(n_52), .A(in_3[0]), .B(in_6[0]), .CI(in_27[0]));
  INVX1 g3227(.Y(n_50), .A(n_48));
  ADDFX1 g3228(.CO(n_49), .S(n_48), .A(in_8[2]), .B(in_14[0]), .CI(n_12));
  ADDFX1 g3229(.CO(n_46), .S(n_47), .A(in_14[0]), .B(in_13[0]), .CI(in_32[0]));
  INVX1 g3230(.Y(n_45), .A(n_43));
  INVX1 g3231(.Y(n_44), .A(n_42));
  ADDFX1 g3232(.CO(n_42), .S(n_43), .A(in_9[1]), .B(in_12[1]), .CI(n_14));
  ADDFX1 g3233(.CO(n_40), .S(n_41), .A(in_10[0]), .B(in_8[0]), .CI(in_15[0]));
  INVX1 g3234(.Y(n_39), .A(n_37));
  INVX1 g3235(.Y(n_38), .A(n_36));
  ADDFX1 g3236(.CO(n_36), .S(n_37), .A(in_2[1]), .B(in_34[1]), .CI(in_18[1]));
  ADDFX1 g3237(.CO(n_34), .S(n_35), .A(in_23), .B(n_10), .CI(n_11));
  ADDFX1 g3238(.CO(n_32), .S(n_33), .A(in_11[0]), .B(n_2), .CI(n_4));
  ADDFX1 g3239(.CO(n_30), .S(n_31), .A(in_29[0]), .B(in_36[0]), .CI(in_12[0]));
  INVX1 g3240(.Y(n_29), .A(n_27));
  INVX1 g3241(.Y(n_28), .A(n_26));
  ADDFX1 g3242(.CO(n_26), .S(n_27), .A(in_25[1]), .B(in_30[1]), .CI(in_37[1]));
  ADDFX1 g3243(.CO(n_24), .S(n_25), .A(in_16[1]), .B(in_19[1]), .CI(in_28[1]));
  ADDFX1 g3244(.CO(n_22), .S(n_23), .A(in_7[0]), .B(n_9), .CI(n_5));
  ADDFX1 g3245(.CO(n_20), .S(n_21), .A(in_0[1]), .B(n_6), .CI(n_1));
  ADDFX1 g3246(.CO(n_18), .S(n_19), .A(in_29[0]), .B(in_8[1]), .CI(in_15[1]));
  ADDFX1 g3247(.CO(n_16), .S(n_17), .A(in_5[0]), .B(in_4[0]), .CI(n_7));
  OAI2BB1X1 g3248(.Y(n_15), .A0N(in_20[2]), .A1N(n_8), .B0(n_13));
  XNOR2X1 g3249(.Y(n_14), .A(in_22[1]), .B(in_36[0]));
  NAND2BX1 g3250(.Y(n_13), .AN(in_20[2]), .B(in_4[0]));
  NAND2X1 g3251(.Y(n_12), .A(in_36[0]), .B(in_22[1]));
  INVX1 g3252(.Y(n_11), .A(in_24[0]));
  INVX1 g3253(.Y(n_10), .A(in_1[0]));
  INVX1 g3254(.Y(n_9), .A(in_31[0]));
  INVXL g3255(.Y(n_8), .A(in_4[0]));
  INVX1 g3256(.Y(n_7), .A(in_26[0]));
  INVX1 g3257(.Y(n_6), .A(in_21[1]));
  INVX1 g3258(.Y(n_5), .A(in_35[0]));
  INVX1 g3259(.Y(n_4), .A(in_33[0]));
  INVX1 g3260(.Y(n_3), .A(in_10[1]));
  INVX1 g3261(.Y(n_2), .A(in_17[0]));
  INVX1 g3262(.Y(n_1), .A(in_7[1]));
endmodule

module WALLACE_CSA_DUMMY_OP130_group_109827(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, out_0);
input  in_5, in_17, in_32;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [1:0] in_4;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [1:0] in_16;
input   [2:0] in_18;
input   [2:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [1:0] in_33;
input   [4:0] in_34;
input   [2:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
output  [9:0] out_0;
wire  n_104, n_101, n_99, n_98, n_97, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, 
    n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, 
    n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, 
    n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_1, in_32, in_17, in_5;
wire   [9:0] out_0;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [1:0] in_41;
wire   [1:0] in_33;
wire   [1:0] in_31;
wire   [1:0] in_16;
wire   [1:0] in_4;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_34;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_35;
wire   [2:0] in_19;
wire   [2:0] in_18;
wire   [2:0] in_3;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  OA21X1 g3106(.Y(out_0[5]), .A0(n_91), .A1(n_104), .B0(out_0[9]));
  NAND2X1 g3107(.Y(out_0[9]), .A(n_91), .B(n_104));
  ADDFX1 g3108(.CO(n_104), .S(out_0[4]), .A(n_94), .B(n_97), .CI(n_101));
  ADDFX1 g3109(.CO(n_101), .S(out_0[3]), .A(n_92), .B(n_98), .CI(n_99));
  ADDFX1 g3110(.CO(n_99), .S(out_0[2]), .A(n_90), .B(n_93), .CI(n_95));
  ADDFX1 g3111(.CO(n_97), .S(n_98), .A(n_75), .B(n_89), .CI(n_87));
  ADDFX1 g3112(.CO(n_95), .S(out_0[1]), .A(n_74), .B(n_83), .CI(n_86));
  OAI2BB1X1 g3113(.Y(n_94), .A0N(n_80), .A1N(n_88), .B0(n_91));
  ADDFX1 g3114(.CO(n_92), .S(n_93), .A(n_78), .B(n_76), .CI(n_85));
  OR2X1 g3115(.Y(n_91), .A(n_80), .B(n_88));
  ADDFX1 g3116(.CO(n_89), .S(n_90), .A(n_72), .B(n_73), .CI(n_81));
  ADDFX1 g3117(.CO(n_88), .S(n_87), .A(n_71), .B(n_79), .CI(n_77));
  ADDFX1 g3118(.CO(n_85), .S(n_86), .A(n_64), .B(n_54), .CI(n_82));
  ADDFX1 g3119(.CO(n_83), .S(out_0[0]), .A(n_52), .B(n_68), .CI(n_58));
  ADDFX1 g3120(.CO(n_81), .S(n_82), .A(n_70), .B(n_60), .CI(n_67));
  ADDFX1 g3121(.CO(n_80), .S(n_79), .A(n_17), .B(n_61), .CI(n_55));
  ADDFX1 g3122(.CO(n_77), .S(n_78), .A(n_65), .B(n_56), .CI(n_63));
  ADDFX1 g3123(.CO(n_75), .S(n_76), .A(n_62), .B(n_59), .CI(n_53));
  ADDFX1 g3124(.CO(n_73), .S(n_74), .A(n_51), .B(n_66), .CI(n_57));
  ADDFX1 g3125(.CO(n_71), .S(n_72), .A(n_29), .B(n_18), .CI(n_69));
  ADDFX1 g3126(.CO(n_69), .S(n_70), .A(in_34[0]), .B(n_39), .CI(n_31));
  ADDFX1 g3127(.CO(n_67), .S(n_68), .A(n_40), .B(n_36), .CI(n_44));
  ADDFX1 g3128(.CO(n_65), .S(n_66), .A(n_33), .B(n_43), .CI(n_35));
  ADDFX1 g3129(.CO(n_63), .S(n_64), .A(n_14), .B(n_30), .CI(n_20));
  ADDFX1 g3130(.CO(n_61), .S(n_62), .A(n_13), .B(n_37), .CI(n_41));
  ADDFX1 g3131(.CO(n_59), .S(n_60), .A(n_47), .B(n_49), .CI(n_42));
  ADDFX1 g3132(.CO(n_57), .S(n_58), .A(n_48), .B(n_50), .CI(n_32));
  ADDFX1 g3133(.CO(n_55), .S(n_56), .A(n_23), .B(n_27), .CI(n_19));
  ADDFX1 g3134(.CO(n_53), .S(n_54), .A(n_28), .B(n_38), .CI(n_24));
  ADDFX1 g3135(.CO(n_51), .S(n_52), .A(n_7), .B(in_7[0]), .CI(n_34));
  ADDFX1 g3136(.CO(n_49), .S(n_50), .A(in_33[0]), .B(n_4), .CI(n_11));
  INVX1 g3137(.Y(n_48), .A(n_46));
  INVX1 g3138(.Y(n_47), .A(n_45));
  ADDFX1 g3139(.CO(n_45), .S(n_46), .A(in_30[0]), .B(in_39[0]), .CI(in_40[0]));
  ADDFX1 g3140(.CO(n_43), .S(n_44), .A(in_25[0]), .B(n_5), .CI(n_9));
  ADDFX1 g3141(.CO(n_41), .S(n_42), .A(in_0[1]), .B(in_18[1]), .CI(in_35[1]));
  ADDFX1 g3142(.CO(n_39), .S(n_40), .A(in_9[0]), .B(n_1), .CI(in_41[0]));
  ADDFX1 g3143(.CO(n_37), .S(n_38), .A(in_4[1]), .B(n_2), .CI(n_12));
  ADDFX1 g3144(.CO(n_35), .S(n_36), .A(in_6[0]), .B(n_3), .CI(n_10));
  ADDFX1 g3145(.CO(n_33), .S(n_34), .A(in_17), .B(in_5), .CI(in_32));
  ADDFX1 g3146(.CO(n_31), .S(n_32), .A(in_11[0]), .B(n_8), .CI(in_38[0]));
  ADDFX1 g3147(.CO(n_29), .S(n_30), .A(in_3[1]), .B(n_6), .CI(in_7[1]));
  INVX1 g3148(.Y(n_28), .A(n_26));
  INVX1 g3149(.Y(n_27), .A(n_25));
  ADDFX1 g3150(.CO(n_25), .S(n_26), .A(in_2[1]), .B(in_24[1]), .CI(in_29[1]));
  INVX1 g3151(.Y(n_24), .A(n_22));
  INVX1 g3152(.Y(n_23), .A(n_21));
  ADDFX1 g3153(.CO(n_21), .S(n_22), .A(in_14[1]), .B(in_10[1]), .CI(in_28[1]));
  ADDFX1 g3154(.CO(n_19), .S(n_20), .A(in_19[1]), .B(in_16[1]), .CI(in_31[1]));
  INVX1 g3155(.Y(n_18), .A(n_16));
  INVX1 g3156(.Y(n_17), .A(n_15));
  ADDFX1 g3157(.CO(n_15), .S(n_16), .A(in_34[0]), .B(in_25[0]), .CI(in_38[0]));
  OAI21X1 g3158(.Y(n_14), .A0(in_22[1]), .A1(in_36[1]), .B0(n_13));
  NAND2X1 g3159(.Y(n_13), .A(in_36[1]), .B(in_22[1]));
  INVX1 g3160(.Y(n_12), .A(in_26[1]));
  INVX1 g3161(.Y(n_11), .A(in_37[0]));
  INVX1 g3162(.Y(n_10), .A(in_12[0]));
  INVX1 g3163(.Y(n_9), .A(in_1[0]));
  INVX1 g3164(.Y(n_8), .A(in_15[0]));
  INVX1 g3165(.Y(n_7), .A(in_34[0]));
  INVX1 g3166(.Y(n_6), .A(in_13[1]));
  INVX1 g3167(.Y(n_5), .A(in_27[0]));
  INVX1 g3168(.Y(n_4), .A(in_23[0]));
  INVX1 g3169(.Y(n_3), .A(in_8[0]));
  INVX1 g3170(.Y(n_2), .A(in_21[1]));
  INVX1 g3171(.Y(n_1), .A(in_20[0]));
endmodule

module WALLACE_CSA_DUMMY_OP131_group_106210(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , out_0);
input  in_23, in_30, in_35, in_46;
input   [4:0] in_0;
input   [2:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [9:0] in_4;
input   [6:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [2:0] in_12;
input   [4:0] in_13;
input   [1:0] in_14;
input   [1:0] in_15;
input   [2:0] in_16;
input   [4:0] in_17;
input   [3:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [2:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [1:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [1:0] in_34;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
input   [2:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [4:0] in_47;
input   [4:0] in_48;
output  [9:0] out_0;
wire  n_171, n_168, n_166, n_164, n_162, n_161, n_160, n_159, n_158, n_157, 
    n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_148, n_147, n_146, 
    n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, 
    n_135, n_134, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, 
    n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, 
    n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, 
    n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, 
    n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, 
    n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, 
    n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
    n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
    n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, 
    n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
    n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
    n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_46, in_35, in_30, 
    in_23;
wire   [9:0] out_0;
wire   [3:0] in_18;
wire   [1:0] in_45;
wire   [1:0] in_41;
wire   [1:0] in_34;
wire   [1:0] in_33;
wire   [1:0] in_31;
wire   [1:0] in_25;
wire   [1:0] in_21;
wire   [1:0] in_15;
wire   [1:0] in_14;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_5;
wire   [9:0] in_4;
wire   [2:0] in_42;
wire   [2:0] in_24;
wire   [2:0] in_16;
wire   [2:0] in_12;
wire   [2:0] in_1;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_32;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_17;
wire   [4:0] in_13;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  AOI22X1 g5380(.Y(out_0[9]), .A0(n_126), .A1(n_171), .B0(n_22), .B1(n_109));
  XNOR2X1 g5381(.Y(out_0[7]), .A(n_131), .B(n_171));
  ADDFX1 g5382(.CO(n_171), .S(out_0[6]), .A(n_158), .B(n_116), .CI(n_168));
  ADDFX1 g5383(.CO(n_168), .S(out_0[5]), .A(n_160), .B(n_159), .CI(n_166));
  ADDFX1 g5384(.CO(n_166), .S(out_0[4]), .A(n_156), .B(n_161), .CI(n_164));
  ADDFX1 g5385(.CO(n_164), .S(out_0[3]), .A(n_153), .B(n_157), .CI(n_162));
  ADDFX1 g5386(.CO(n_162), .S(out_0[2]), .A(n_137), .B(n_148), .CI(n_151));
  ADDFX1 g5387(.CO(n_160), .S(n_161), .A(n_145), .B(n_152), .CI(n_155));
  ADDFX1 g5388(.CO(n_158), .S(n_159), .A(n_144), .B(n_154), .CI(n_108));
  ADDFX1 g5389(.CO(n_156), .S(n_157), .A(n_136), .B(n_147), .CI(n_150));
  ADDFX1 g5390(.CO(n_154), .S(n_155), .A(n_142), .B(in_4[4]), .CI(n_146));
  ADDFX1 g5391(.CO(n_152), .S(n_153), .A(n_134), .B(n_143), .CI(n_140));
  ADDFX1 g5392(.CO(n_150), .S(n_151), .A(n_135), .B(n_138), .CI(n_141));
  ADDFX1 g5393(.CO(n_148), .S(out_0[1]), .A(n_139), .B(n_132), .CI(n_119));
  ADDFX1 g5394(.CO(n_146), .S(n_147), .A(n_124), .B(n_130), .CI(in_4[3]));
  ADDFX1 g5395(.CO(n_144), .S(n_145), .A(n_106), .B(n_114), .CI(n_129));
  ADDFX1 g5396(.CO(n_142), .S(n_143), .A(n_127), .B(n_115), .CI(n_112));
  ADDFX1 g5397(.CO(n_140), .S(n_141), .A(n_120), .B(n_110), .CI(in_4[2]));
  ADDFX1 g5398(.CO(n_138), .S(n_139), .A(n_121), .B(n_123), .CI(n_111));
  ADDFX1 g5399(.CO(n_136), .S(n_137), .A(n_113), .B(n_125), .CI(n_118));
  ADDFX1 g5400(.CO(n_134), .S(n_135), .A(n_102), .B(n_128), .CI(n_122));
  ADDFX1 g5401(.CO(n_132), .S(out_0[0]), .A(n_79), .B(n_75), .CI(n_105));
  NAND2X1 g5402(.Y(n_131), .A(n_117), .B(n_126));
  ADDFX1 g5403(.CO(n_129), .S(n_130), .A(n_94), .B(n_92), .CI(n_101));
  ADDFX1 g5404(.CO(n_127), .S(n_128), .A(n_96), .B(n_98), .CI(n_82));
  OAI2BB1X1 g5405(.Y(n_126), .A0N(in_4[6]), .A1N(n_109), .B0(in_4[7]));
  ADDFX1 g5406(.CO(n_124), .S(n_125), .A(n_89), .B(n_93), .CI(n_90));
  ADDFX1 g5407(.CO(n_122), .S(n_123), .A(n_86), .B(n_99), .CI(n_74));
  ADDFX1 g5408(.CO(n_120), .S(n_121), .A(n_72), .B(n_97), .CI(n_83));
  ADDFX1 g5409(.CO(n_118), .S(n_119), .A(n_91), .B(n_104), .CI(in_4[1]));
  NAND2X1 g5410(.Y(n_117), .A(n_22), .B(n_109));
  XNOR2X1 g5411(.Y(n_116), .A(n_107), .B(n_26));
  ADDFX1 g5412(.CO(n_114), .S(n_115), .A(n_69), .B(n_76), .CI(n_88));
  ADDFX1 g5413(.CO(n_112), .S(n_113), .A(n_77), .B(n_84), .CI(n_80));
  ADDFX1 g5414(.CO(n_110), .S(n_111), .A(n_78), .B(n_85), .CI(n_81));
  NAND2X1 g5415(.Y(n_109), .A(in_37[0]), .B(n_107));
  XNOR2X1 g5416(.Y(n_108), .A(n_103), .B(in_4[5]));
  OAI21X1 g5417(.Y(n_107), .A0(n_100), .A1(in_4[5]), .B0(in_37[0]));
  OAI2BB1X1 g5418(.Y(n_106), .A0N(n_68), .A1N(n_95), .B0(n_103));
  ADDFX1 g5419(.CO(n_104), .S(n_105), .A(n_73), .B(n_87), .CI(in_4[0]));
  NAND2BX1 g5420(.Y(n_103), .AN(n_100), .B(in_37[0]));
  ADDFX1 g5421(.CO(n_101), .S(n_102), .A(n_57), .B(n_70), .CI(n_50));
  NAND2BX1 g5422(.Y(n_100), .AN(n_95), .B(n_56));
  ADDFX1 g5423(.CO(n_98), .S(n_99), .A(n_41), .B(n_64), .CI(n_53));
  ADDFX1 g5424(.CO(n_96), .S(n_97), .A(n_23), .B(n_60), .CI(n_62));
  ADDFX1 g5425(.CO(n_95), .S(n_94), .A(n_66), .B(n_29), .CI(n_49));
  ADDFX1 g5426(.CO(n_92), .S(n_93), .A(n_67), .B(n_32), .CI(n_37));
  ADDFX1 g5427(.CO(n_90), .S(n_91), .A(n_39), .B(n_38), .CI(n_71));
  ADDFX1 g5428(.CO(n_88), .S(n_89), .A(n_45), .B(n_47), .CI(n_14));
  ADDFX1 g5429(.CO(n_86), .S(n_87), .A(n_63), .B(n_52), .CI(n_54));
  ADDFX1 g5430(.CO(n_84), .S(n_85), .A(n_48), .B(n_59), .CI(n_46));
  ADDFX1 g5431(.CO(n_82), .S(n_83), .A(n_51), .B(n_30), .CI(n_35));
  ADDFX1 g5432(.CO(n_80), .S(n_81), .A(n_44), .B(n_34), .CI(in_5[1]));
  ADDFX1 g5433(.CO(n_78), .S(n_79), .A(n_27), .B(n_61), .CI(n_40));
  ADDFX1 g5434(.CO(n_76), .S(n_77), .A(n_58), .B(n_43), .CI(n_33));
  ADDFX1 g5435(.CO(n_74), .S(n_75), .A(n_36), .B(n_65), .CI(n_31));
  ADDFX1 g5436(.CO(n_72), .S(n_73), .A(in_6[0]), .B(in_7[0]), .CI(n_42));
  ADDFX1 g5437(.CO(n_70), .S(n_71), .A(n_16), .B(n_24), .CI(in_9[1]));
  OAI21X1 g5438(.Y(n_69), .A0(in_37[0]), .A1(n_56), .B0(n_68));
  NAND2X1 g5439(.Y(n_68), .A(in_37[0]), .B(n_56));
  ADDFX1 g5440(.CO(n_66), .S(n_67), .A(in_18[2]), .B(n_1), .CI(in_42[1]));
  ADDFX1 g5441(.CO(n_64), .S(n_65), .A(in_10[0]), .B(n_17), .CI(in_11[0]));
  ADDFX1 g5442(.CO(n_62), .S(n_63), .A(in_15[0]), .B(in_26[0]), .CI(in_38[0]));
  ADDFX1 g5443(.CO(n_60), .S(n_61), .A(in_25[0]), .B(n_5), .CI(n_8));
  ADDFX1 g5444(.CO(n_58), .S(n_59), .A(in_15[0]), .B(n_2), .CI(n_7));
  INVX1 g5445(.Y(n_57), .A(n_55));
  ADDFX1 g5446(.CO(n_56), .S(n_55), .A(in_26[0]), .B(in_38[0]), .CI(in_44[2]));
  ADDFX1 g5447(.CO(n_53), .S(n_54), .A(in_3[0]), .B(in_21[0]), .CI(in_46));
  ADDFX1 g5448(.CO(n_51), .S(n_52), .A(in_43[0]), .B(n_11), .CI(n_4));
  ADDFX1 g5449(.CO(n_49), .S(n_50), .A(n_21), .B(n_12), .CI(n_13));
  ADDFX1 g5450(.CO(n_47), .S(n_48), .A(in_31[1]), .B(n_6), .CI(in_37[0]));
  ADDFX1 g5451(.CO(n_45), .S(n_46), .A(in_34[1]), .B(in_41[1]), .CI(in_45[1]));
  ADDFX1 g5452(.CO(n_43), .S(n_44), .A(in_14[1]), .B(in_16[1]), .CI(n_19));
  ADDFX1 g5453(.CO(n_41), .S(n_42), .A(n_10), .B(n_15), .CI(in_30));
  ADDFX1 g5454(.CO(n_39), .S(n_40), .A(in_9[0]), .B(in_37[0]), .CI(in_8[0]));
  ADDFX1 g5455(.CO(n_37), .S(n_38), .A(in_42[1]), .B(in_8[1]), .CI(n_3));
  ADDFX1 g5456(.CO(n_35), .S(n_36), .A(in_5[0]), .B(in_23), .CI(in_33[0]));
  ADDFX1 g5457(.CO(n_33), .S(n_34), .A(in_12[1]), .B(in_1[1]), .CI(n_18));
  XNOR2X1 g5458(.Y(n_32), .A(in_43[0]), .B(n_25));
  XOR2XL g5459(.Y(n_31), .A(in_27[0]), .B(n_25));
  OAI21X1 g5460(.Y(n_30), .A0(in_27[0]), .A1(n_9), .B0(n_28));
  OAI22X1 g5461(.Y(n_29), .A0(in_48[0]), .A1(n_0), .B0(in_43[0]), .B1(n_9));
  OAI2BB1X1 g5462(.Y(n_28), .A0N(in_27[0]), .A1N(n_9), .B0(in_48[0]));
  OAI2BB1X1 g5463(.Y(n_27), .A0N(in_35), .A1N(n_20), .B0(n_23));
  XNOR2X1 g5464(.Y(n_26), .A(in_37[0]), .B(in_4[6]));
  MX2XL g5465(.Y(n_25), .A(n_9), .B(in_24[0]), .S0(in_48[0]));
  XOR2XL g5466(.Y(n_24), .A(in_36[1]), .B(in_19[1]));
  OR2X1 g5467(.Y(n_23), .A(in_35), .B(n_20));
  NOR2BX1 g5468(.Y(n_22), .AN(in_4[6]), .B(in_4[7]));
  NOR2X1 g5469(.Y(n_21), .A(in_36[1]), .B(in_19[1]));
  INVX1 g5471(.Y(n_20), .A(in_47[0]));
  INVX1 g5472(.Y(n_19), .A(in_22[1]));
  INVX1 g5473(.Y(n_18), .A(in_32[1]));
  INVX1 g5474(.Y(n_17), .A(in_17[0]));
  INVX1 g5475(.Y(n_16), .A(in_7[1]));
  INVX1 g5476(.Y(n_15), .A(in_13[0]));
  INVX1 g5477(.Y(n_14), .A(in_5[2]));
  INVX1 g5478(.Y(n_13), .A(in_8[2]));
  INVX1 g5479(.Y(n_12), .A(in_9[2]));
  INVX1 g5480(.Y(n_11), .A(in_0[0]));
  INVX1 g5481(.Y(n_10), .A(in_29[0]));
  INVX1 g5482(.Y(n_9), .A(in_24[0]));
  INVX1 g5483(.Y(n_8), .A(in_28[0]));
  INVX1 g5484(.Y(n_7), .A(in_40[1]));
  INVX1 g5485(.Y(n_6), .A(in_10[1]));
  INVX1 g5486(.Y(n_5), .A(in_2[0]));
  INVX1 g5487(.Y(n_4), .A(in_39[0]));
  INVX1 g5488(.Y(n_3), .A(in_6[1]));
  INVX1 g5489(.Y(n_2), .A(in_20[1]));
  INVX1 g5491(.Y(n_1), .A(in_3[0]));
  NOR2BX1 g2(.Y(n_0), .AN(in_43[0]), .B(in_24[0]));
endmodule

module WALLACE_CSA_DUMMY_OP140_group_106218(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, out_0);
input  in_67, in_70, in_71, in_76, in_82;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [9:0] in_4;
input   [7:0] in_5;
input   [7:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [2:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [2:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [4:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [4:0] in_56;
input   [2:0] in_57;
input   [3:0] in_58;
input   [1:0] in_59;
input   [4:0] in_60;
input   [1:0] in_61;
input   [4:0] in_62;
input   [1:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [2:0] in_66;
input   [1:0] in_68;
input   [2:0] in_69;
input   [1:0] in_72;
input   [4:0] in_73;
input   [3:0] in_74;
input   [1:0] in_75;
input   [2:0] in_77;
input   [1:0] in_78;
input   [4:0] in_79;
input   [1:0] in_80;
input   [1:0] in_81;
input   [3:0] in_83;
input   [4:0] in_84;
output  [9:0] out_0;
wire  n_294, n_291, n_289, n_287, n_285, n_284, n_283, n_282, n_281, n_279, 
    n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, 
    n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, 
    n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, n_249, n_248, 
    n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, 
    n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, 
    n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_219, n_218, n_217, 
    n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, n_207, 
    n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
    n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, n_187, 
    n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, 
    n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
    n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, 
    n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, 
    n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
    n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, 
    n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_82, in_76, 
    in_71, in_70, in_67;
wire   [9:0] out_0;
wire   [3:0] in_83;
wire   [3:0] in_74;
wire   [3:0] in_58;
wire   [1:0] in_81;
wire   [1:0] in_80;
wire   [1:0] in_78;
wire   [1:0] in_75;
wire   [1:0] in_72;
wire   [1:0] in_68;
wire   [1:0] in_63;
wire   [1:0] in_61;
wire   [1:0] in_59;
wire   [1:0] in_32;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [7:0] in_6;
wire   [7:0] in_5;
wire   [9:0] in_4;
wire   [4:0] in_84;
wire   [4:0] in_79;
wire   [4:0] in_73;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_62;
wire   [4:0] in_60;
wire   [4:0] in_56;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_51;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_77;
wire   [2:0] in_69;
wire   [2:0] in_66;
wire   [2:0] in_57;
wire   [2:0] in_42;
wire   [2:0] in_30;
wire   [2:0] in_22;
wire   [2:0] in_0;
  OA21X1 g8885(.Y(out_0[8]), .A0(n_263), .A1(n_294), .B0(out_0[9]));
  NAND2X1 g8886(.Y(out_0[9]), .A(n_263), .B(n_294));
  ADDFX1 g8887(.CO(n_294), .S(out_0[7]), .A(n_266), .B(n_277), .CI(n_291));
  ADDFX1 g8888(.CO(n_291), .S(out_0[6]), .A(n_281), .B(n_278), .CI(n_289));
  ADDFX1 g8889(.CO(n_289), .S(out_0[5]), .A(n_283), .B(n_282), .CI(n_287));
  ADDFX1 g8890(.CO(n_287), .S(out_0[4]), .A(n_275), .B(n_284), .CI(n_285));
  ADDFX1 g8891(.CO(n_285), .S(out_0[3]), .A(n_269), .B(n_279), .CI(n_276));
  ADDFX1 g8892(.CO(n_283), .S(n_284), .A(n_265), .B(n_271), .CI(n_274));
  ADDFX1 g8893(.CO(n_281), .S(n_282), .A(n_264), .B(n_273), .CI(n_268));
  ADDFX1 g8894(.CO(n_279), .S(out_0[2]), .A(n_270), .B(n_257), .CI(n_250));
  ADDFX1 g8895(.CO(n_277), .S(n_278), .A(n_261), .B(in_4[6]), .CI(n_267));
  ADDFX1 g8896(.CO(n_275), .S(n_276), .A(n_260), .B(n_249), .CI(n_272));
  ADDFX1 g8897(.CO(n_273), .S(n_274), .A(n_245), .B(n_259), .CI(in_4[4]));
  ADDFX1 g8898(.CO(n_271), .S(n_272), .A(n_253), .B(n_246), .CI(in_4[3]));
  ADDFX1 g8899(.CO(n_269), .S(n_270), .A(n_242), .B(n_254), .CI(n_243));
  ADDFX1 g8900(.CO(n_267), .S(n_268), .A(n_252), .B(n_255), .CI(in_4[5]));
  OAI2BB1X1 g8901(.Y(n_266), .A0N(n_262), .A1N(n_36), .B0(n_263));
  ADDFX1 g8902(.CO(n_264), .S(n_265), .A(n_240), .B(n_247), .CI(n_256));
  NAND2BX1 g8903(.Y(n_263), .AN(n_262), .B(in_4[7]));
  ADDFX1 g8904(.CO(n_262), .S(n_261), .A(n_182), .B(n_225), .CI(n_251));
  ADDFX1 g8905(.CO(n_259), .S(n_260), .A(n_241), .B(n_224), .CI(n_248));
  ADDFX1 g8906(.CO(n_257), .S(out_0[1]), .A(n_219), .B(n_238), .CI(n_244));
  ADDFX1 g8907(.CO(n_255), .S(n_256), .A(n_232), .B(n_233), .CI(n_223));
  ADDFX1 g8908(.CO(n_253), .S(n_254), .A(n_222), .B(n_227), .CI(n_236));
  ADDFX1 g8909(.CO(n_251), .S(n_252), .A(n_231), .B(n_226), .CI(n_239));
  ADDFX1 g8910(.CO(n_249), .S(n_250), .A(n_230), .B(n_237), .CI(in_4[2]));
  ADDFX1 g8911(.CO(n_247), .S(n_248), .A(n_215), .B(n_218), .CI(n_235));
  ADDFX1 g8912(.CO(n_245), .S(n_246), .A(n_221), .B(n_234), .CI(n_229));
  ADDFX1 g8913(.CO(n_243), .S(n_244), .A(n_228), .B(n_212), .CI(in_4[1]));
  ADDFX1 g8914(.CO(n_241), .S(n_242), .A(n_216), .B(n_204), .CI(n_211));
  ADDFX1 g8915(.CO(n_239), .S(n_240), .A(n_195), .B(n_198), .CI(n_217));
  ADDFX1 g8916(.CO(n_237), .S(n_238), .A(n_210), .B(n_208), .CI(n_187));
  ADDFX1 g8917(.CO(n_235), .S(n_236), .A(n_139), .B(n_209), .CI(n_186));
  ADDFX1 g8918(.CO(n_233), .S(n_234), .A(n_206), .B(n_196), .CI(n_203));
  ADDFX1 g8919(.CO(n_231), .S(n_232), .A(n_165), .B(n_205), .CI(n_213));
  ADDFX1 g8920(.CO(n_229), .S(n_230), .A(n_200), .B(n_207), .CI(n_183));
  ADDFX1 g8921(.CO(n_227), .S(n_228), .A(n_189), .B(n_192), .CI(n_194));
  ADDFX1 g8922(.CO(n_225), .S(n_226), .A(n_164), .B(n_133), .CI(n_197));
  ADDFX1 g8923(.CO(n_223), .S(n_224), .A(n_214), .B(n_199), .CI(n_185));
  ADDFX1 g8924(.CO(n_221), .S(n_222), .A(n_202), .B(n_191), .CI(n_193));
  ADDFX1 g8925(.CO(n_219), .S(out_0[0]), .A(n_190), .B(n_171), .CI(n_188));
  ADDFX1 g8926(.CO(n_217), .S(n_218), .A(n_141), .B(n_201), .CI(n_172));
  ADDFX1 g8927(.CO(n_215), .S(n_216), .A(n_159), .B(n_176), .CI(n_173));
  ADDFX1 g8928(.CO(n_213), .S(n_214), .A(n_128), .B(n_180), .CI(n_158));
  ADDFX1 g8929(.CO(n_211), .S(n_212), .A(n_177), .B(n_170), .CI(n_184));
  ADDFX1 g8930(.CO(n_209), .S(n_210), .A(n_175), .B(n_163), .CI(n_134));
  ADDFX1 g8931(.CO(n_207), .S(n_208), .A(n_157), .B(n_155), .CI(n_179));
  ADDFX1 g8932(.CO(n_205), .S(n_206), .A(n_87), .B(n_168), .CI(n_166));
  ADDFX1 g8933(.CO(n_203), .S(n_204), .A(n_154), .B(n_169), .CI(n_178));
  ADDFX1 g8934(.CO(n_201), .S(n_202), .A(n_144), .B(n_162), .CI(n_174));
  ADDFX1 g8935(.CO(n_199), .S(n_200), .A(n_181), .B(n_167), .CI(n_156));
  ADDFX1 g8936(.CO(n_197), .S(n_198), .A(n_130), .B(n_160), .CI(n_140));
  ADDFX1 g8937(.CO(n_195), .S(n_196), .A(n_14), .B(n_161), .CI(n_138));
  ADDFX1 g8938(.CO(n_193), .S(n_194), .A(n_151), .B(n_145), .CI(n_148));
  ADDFX1 g8939(.CO(n_191), .S(n_192), .A(n_146), .B(n_137), .CI(n_142));
  ADDFX1 g8940(.CO(n_189), .S(n_190), .A(n_143), .B(n_147), .CI(n_135));
  ADDFX1 g8941(.CO(n_187), .S(n_188), .A(n_153), .B(n_149), .CI(in_4[0]));
  ADDFX1 g8942(.CO(n_185), .S(n_186), .A(n_136), .B(n_150), .CI(in_6[2]));
  ADDFX1 g8943(.CO(n_183), .S(n_184), .A(n_115), .B(n_152), .CI(in_6[1]));
  OAI211X1 g8944(.Y(n_182), .A0(in_49[1]), .A1(n_45), .B0(n_46), .C0(n_132));
  ADDFX1 g8945(.CO(n_180), .S(n_181), .A(in_81[0]), .B(n_90), .CI(n_124));
  ADDFX1 g8946(.CO(n_178), .S(n_179), .A(n_69), .B(n_117), .CI(in_5[1]));
  ADDFX1 g8947(.CO(n_176), .S(n_177), .A(n_105), .B(n_81), .CI(n_78));
  ADDFX1 g8948(.CO(n_174), .S(n_175), .A(n_58), .B(n_50), .CI(n_52));
  ADDFX1 g8949(.CO(n_172), .S(n_173), .A(n_107), .B(n_114), .CI(n_16));
  ADDFX1 g8950(.CO(n_170), .S(n_171), .A(n_119), .B(n_79), .CI(in_6[0]));
  ADDFX1 g8951(.CO(n_168), .S(n_169), .A(n_94), .B(n_122), .CI(n_104));
  ADDFX1 g8952(.CO(n_166), .S(n_167), .A(n_68), .B(n_116), .CI(n_80));
  ADDFX1 g8953(.CO(n_164), .S(n_165), .A(n_47), .B(n_48), .CI(n_129));
  ADDFX1 g8954(.CO(n_162), .S(n_163), .A(n_118), .B(n_66), .CI(n_120));
  ADDFX1 g8955(.CO(n_160), .S(n_161), .A(n_96), .B(n_82), .CI(n_106));
  ADDFX1 g8956(.CO(n_158), .S(n_159), .A(n_108), .B(n_110), .CI(n_63));
  ADDFX1 g8957(.CO(n_156), .S(n_157), .A(n_91), .B(n_109), .CI(n_125));
  ADDFX1 g8958(.CO(n_154), .S(n_155), .A(n_74), .B(n_95), .CI(n_123));
  ADDFX1 g8959(.CO(n_152), .S(n_153), .A(n_121), .B(n_67), .CI(n_73));
  ADDFX1 g8960(.CO(n_150), .S(n_151), .A(in_15[1]), .B(n_76), .CI(n_72));
  ADDFX1 g8961(.CO(n_148), .S(n_149), .A(n_59), .B(n_75), .CI(in_5[0]));
  ADDFX1 g8962(.CO(n_146), .S(n_147), .A(n_93), .B(n_71), .CI(n_99));
  ADDFX1 g8963(.CO(n_144), .S(n_145), .A(n_40), .B(n_70), .CI(n_84));
  ADDFX1 g8964(.CO(n_142), .S(n_143), .A(n_43), .B(n_101), .CI(n_51));
  ADDFX1 g8965(.CO(n_140), .S(n_141), .A(n_102), .B(n_44), .CI(n_62));
  ADDFX1 g8966(.CO(n_138), .S(n_139), .A(n_103), .B(n_97), .CI(n_83));
  ADDFX1 g8967(.CO(n_136), .S(n_137), .A(n_98), .B(n_100), .CI(n_92));
  ADDFX1 g8968(.CO(n_134), .S(n_135), .A(n_53), .B(n_85), .CI(n_77));
  XNOR2X1 g8969(.Y(n_133), .A(n_131), .B(n_126));
  NAND2BXL g8970(.Y(n_132), .AN(n_126), .B(n_131));
  ADDFX1 g8971(.CO(n_131), .S(n_130), .A(in_49[1]), .B(n_38), .CI(n_86));
  OAI2BB1X1 g8972(.Y(n_129), .A0N(in_38[0]), .A1N(in_39[0]), .B0(n_127));
  XNOR2X1 g8973(.Y(n_128), .A(n_42), .B(n_111));
  OAI21X1 g8974(.Y(n_127), .A0(in_38[0]), .A1(in_39[0]), .B0(n_111));
  XNOR2X1 g8975(.Y(n_126), .A(n_45), .B(n_49));
  ADDFX1 g8976(.CO(n_124), .S(n_125), .A(in_31[0]), .B(in_42[1]), .CI(in_69[1]));
  ADDFX1 g8977(.CO(n_122), .S(n_123), .A(in_41[0]), .B(in_68[1]), .CI(in_39[0]));
  ADDFX1 g8978(.CO(n_120), .S(n_121), .A(in_64[0]), .B(in_80[0]), .CI(in_75[0]));
  ADDFX1 g8979(.CO(n_118), .S(n_119), .A(in_25[0]), .B(in_32[0]), .CI(in_72[0]));
  ADDFX1 g8980(.CO(n_116), .S(n_117), .A(n_8), .B(in_57[1]), .CI(n_9));
  INVX1 g8981(.Y(n_115), .A(n_113));
  INVX1 g8982(.Y(n_114), .A(n_112));
  ADDFX1 g8983(.CO(n_112), .S(n_113), .A(in_81[0]), .B(in_14[1]), .CI(in_21[1]));
  ADDFX1 g8984(.CO(n_111), .S(n_110), .A(n_21), .B(n_24), .CI(in_83[2]));
  ADDFX1 g8985(.CO(n_108), .S(n_109), .A(in_66[1]), .B(in_75[0]), .CI(in_78[1]));
  ADDFX1 g8986(.CO(n_106), .S(n_107), .A(n_4), .B(n_6), .CI(in_58[2]));
  ADDFX1 g8987(.CO(n_104), .S(n_105), .A(in_49[1]), .B(n_31), .CI(n_19));
  INVX1 g8988(.Y(n_103), .A(n_89));
  INVX1 g8989(.Y(n_102), .A(n_88));
  INVX1 g8990(.Y(n_101), .A(n_65));
  INVX1 g8991(.Y(n_100), .A(n_64));
  INVX1 g8992(.Y(n_99), .A(n_61));
  INVX1 g8993(.Y(n_98), .A(n_60));
  INVX1 g8994(.Y(n_97), .A(n_57));
  INVX1 g8995(.Y(n_96), .A(n_56));
  INVX1 g8996(.Y(n_95), .A(n_55));
  INVX1 g8997(.Y(n_94), .A(n_54));
  ADDFX1 g8998(.CO(n_92), .S(n_93), .A(in_39[0]), .B(in_76), .CI(in_81[0]));
  ADDFX1 g8999(.CO(n_90), .S(n_91), .A(in_0[1]), .B(n_34), .CI(n_28));
  ADDFX1 g9000(.CO(n_88), .S(n_89), .A(in_34[2]), .B(in_45[0]), .CI(in_51[2]));
  ADDFX1 g9001(.CO(n_86), .S(n_87), .A(in_26[3]), .B(in_49[1]), .CI(in_41[0]));
  ADDFX1 g9002(.CO(n_84), .S(n_85), .A(n_13), .B(n_26), .CI(in_41[0]));
  ADDFX1 g9003(.CO(n_82), .S(n_83), .A(n_25), .B(in_74[2]), .CI(n_20));
  ADDFX1 g9004(.CO(n_80), .S(n_81), .A(in_30[1]), .B(n_30), .CI(n_32));
  ADDFX1 g9005(.CO(n_78), .S(n_79), .A(in_67), .B(in_21[0]), .CI(in_14[0]));
  ADDFX1 g9006(.CO(n_76), .S(n_77), .A(in_31[0]), .B(in_45[0]), .CI(n_35));
  ADDFX1 g9007(.CO(n_74), .S(n_75), .A(in_40[0]), .B(n_11), .CI(in_61[0]));
  ADDFX1 g9008(.CO(n_72), .S(n_73), .A(in_63[0]), .B(in_70), .CI(in_56[0]));
  ADDFX1 g9009(.CO(n_70), .S(n_71), .A(n_10), .B(in_50[0]), .CI(n_5));
  ADDFX1 g9010(.CO(n_68), .S(n_69), .A(in_22[1]), .B(n_29), .CI(n_33));
  ADDFX1 g9011(.CO(n_66), .S(n_67), .A(in_38[0]), .B(n_15), .CI(in_82));
  ADDFX1 g9012(.CO(n_64), .S(n_65), .A(in_3[0]), .B(in_20[0]), .CI(in_84[0]));
  ADDFX1 g9013(.CO(n_62), .S(n_63), .A(in_77[2]), .B(n_23), .CI(n_7));
  ADDFX1 g9014(.CO(n_60), .S(n_61), .A(in_23[0]), .B(in_9[0]), .CI(in_33[0]));
  ADDFX1 g9015(.CO(n_58), .S(n_59), .A(n_27), .B(n_12), .CI(in_59[0]));
  ADDFX1 g9016(.CO(n_56), .S(n_57), .A(in_27[2]), .B(in_24[2]), .CI(in_65[2]));
  ADDFX1 g9017(.CO(n_54), .S(n_55), .A(in_13[1]), .B(in_17[1]), .CI(in_36[1]));
  ADDFX1 g9018(.CO(n_52), .S(n_53), .A(in_15[0]), .B(n_17), .CI(in_60[0]));
  ADDFX1 g9019(.CO(n_50), .S(n_51), .A(in_7[0]), .B(in_71), .CI(n_18));
  XNOR2X1 g9020(.Y(n_49), .A(in_49[1]), .B(n_46));
  MXI2XL g9021(.Y(n_48), .A(n_22), .B(in_26[3]), .S0(n_42));
  XNOR2X1 g9022(.Y(n_47), .A(in_25[0]), .B(n_0));
  AOI22X1 g9023(.Y(n_46), .A0(n_2), .A1(n_41), .B0(n_22), .B1(n_3));
  AOI21X1 g9024(.Y(n_45), .A0(n_1), .A1(n_39), .B0(n_37));
  NAND2X1 g9025(.Y(n_44), .A(n_39), .B(n_38));
  OAI21X1 g9026(.Y(n_43), .A0(in_1[0]), .A1(in_19[0]), .B0(n_40));
  AOI22X1 g9028(.Y(n_42), .A0(in_38[0]), .A1(n_2), .B0(n_3), .B1(in_39[0]));
  NAND2XL g9029(.Y(n_41), .A(in_26[3]), .B(in_38[0]));
  NAND2X1 g9030(.Y(n_40), .A(in_19[0]), .B(in_1[0]));
  NAND2X1 g9031(.Y(n_39), .A(in_25[0]), .B(in_31[0]));
  INVX1 g9032(.Y(n_38), .A(n_37));
  NOR2X1 g9033(.Y(n_37), .A(in_25[0]), .B(in_31[0]));
  INVX1 g9034(.Y(n_36), .A(in_4[7]));
  INVX1 g9035(.Y(n_35), .A(in_62[0]));
  INVX1 g9036(.Y(n_34), .A(in_73[1]));
  INVX1 g9037(.Y(n_33), .A(in_53[1]));
  INVX1 g9038(.Y(n_32), .A(in_47[1]));
  INVX1 g9039(.Y(n_31), .A(in_8[1]));
  INVX1 g9040(.Y(n_30), .A(in_29[1]));
  INVX1 g9041(.Y(n_29), .A(in_48[1]));
  INVX1 g9042(.Y(n_28), .A(in_18[1]));
  INVX1 g9043(.Y(n_27), .A(in_11[0]));
  INVX1 g9044(.Y(n_26), .A(in_10[0]));
  INVX1 g9045(.Y(n_25), .A(in_46[2]));
  INVX1 g9046(.Y(n_24), .A(in_60[0]));
  INVX1 g9047(.Y(n_23), .A(in_64[0]));
  INVX1 g9048(.Y(n_22), .A(in_26[3]));
  INVX1 g9049(.Y(n_21), .A(in_56[0]));
  INVX1 g9050(.Y(n_20), .A(in_40[0]));
  INVX1 g9051(.Y(n_19), .A(in_52[1]));
  INVX1 g9052(.Y(n_18), .A(in_79[0]));
  INVX1 g9053(.Y(n_17), .A(in_28[0]));
  INVX1 g9054(.Y(n_16), .A(in_5[2]));
  INVX1 g9055(.Y(n_15), .A(in_12[0]));
  INVX1 g9056(.Y(n_14), .A(in_6[3]));
  INVX1 g9057(.Y(n_13), .A(in_16[0]));
  INVX1 g9058(.Y(n_12), .A(in_43[0]));
  INVX1 g9059(.Y(n_11), .A(in_2[0]));
  INVX1 g9060(.Y(n_10), .A(in_37[0]));
  INVX1 g9061(.Y(n_9), .A(in_35[1]));
  INVX1 g9062(.Y(n_8), .A(in_55[1]));
  INVX1 g9063(.Y(n_7), .A(in_15[2]));
  INVX1 g9064(.Y(n_6), .A(in_54[2]));
  INVX1 g9065(.Y(n_5), .A(in_44[0]));
  INVX1 g9066(.Y(n_4), .A(in_50[0]));
  INVX1 g9067(.Y(n_3), .A(in_38[0]));
  INVX1 g9069(.Y(n_2), .A(in_39[0]));
  INVX1 g9070(.Y(n_1), .A(in_41[0]));
  MXI2XL g2(.Y(n_0), .A(n_1), .B(in_41[0]), .S0(in_31[0]));
endmodule

module WALLACE_CSA_DUMMY_OP144_group_106215(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, out_0);
input  in_36, in_38, in_51, in_52, in_53, in_54, in_72, in_73, in_74;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [9:0] in_4;
input   [8:0] in_5;
input   [7:0] in_6;
input   [6:0] in_7;
input   [4:0] in_8;
input   [4:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [3:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [1:0] in_33;
input   [4:0] in_34;
input   [1:0] in_35;
input   [1:0] in_37;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [2:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [4:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [1:0] in_58;
input   [3:0] in_59;
input   [1:0] in_60;
input   [1:0] in_61;
input   [4:0] in_62;
input   [4:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [3:0] in_66;
input   [4:0] in_67;
input   [1:0] in_68;
input   [1:0] in_69;
input   [4:0] in_70;
input   [2:0] in_71;
input   [1:0] in_75;
output  [9:0] out_0;
wire  n_244, n_242, n_240, n_238, n_236, n_235, n_234, n_233, n_232, n_231, 
    n_230, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, 
    n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_210, n_209, 
    n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, 
    n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, 
    n_188, n_187, n_186, n_185, n_184, n_182, n_181, n_180, n_179, n_178, 
    n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, 
    n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_74, 
    in_73, in_72, in_54, in_53, in_52, in_51, in_38, in_36;
wire   [9:0] out_0;
wire   [1:0] in_75;
wire   [1:0] in_69;
wire   [1:0] in_68;
wire   [1:0] in_61;
wire   [1:0] in_60;
wire   [1:0] in_58;
wire   [1:0] in_37;
wire   [1:0] in_35;
wire   [1:0] in_33;
wire   [3:0] in_66;
wire   [3:0] in_59;
wire   [3:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [6:0] in_7;
wire   [7:0] in_6;
wire   [8:0] in_5;
wire   [9:0] in_4;
wire   [4:0] in_70;
wire   [4:0] in_67;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_63;
wire   [4:0] in_62;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_55;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_34;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_9;
wire   [4:0] in_8;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_71;
wire   [2:0] in_44;
wire   [2:0] in_32;
wire   [2:0] in_3;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g3079(.Y(out_0[9]), .A(n_244));
  ADDFX1 g3080(.CO(n_244), .S(out_0[7]), .A(n_29), .B(n_230), .CI(n_242));
  ADDFX1 g3081(.CO(n_242), .S(out_0[6]), .A(n_234), .B(n_231), .CI(n_240));
  ADDFX1 g3082(.CO(n_240), .S(out_0[5]), .A(n_232), .B(n_235), .CI(n_238));
  ADDFX1 g3083(.CO(n_238), .S(out_0[4]), .A(n_226), .B(n_233), .CI(n_236));
  ADDFX1 g3084(.CO(n_236), .S(out_0[3]), .A(n_216), .B(n_228), .CI(n_227));
  ADDFX1 g3085(.CO(n_234), .S(n_235), .A(n_220), .B(n_224), .CI(n_223));
  ADDFX1 g3086(.CO(n_232), .S(n_233), .A(n_221), .B(n_218), .CI(n_225));
  ADDFX1 g3087(.CO(n_230), .S(n_231), .A(n_202), .B(in_4[6]), .CI(n_222));
  ADDFX1 g3088(.CO(n_228), .S(out_0[2]), .A(n_217), .B(n_205), .CI(n_210));
  ADDFX1 g3089(.CO(n_226), .S(n_227), .A(n_209), .B(n_204), .CI(n_219));
  ADDFX1 g3090(.CO(n_224), .S(n_225), .A(n_212), .B(n_208), .CI(in_4[4]));
  ADDFX1 g3091(.CO(n_222), .S(n_223), .A(n_214), .B(n_203), .CI(in_4[5]));
  ADDFX1 g3092(.CO(n_220), .S(n_221), .A(n_186), .B(n_193), .CI(n_215));
  ADDFX1 g3093(.CO(n_218), .S(n_219), .A(n_206), .B(n_213), .CI(in_4[3]));
  ADDFX1 g3094(.CO(n_216), .S(n_217), .A(n_178), .B(n_207), .CI(n_198));
  ADDFX1 g3095(.CO(n_214), .S(n_215), .A(n_139), .B(n_200), .CI(n_194));
  ADDFX1 g3096(.CO(n_212), .S(n_213), .A(n_201), .B(n_184), .CI(n_196));
  ADDFX1 g3097(.CO(n_210), .S(out_0[1]), .A(n_179), .B(n_182), .CI(n_199));
  ADDFX1 g3098(.CO(n_208), .S(n_209), .A(n_190), .B(n_187), .CI(n_195));
  ADDFX1 g3099(.CO(n_206), .S(n_207), .A(n_154), .B(n_188), .CI(n_197));
  ADDFX1 g3100(.CO(n_204), .S(n_205), .A(n_185), .B(n_191), .CI(in_4[2]));
  ADDFX1 g3101(.CO(n_202), .S(n_203), .A(n_0), .B(n_138), .CI(n_192));
  ADDFX1 g3102(.CO(n_200), .S(n_201), .A(n_164), .B(n_180), .CI(n_157));
  ADDFX1 g3103(.CO(n_198), .S(n_199), .A(n_149), .B(n_189), .CI(in_4[1]));
  ADDFX1 g3104(.CO(n_196), .S(n_197), .A(n_144), .B(n_172), .CI(n_181));
  ADDFX1 g3105(.CO(n_194), .S(n_195), .A(n_140), .B(n_170), .CI(n_177));
  ADDFX1 g3106(.CO(n_192), .S(n_193), .A(n_156), .B(n_176), .CI(n_142));
  ADDFX1 g3107(.CO(n_190), .S(n_191), .A(n_175), .B(n_141), .CI(n_171));
  ADDFX1 g3108(.CO(n_188), .S(n_189), .A(n_145), .B(n_168), .CI(n_173));
  ADDFX1 g3109(.CO(n_186), .S(n_187), .A(n_166), .B(n_174), .CI(n_143));
  ADDFX1 g3110(.CO(n_184), .S(n_185), .A(n_167), .B(n_148), .CI(n_162));
  ADDFX1 g3111(.CO(n_182), .S(out_0[0]), .A(n_153), .B(n_169), .CI(in_4[0]));
  ADDFX1 g3112(.CO(n_180), .S(n_181), .A(n_116), .B(n_108), .CI(n_160));
  ADDFX1 g3113(.CO(n_178), .S(n_179), .A(n_155), .B(n_152), .CI(n_163));
  ADDFX1 g3114(.CO(n_176), .S(n_177), .A(n_128), .B(n_150), .CI(n_158));
  ADDFX1 g3115(.CO(n_174), .S(n_175), .A(n_113), .B(n_110), .CI(n_165));
  ADDFX1 g3116(.CO(n_172), .S(n_173), .A(n_115), .B(n_137), .CI(n_161));
  ADDFX1 g3117(.CO(n_170), .S(n_171), .A(n_123), .B(n_126), .CI(n_159));
  ADDFX1 g3118(.CO(n_168), .S(n_169), .A(n_57), .B(n_107), .CI(n_147));
  ADDFX1 g3119(.CO(n_166), .S(n_167), .A(n_114), .B(n_129), .CI(n_136));
  ADDFX1 g3120(.CO(n_164), .S(n_165), .A(n_77), .B(n_40), .CI(n_151));
  ADDFX1 g3121(.CO(n_162), .S(n_163), .A(n_104), .B(n_146), .CI(in_5[1]));
  ADDFX1 g3122(.CO(n_160), .S(n_161), .A(n_64), .B(n_50), .CI(n_135));
  ADDFX1 g3123(.CO(n_158), .S(n_159), .A(n_44), .B(n_86), .CI(n_133));
  ADDFX1 g3124(.CO(n_156), .S(n_157), .A(n_78), .B(n_122), .CI(n_132));
  ADDFX1 g3125(.CO(n_154), .S(n_155), .A(n_127), .B(n_119), .CI(n_111));
  ADDFX1 g3126(.CO(n_152), .S(n_153), .A(n_131), .B(n_105), .CI(n_101));
  ADDFX1 g3127(.CO(n_150), .S(n_151), .A(n_14), .B(n_21), .CI(n_134));
  ADDFX1 g3128(.CO(n_148), .S(n_149), .A(n_117), .B(n_100), .CI(n_103));
  ADDFX1 g3129(.CO(n_146), .S(n_147), .A(n_83), .B(in_6[0]), .CI(n_121));
  ADDFX1 g3130(.CO(n_144), .S(n_145), .A(n_109), .B(n_130), .CI(n_106));
  ADDFX1 g3131(.CO(n_142), .S(n_143), .A(n_112), .B(n_125), .CI(in_5[3]));
  ADDFX1 g3132(.CO(n_140), .S(n_141), .A(n_118), .B(n_102), .CI(in_5[2]));
  ADDFX1 g3133(.CO(n_138), .S(n_139), .A(n_34), .B(n_124), .CI(n_4));
  ADDFX1 g3134(.CO(n_136), .S(n_137), .A(n_38), .B(n_43), .CI(n_120));
  ADDFX1 g3135(.CO(n_134), .S(n_135), .A(in_60[1]), .B(n_96), .CI(n_99));
  ADDFX1 g3136(.CO(n_132), .S(n_133), .A(n_15), .B(n_98), .CI(n_35));
  ADDFX1 g3137(.CO(n_130), .S(n_131), .A(n_93), .B(n_51), .CI(n_47));
  ADDFX1 g3138(.CO(n_128), .S(n_129), .A(n_94), .B(n_42), .CI(n_90));
  ADDFX1 g3139(.CO(n_126), .S(n_127), .A(n_37), .B(n_87), .CI(n_91));
  ADDFX1 g3140(.CO(n_124), .S(n_125), .A(n_76), .B(n_84), .CI(n_34));
  ADDFX1 g3141(.CO(n_122), .S(n_123), .A(n_58), .B(n_54), .CI(n_36));
  ADDFX1 g3142(.CO(n_120), .S(n_121), .A(in_72), .B(n_97), .CI(n_75));
  ADDFX1 g3143(.CO(n_118), .S(n_119), .A(n_55), .B(n_95), .CI(n_67));
  ADDFX1 g3144(.CO(n_116), .S(n_117), .A(n_46), .B(n_52), .CI(n_88));
  ADDFX1 g3145(.CO(n_114), .S(n_115), .A(in_21[1]), .B(n_92), .CI(n_82));
  ADDFX1 g3146(.CO(n_112), .S(n_113), .A(n_85), .B(n_66), .CI(n_79));
  ADDFX1 g3147(.CO(n_110), .S(n_111), .A(n_70), .B(n_56), .CI(n_41));
  ADDFX1 g3148(.CO(n_108), .S(n_109), .A(n_60), .B(n_62), .CI(n_48));
  ADDFX1 g3149(.CO(n_106), .S(n_107), .A(n_39), .B(n_89), .CI(n_49));
  ADDFX1 g3150(.CO(n_104), .S(n_105), .A(n_63), .B(n_61), .CI(n_65));
  ADDFX1 g3151(.CO(n_102), .S(n_103), .A(n_59), .B(n_45), .CI(in_6[1]));
  ADDFX1 g3152(.CO(n_100), .S(n_101), .A(n_71), .B(n_53), .CI(in_5[0]));
  ADDFX1 g3153(.CO(n_98), .S(n_99), .A(n_30), .B(n_33), .CI(n_74));
  INVX1 g3155(.Y(n_97), .A(n_81));
  INVX1 g3156(.Y(n_96), .A(n_80));
  ADDFX1 g3157(.CO(n_94), .S(n_95), .A(n_6), .B(n_5), .CI(in_75[0]));
  ADDFX1 g3158(.CO(n_92), .S(n_93), .A(in_19[0]), .B(in_53), .CI(in_58[0]));
  ADDFX1 g3159(.CO(n_90), .S(n_91), .A(in_32[1]), .B(n_1), .CI(in_69[0]));
  ADDFX1 g3160(.CO(n_88), .S(n_89), .A(in_54), .B(in_63[0]), .CI(in_75[0]));
  ADDFX1 g3161(.CO(n_86), .S(n_87), .A(in_37[0]), .B(n_2), .CI(n_10));
  ADDFX1 g3162(.CO(n_84), .S(n_85), .A(in_16[2]), .B(n_16), .CI(in_66[2]));
  ADDFX1 g3163(.CO(n_82), .S(n_83), .A(in_36), .B(in_21[0]), .CI(in_44[0]));
  ADDFX1 g3164(.CO(n_80), .S(n_81), .A(in_18[0]), .B(in_23[0]), .CI(n_32));
  ADDFX1 g3165(.CO(n_78), .S(n_79), .A(in_29[0]), .B(n_17), .CI(in_59[2]));
  INVX1 g3166(.Y(n_77), .A(n_73));
  INVX1 g3167(.Y(n_76), .A(n_72));
  INVX1 g3168(.Y(n_75), .A(n_69));
  INVX1 g3169(.Y(n_74), .A(n_68));
  ADDFX1 g3170(.CO(n_72), .S(n_73), .A(in_8[0]), .B(in_48[0]), .CI(in_70[0]));
  ADDFX1 g3171(.CO(n_70), .S(n_71), .A(in_37[0]), .B(in_38), .CI(in_22[0]));
  ADDFX1 g3172(.CO(n_68), .S(n_69), .A(in_12[0]), .B(in_10[0]), .CI(in_14[0]));
  ADDFX1 g3173(.CO(n_66), .S(n_67), .A(in_71[1]), .B(n_23), .CI(n_18));
  ADDFX1 g3174(.CO(n_64), .S(n_65), .A(in_51), .B(in_73), .CI(n_8));
  ADDFX1 g3175(.CO(n_62), .S(n_63), .A(in_41[0]), .B(n_26), .CI(n_28));
  ADDFX1 g3176(.CO(n_60), .S(n_61), .A(in_35[0]), .B(in_25[0]), .CI(in_65[0]));
  ADDFX1 g3177(.CO(n_58), .S(n_59), .A(in_3[1]), .B(in_35[0]), .CI(n_11));
  ADDFX1 g3178(.CO(n_56), .S(n_57), .A(in_15[0]), .B(in_17[0]), .CI(in_20[0]));
  ADDFX1 g3179(.CO(n_54), .S(n_55), .A(in_27[1]), .B(n_25), .CI(n_13));
  ADDFX1 g3180(.CO(n_52), .S(n_53), .A(n_3), .B(n_7), .CI(in_52));
  ADDFX1 g3181(.CO(n_50), .S(n_51), .A(in_48[0]), .B(in_29[0]), .CI(in_74));
  ADDFX1 g3182(.CO(n_48), .S(n_49), .A(in_13[0]), .B(in_26[0]), .CI(in_70[0]));
  ADDFX1 g3183(.CO(n_46), .S(n_47), .A(in_33[0]), .B(n_24), .CI(in_69[0]));
  ADDFX1 g3184(.CO(n_44), .S(n_45), .A(in_61[1]), .B(n_20), .CI(n_9));
  ADDFX1 g3185(.CO(n_42), .S(n_43), .A(in_0[1]), .B(in_44[0]), .CI(n_12));
  ADDFX1 g3186(.CO(n_40), .S(n_41), .A(in_20[1]), .B(n_22), .CI(in_17[1]));
  ADDFX1 g3187(.CO(n_38), .S(n_39), .A(in_28[0]), .B(in_8[0]), .CI(n_27));
  ADDFX1 g3188(.CO(n_36), .S(n_37), .A(in_19[0]), .B(n_19), .CI(in_68[1]));
  OAI21X1 g3189(.Y(n_35), .A0(n_31), .A1(in_6[2]), .B0(n_0));
  INVX1 g3190(.Y(n_34), .A(n_0));
  NAND2X1 g3191(.Y(n_0), .A(n_31), .B(in_6[2]));
  XOR2XL g3192(.Y(n_33), .A(in_26[1]), .B(in_11[1]));
  XNOR2X1 g3193(.Y(n_32), .A(in_24[0]), .B(in_7[0]));
  OR2X1 g3194(.Y(n_31), .A(in_26[1]), .B(in_11[1]));
  NOR2X1 g3195(.Y(n_30), .A(in_24[0]), .B(in_7[0]));
  INVX1 g3196(.Y(n_29), .A(in_4[7]));
  INVX1 g3197(.Y(n_28), .A(in_64[0]));
  INVX1 g3198(.Y(n_27), .A(in_56[0]));
  INVX1 g3199(.Y(n_26), .A(in_30[0]));
  INVX1 g3200(.Y(n_25), .A(in_9[1]));
  INVX1 g3201(.Y(n_24), .A(in_2[0]));
  INVX1 g3202(.Y(n_23), .A(in_46[1]));
  INVX1 g3203(.Y(n_22), .A(in_15[1]));
  INVX1 g3204(.Y(n_21), .A(in_21[2]));
  INVX1 g3205(.Y(n_20), .A(in_40[1]));
  INVX1 g3206(.Y(n_19), .A(in_34[1]));
  INVX1 g3207(.Y(n_18), .A(in_22[1]));
  INVX1 g3208(.Y(n_17), .A(in_50[2]));
  INVX1 g3209(.Y(n_16), .A(in_65[0]));
  INVX1 g3210(.Y(n_15), .A(in_63[0]));
  INVX1 g3211(.Y(n_14), .A(in_41[0]));
  INVX1 g3212(.Y(n_13), .A(in_39[1]));
  INVX1 g3213(.Y(n_12), .A(in_62[1]));
  INVX1 g3214(.Y(n_11), .A(in_43[1]));
  INVX1 g3215(.Y(n_10), .A(in_45[1]));
  INVX1 g3216(.Y(n_9), .A(in_67[1]));
  INVX1 g3217(.Y(n_8), .A(in_42[0]));
  INVX1 g3218(.Y(n_7), .A(in_1[0]));
  INVX1 g3219(.Y(n_6), .A(in_49[1]));
  INVX1 g3220(.Y(n_5), .A(in_57[1]));
  INVX1 g3221(.Y(n_4), .A(in_5[4]));
  INVX1 g3222(.Y(n_3), .A(in_47[0]));
  INVX1 g3223(.Y(n_2), .A(in_31[1]));
  INVX1 g3224(.Y(n_1), .A(in_55[1]));
endmodule

module WALLACE_CSA_DUMMY_OP146_group_106214(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, out_0);
input  in_34, in_35, in_37, in_47, in_68;
input   [4:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [7:0] in_3;
input   [6:0] in_4;
input   [6:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [4:0] in_10;
input   [4:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [1:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [1:0] in_36;
input   [1:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [1:0] in_44;
input   [4:0] in_45;
input   [1:0] in_46;
input   [2:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [1:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [1:0] in_54;
input   [4:0] in_55;
input   [1:0] in_56;
input   [1:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [2:0] in_60;
input   [4:0] in_61;
input   [1:0] in_62;
input   [4:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [1:0] in_67;
input   [1:0] in_69;
input   [4:0] in_70;
input   [1:0] in_71;
input   [4:0] in_72;
input   [4:0] in_73;
input   [4:0] in_74;
input   [1:0] in_75;
output  [9:0] out_0;
wire  n_242, n_240, n_238, n_236, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_224, n_223, n_222, n_221, n_220, n_219, n_218, 
    n_217, n_216, n_215, n_214, n_213, n_212, n_210, n_209, n_208, n_207, 
    n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
    n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, n_187, 
    n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_177, n_176, 
    n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, 
    n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156, 
    n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, 
    n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, 
    n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, 
    n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, 
    n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, 
    n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, 
    n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, 
    n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, 
    n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, 
    n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, 
    n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, 
    n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, 
    n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_68, in_47, 
    in_37, in_35, in_34;
wire   [9:0] out_0;
wire   [2:0] in_60;
wire   [2:0] in_48;
wire   [1:0] in_75;
wire   [1:0] in_71;
wire   [1:0] in_69;
wire   [1:0] in_67;
wire   [1:0] in_62;
wire   [1:0] in_57;
wire   [1:0] in_56;
wire   [1:0] in_54;
wire   [1:0] in_51;
wire   [1:0] in_46;
wire   [1:0] in_44;
wire   [1:0] in_38;
wire   [1:0] in_36;
wire   [1:0] in_14;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_5;
wire   [6:0] in_4;
wire   [7:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_74;
wire   [4:0] in_73;
wire   [4:0] in_72;
wire   [4:0] in_70;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_63;
wire   [4:0] in_61;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_55;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_45;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_11;
wire   [4:0] in_10;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g7683(.Y(out_0[9]), .A(n_242));
  ADDFX1 g7684(.CO(n_242), .S(out_0[7]), .A(n_11), .B(n_228), .CI(n_240));
  ADDFX1 g7685(.CO(n_240), .S(out_0[6]), .A(n_232), .B(n_229), .CI(n_238));
  ADDFX1 g7686(.CO(n_238), .S(out_0[5]), .A(n_233), .B(n_230), .CI(n_236));
  ADDFX1 g7687(.CO(n_236), .S(out_0[4]), .A(n_226), .B(n_231), .CI(n_234));
  ADDFX1 g7688(.CO(n_234), .S(out_0[3]), .A(n_212), .B(n_224), .CI(n_227));
  ADDFX1 g7689(.CO(n_232), .S(n_233), .A(n_221), .B(in_2[5]), .CI(n_222));
  ADDFX1 g7690(.CO(n_230), .S(n_231), .A(n_219), .B(n_216), .CI(n_223));
  ADDFX1 g7691(.CO(n_228), .S(n_229), .A(n_176), .B(n_220), .CI(in_2[6]));
  ADDFX1 g7692(.CO(n_226), .S(n_227), .A(n_215), .B(n_206), .CI(n_217));
  ADDFX1 g7693(.CO(n_224), .S(out_0[2]), .A(n_213), .B(n_210), .CI(n_207));
  ADDFX1 g7694(.CO(n_222), .S(n_223), .A(n_208), .B(n_214), .CI(in_2[4]));
  ADDFX1 g7695(.CO(n_220), .S(n_221), .A(n_181), .B(n_200), .CI(n_218));
  ADDFX1 g7696(.CO(n_218), .S(n_219), .A(n_184), .B(n_196), .CI(n_201));
  ADDFX1 g7697(.CO(n_216), .S(n_217), .A(n_198), .B(n_204), .CI(in_2[3]));
  ADDFX1 g7698(.CO(n_214), .S(n_215), .A(n_197), .B(n_190), .CI(n_209));
  ADDFX1 g7699(.CO(n_212), .S(n_213), .A(n_199), .B(n_205), .CI(n_202));
  ADDFX1 g7700(.CO(n_210), .S(out_0[1]), .A(n_177), .B(n_203), .CI(n_189));
  ADDFX1 g7701(.CO(n_208), .S(n_209), .A(n_185), .B(n_194), .CI(n_193));
  ADDFX1 g7702(.CO(n_206), .S(n_207), .A(n_191), .B(n_188), .CI(in_2[2]));
  ADDFX1 g7703(.CO(n_204), .S(n_205), .A(n_186), .B(n_179), .CI(n_195));
  ADDFX1 g7704(.CO(n_202), .S(n_203), .A(n_180), .B(n_187), .CI(n_148));
  ADDFX1 g7705(.CO(n_200), .S(n_201), .A(n_160), .B(n_174), .CI(n_192));
  ADDFX1 g7706(.CO(n_198), .S(n_199), .A(n_147), .B(n_183), .CI(n_150));
  ADDFX1 g7707(.CO(n_196), .S(n_197), .A(n_182), .B(n_146), .CI(n_164));
  ADDFX1 g7708(.CO(n_194), .S(n_195), .A(n_171), .B(n_172), .CI(n_159));
  ADDFX1 g7709(.CO(n_192), .S(n_193), .A(n_126), .B(n_158), .CI(n_167));
  ADDFX1 g7710(.CO(n_190), .S(n_191), .A(n_169), .B(n_152), .CI(n_165));
  ADDFX1 g7711(.CO(n_188), .S(n_189), .A(n_153), .B(n_151), .CI(in_2[1]));
  ADDFX1 g7712(.CO(n_186), .S(n_187), .A(n_157), .B(n_163), .CI(n_154));
  ADDFX1 g7713(.CO(n_184), .S(n_185), .A(n_170), .B(n_168), .CI(n_161));
  ADDFX1 g7714(.CO(n_182), .S(n_183), .A(n_127), .B(n_162), .CI(n_156));
  XNOR2X1 g7715(.Y(n_181), .A(in_3[4]), .B(n_175));
  ADDFX1 g7716(.CO(n_179), .S(n_180), .A(n_144), .B(n_115), .CI(n_173));
  ADDFX1 g7717(.CO(n_177), .S(out_0[0]), .A(n_145), .B(n_155), .CI(n_149));
  NOR2BX1 g7718(.Y(n_176), .AN(n_175), .B(in_3[4]));
  ADDFX1 g7719(.CO(n_175), .S(n_174), .A(n_140), .B(in_3[4]), .CI(n_166));
  ADDFX1 g7720(.CO(n_172), .S(n_173), .A(n_143), .B(n_134), .CI(n_124));
  ADDFX1 g7721(.CO(n_170), .S(n_171), .A(n_132), .B(n_142), .CI(n_131));
  ADDFX1 g7722(.CO(n_168), .S(n_169), .A(n_128), .B(n_119), .CI(n_106));
  ADDFX1 g7723(.CO(n_166), .S(n_167), .A(n_118), .B(n_130), .CI(in_3[3]));
  ADDFX1 g7724(.CO(n_164), .S(n_165), .A(n_114), .B(n_104), .CI(n_122));
  ADDFX1 g7725(.CO(n_162), .S(n_163), .A(n_109), .B(n_129), .CI(n_116));
  ADDFX1 g7726(.CO(n_160), .S(n_161), .A(n_141), .B(n_112), .CI(n_136));
  ADDFX1 g7727(.CO(n_158), .S(n_159), .A(n_108), .B(n_120), .CI(in_3[2]));
  ADDFX1 g7728(.CO(n_156), .S(n_157), .A(n_121), .B(n_133), .CI(n_138));
  ADDFX1 g7729(.CO(n_154), .S(n_155), .A(n_125), .B(n_117), .CI(n_139));
  ADDFX1 g7730(.CO(n_152), .S(n_153), .A(n_103), .B(n_107), .CI(n_100));
  ADDFX1 g7731(.CO(n_150), .S(n_151), .A(n_110), .B(n_105), .CI(n_123));
  ADDFX1 g7732(.CO(n_148), .S(n_149), .A(n_111), .B(n_101), .CI(in_2[0]));
  ADDFX1 g7733(.CO(n_146), .S(n_147), .A(n_102), .B(n_113), .CI(n_137));
  ADDFX1 g7734(.CO(n_144), .S(n_145), .A(n_49), .B(n_71), .CI(n_135));
  ADDFX1 g7735(.CO(n_142), .S(n_143), .A(n_44), .B(n_98), .CI(n_46));
  ADDFX1 g7736(.CO(n_140), .S(n_141), .A(n_26), .B(n_96), .CI(n_78));
  ADDFX1 g7737(.CO(n_138), .S(n_139), .A(n_41), .B(n_47), .CI(n_93));
  ADDFX1 g7738(.CO(n_136), .S(n_137), .A(n_34), .B(n_76), .CI(n_15));
  ADDFX1 g7739(.CO(n_134), .S(n_135), .A(n_85), .B(n_83), .CI(n_45));
  ADDFX1 g7740(.CO(n_132), .S(n_133), .A(n_66), .B(n_82), .CI(n_84));
  ADDFX1 g7741(.CO(n_130), .S(n_131), .A(n_74), .B(n_50), .CI(n_68));
  ADDFX1 g7742(.CO(n_128), .S(n_129), .A(n_60), .B(n_92), .CI(n_69));
  ADDFX1 g7743(.CO(n_126), .S(n_127), .A(n_97), .B(n_58), .CI(n_79));
  ADDFX1 g7744(.CO(n_124), .S(n_125), .A(in_7[0]), .B(n_67), .CI(n_99));
  ADDFX1 g7745(.CO(n_122), .S(n_123), .A(n_77), .B(n_70), .CI(in_3[1]));
  ADDFX1 g7746(.CO(n_120), .S(n_121), .A(n_30), .B(n_86), .CI(n_52));
  ADDFX1 g7747(.CO(n_118), .S(n_119), .A(n_36), .B(n_90), .CI(n_42));
  ADDFX1 g7748(.CO(n_116), .S(n_117), .A(n_29), .B(n_53), .CI(n_87));
  ADDFX1 g7749(.CO(n_114), .S(n_115), .A(n_37), .B(n_32), .CI(n_81));
  ADDFX1 g7750(.CO(n_112), .S(n_113), .A(n_27), .B(n_56), .CI(n_80));
  ADDFX1 g7751(.CO(n_110), .S(n_111), .A(n_61), .B(n_65), .CI(n_33));
  ADDFX1 g7752(.CO(n_108), .S(n_109), .A(n_64), .B(n_40), .CI(n_28));
  ADDFX1 g7753(.CO(n_106), .S(n_107), .A(n_35), .B(n_51), .CI(in_4[1]));
  ADDFX1 g7754(.CO(n_104), .S(n_105), .A(n_57), .B(n_48), .CI(n_59));
  ADDFX1 g7755(.CO(n_102), .S(n_103), .A(n_43), .B(n_91), .CI(n_75));
  ADDFX1 g7756(.CO(n_100), .S(n_101), .A(n_31), .B(in_4[0]), .CI(in_3[0]));
  ADDFX1 g7757(.CO(n_98), .S(n_99), .A(in_15[0]), .B(n_24), .CI(in_39[0]));
  INVX1 g7758(.Y(n_97), .A(n_95));
  INVX1 g7759(.Y(n_96), .A(n_94));
  ADDFX1 g7760(.CO(n_94), .S(n_95), .A(in_9[0]), .B(in_39[0]), .CI(in_73[0]));
  ADDFX1 g7761(.CO(n_92), .S(n_93), .A(in_35), .B(n_22), .CI(n_2));
  INVX1 g7762(.Y(n_91), .A(n_89));
  INVX1 g7763(.Y(n_90), .A(n_88));
  ADDFX1 g7764(.CO(n_88), .S(n_89), .A(in_8[1]), .B(in_58[1]), .CI(in_1[1]));
  ADDFX1 g7765(.CO(n_86), .S(n_87), .A(n_14), .B(n_1), .CI(in_75[0]));
  ADDFX1 g7766(.CO(n_84), .S(n_85), .A(in_37), .B(in_62[0]), .CI(n_0));
  ADDFX1 g7767(.CO(n_82), .S(n_83), .A(in_27[0]), .B(in_51[0]), .CI(n_18));
  INVX1 g7768(.Y(n_81), .A(n_73));
  INVX1 g7769(.Y(n_80), .A(n_72));
  INVX1 g7770(.Y(n_79), .A(n_63));
  INVX1 g7771(.Y(n_78), .A(n_62));
  INVX1 g7772(.Y(n_77), .A(n_55));
  INVX1 g7773(.Y(n_76), .A(n_54));
  INVX1 g7774(.Y(n_75), .A(n_39));
  INVX1 g7775(.Y(n_74), .A(n_38));
  ADDFX1 g7776(.CO(n_72), .S(n_73), .A(in_29[1]), .B(in_21[1]), .CI(in_19[1]));
  ADDFX1 g7777(.CO(n_70), .S(n_71), .A(in_69[0]), .B(in_25[0]), .CI(in_19[0]));
  ADDFX1 g7778(.CO(n_68), .S(n_69), .A(in_56[1]), .B(in_36[1]), .CI(in_67[1]));
  ADDFX1 g7779(.CO(n_66), .S(n_67), .A(in_47), .B(n_19), .CI(in_73[0]));
  ADDFX1 g7780(.CO(n_64), .S(n_65), .A(in_24[0]), .B(n_13), .CI(in_55[0]));
  ADDFX1 g7781(.CO(n_62), .S(n_63), .A(in_6[2]), .B(in_28[2]), .CI(in_24[2]));
  ADDFX1 g7782(.CO(n_60), .S(n_61), .A(in_18[0]), .B(in_44[0]), .CI(in_71[0]));
  ADDFX1 g7783(.CO(n_58), .S(n_59), .A(n_12), .B(in_28[1]), .CI(in_24[1]));
  ADDFX1 g7784(.CO(n_56), .S(n_57), .A(in_6[1]), .B(in_25[1]), .CI(in_12[1]));
  ADDFX1 g7785(.CO(n_54), .S(n_55), .A(in_26[1]), .B(in_7[1]), .CI(in_33[1]));
  ADDFX1 g7786(.CO(n_52), .S(n_53), .A(in_5[0]), .B(n_5), .CI(in_54[0]));
  ADDFX1 g7787(.CO(n_50), .S(n_51), .A(in_57[1]), .B(n_6), .CI(in_60[1]));
  ADDFX1 g7788(.CO(n_48), .S(n_49), .A(in_12[0]), .B(in_29[0]), .CI(in_21[0]));
  ADDFX1 g7789(.CO(n_46), .S(n_47), .A(in_38[0]), .B(in_26[0]), .CI(n_23));
  ADDFX1 g7790(.CO(n_44), .S(n_45), .A(in_9[0]), .B(in_16[0]), .CI(n_25));
  ADDFX1 g7791(.CO(n_42), .S(n_43), .A(n_7), .B(in_20[1]), .CI(n_10));
  ADDFX1 g7792(.CO(n_40), .S(n_41), .A(in_14[0]), .B(in_11[0]), .CI(in_68));
  ADDFX1 g7793(.CO(n_38), .S(n_39), .A(in_65[1]), .B(in_59[1]), .CI(in_72[1]));
  ADDFX1 g7794(.CO(n_36), .S(n_37), .A(in_48[1]), .B(n_3), .CI(n_20));
  ADDFX1 g7795(.CO(n_34), .S(n_35), .A(in_46[1]), .B(n_4), .CI(n_9));
  ADDFX1 g7796(.CO(n_32), .S(n_33), .A(in_70[0]), .B(in_33[0]), .CI(in_6[0]));
  ADDFX1 g7797(.CO(n_30), .S(n_31), .A(in_28[0]), .B(n_21), .CI(n_17));
  ADDFX1 g7798(.CO(n_28), .S(n_29), .A(in_34), .B(n_16), .CI(n_8));
  OAI21X1 g7799(.Y(n_27), .A0(in_55[0]), .A1(in_11[0]), .B0(n_26));
  NAND2X1 g7800(.Y(n_26), .A(in_55[0]), .B(in_11[0]));
  INVX1 g7801(.Y(n_25), .A(in_49[0]));
  INVX1 g7802(.Y(n_24), .A(in_66[0]));
  INVX1 g7803(.Y(n_23), .A(in_45[0]));
  INVX1 g7804(.Y(n_22), .A(in_63[0]));
  INVX1 g7805(.Y(n_21), .A(in_31[0]));
  INVX1 g7806(.Y(n_20), .A(in_74[1]));
  INVX1 g7807(.Y(n_19), .A(in_64[0]));
  INVX1 g7808(.Y(n_18), .A(in_17[0]));
  INVX1 g7809(.Y(n_17), .A(in_13[0]));
  INVX1 g7810(.Y(n_16), .A(in_30[0]));
  INVX1 g7811(.Y(n_15), .A(in_4[2]));
  INVX1 g7812(.Y(n_14), .A(in_0[0]));
  INVX1 g7813(.Y(n_13), .A(in_41[0]));
  INVX1 g7814(.Y(n_12), .A(in_70[0]));
  INVX1 g7815(.Y(n_11), .A(in_2[7]));
  INVX1 g7816(.Y(n_10), .A(in_50[1]));
  INVX1 g7817(.Y(n_9), .A(in_61[1]));
  INVX1 g7818(.Y(n_8), .A(in_52[0]));
  INVX1 g7819(.Y(n_7), .A(in_10[1]));
  INVX1 g7820(.Y(n_6), .A(in_43[1]));
  INVX1 g7821(.Y(n_5), .A(in_22[0]));
  INVX1 g7822(.Y(n_4), .A(in_32[1]));
  INVX1 g7823(.Y(n_3), .A(in_53[1]));
  INVX1 g7824(.Y(n_2), .A(in_23[0]));
  INVX1 g7825(.Y(n_1), .A(in_40[0]));
  INVX1 g7826(.Y(n_0), .A(in_42[0]));
endmodule

module WALLACE_CSA_DUMMY_OP149_group_109835(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, out_0);
input  in_22, in_23, in_27;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [2:0] in_5;
input   [9:0] in_6;
input   [9:0] in_7;
input   [6:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [1:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [2:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [4:0] in_40;
input   [2:0] in_41;
input   [2:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
output  [9:0] out_0;
wire  n_157, n_154, n_152, n_150, n_149, n_148, n_147, n_146, n_145, n_144, 
    n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_135, n_134, n_133, 
    n_132, n_131, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, 
    n_111, n_110, n_109, n_108, n_107, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, n_0, in_27, in_23, in_22;
wire   [9:0] out_0;
wire   [1:0] in_37;
wire   [1:0] in_31;
wire   [1:0] in_29;
wire   [1:0] in_28;
wire   [1:0] in_24;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [6:0] in_8;
wire   [9:0] in_7;
wire   [9:0] in_6;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_30;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_42;
wire   [2:0] in_41;
wire   [2:0] in_39;
wire   [2:0] in_34;
wire   [2:0] in_32;
wire   [2:0] in_5;
wire   [2:0] in_3;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  OAI21X1 g4956(.Y(out_0[9]), .A0(n_143), .A1(n_157), .B0(n_144));
  XNOR2X1 g4957(.Y(out_0[7]), .A(n_145), .B(n_157));
  ADDFX1 g4958(.CO(n_157), .S(out_0[6]), .A(n_146), .B(n_141), .CI(n_154));
  ADDFX1 g4959(.CO(n_154), .S(out_0[5]), .A(n_148), .B(n_147), .CI(n_152));
  ADDFX1 g4960(.CO(n_152), .S(out_0[4]), .A(n_137), .B(n_149), .CI(n_150));
  ADDFX1 g4961(.CO(n_150), .S(out_0[3]), .A(n_135), .B(n_138), .CI(n_126));
  ADDFX1 g4962(.CO(n_148), .S(n_149), .A(n_140), .B(in_6[4]), .CI(n_125));
  ADDFX1 g4963(.CO(n_146), .S(n_147), .A(n_124), .B(n_139), .CI(in_6[5]));
  NAND2BX1 g4964(.Y(n_145), .AN(n_143), .B(n_144));
  NAND2BX1 g4965(.Y(n_144), .AN(n_142), .B(in_6[7]));
  NOR2BX1 g4966(.Y(n_143), .AN(n_142), .B(in_6[7]));
  ADDFX1 g4967(.CO(n_142), .S(n_141), .A(n_11), .B(n_123), .CI(in_6[6]));
  ADDFX1 g4968(.CO(n_139), .S(n_140), .A(n_111), .B(n_121), .CI(n_133));
  ADDFX1 g4969(.CO(n_137), .S(n_138), .A(n_134), .B(n_127), .CI(n_131));
  ADDFX1 g4970(.CO(n_135), .S(out_0[2]), .A(n_129), .B(n_128), .CI(n_132));
  ADDFX1 g4971(.CO(n_133), .S(n_134), .A(n_108), .B(n_119), .CI(n_109));
  ADDFX1 g4972(.CO(n_131), .S(n_132), .A(n_120), .B(n_110), .CI(in_6[2]));
  ADDFX1 g4973(.CO(n_129), .S(out_0[1]), .A(n_116), .B(n_105), .CI(n_118));
  ADDFX1 g4974(.CO(n_127), .S(n_128), .A(n_115), .B(n_114), .CI(n_117));
  ADDFX1 g4975(.CO(n_125), .S(n_126), .A(n_113), .B(n_112), .CI(in_6[3]));
  OAI2BB1X1 g4976(.Y(n_124), .A0N(in_7[5]), .A1N(n_122), .B0(n_123));
  OR2X1 g4977(.Y(n_123), .A(in_7[5]), .B(n_122));
  ADDFX1 g4978(.CO(n_122), .S(n_121), .A(n_85), .B(n_107), .CI(in_7[4]));
  ADDFX1 g4979(.CO(n_119), .S(n_120), .A(n_94), .B(n_88), .CI(n_101));
  ADDFX1 g4980(.CO(n_117), .S(n_118), .A(n_91), .B(n_104), .CI(in_6[1]));
  ADDFX1 g4981(.CO(n_115), .S(n_116), .A(n_102), .B(n_96), .CI(n_89));
  ADDFX1 g4982(.CO(n_113), .S(n_114), .A(n_98), .B(n_95), .CI(n_103));
  ADDFX1 g4983(.CO(n_111), .S(n_112), .A(n_93), .B(n_97), .CI(in_7[3]));
  ADDFX1 g4984(.CO(n_109), .S(n_110), .A(n_81), .B(n_99), .CI(in_7[2]));
  ADDFX1 g4985(.CO(n_107), .S(n_108), .A(n_83), .B(n_86), .CI(n_87));
  ADDHX1 g4986(.CO(n_105), .S(out_0[0]), .A(n_90), .B(n_92));
  ADDFX1 g4987(.CO(n_103), .S(n_104), .A(n_78), .B(n_100), .CI(in_7[1]));
  ADDFX1 g4988(.CO(n_101), .S(n_102), .A(n_79), .B(n_72), .CI(n_67));
  ADDFX1 g4989(.CO(n_99), .S(n_100), .A(n_61), .B(n_70), .CI(n_74));
  ADDFX1 g4990(.CO(n_97), .S(n_98), .A(n_65), .B(n_84), .CI(n_77));
  ADDFX1 g4991(.CO(n_95), .S(n_96), .A(n_66), .B(n_75), .CI(n_82));
  ADDFX1 g4992(.CO(n_93), .S(n_94), .A(n_73), .B(n_69), .CI(n_64));
  ADDFX1 g4993(.CO(n_91), .S(n_92), .A(n_80), .B(n_76), .CI(in_6[0]));
  ADDFX1 g4994(.CO(n_89), .S(n_90), .A(n_62), .B(n_68), .CI(in_7[0]));
  ADDFX1 g4995(.CO(n_87), .S(n_88), .A(n_71), .B(n_58), .CI(n_31));
  ADDFX1 g4996(.CO(n_85), .S(n_86), .A(n_18), .B(n_57), .CI(n_63));
  ADDFX1 g4997(.CO(n_83), .S(n_84), .A(n_37), .B(n_59), .CI(n_53));
  ADDFX1 g4998(.CO(n_81), .S(n_82), .A(n_55), .B(n_54), .CI(n_32));
  ADDFX1 g4999(.CO(n_79), .S(n_80), .A(n_46), .B(n_30), .CI(n_48));
  ADDFX1 g5000(.CO(n_77), .S(n_78), .A(n_22), .B(n_60), .CI(n_27));
  ADDFX1 g5001(.CO(n_75), .S(n_76), .A(n_34), .B(n_28), .CI(n_56));
  ADDFX1 g5002(.CO(n_73), .S(n_74), .A(n_17), .B(n_49), .CI(n_23));
  ADDFX1 g5003(.CO(n_71), .S(n_72), .A(n_25), .B(n_47), .CI(n_33));
  ADDFX1 g5004(.CO(n_69), .S(n_70), .A(n_45), .B(n_43), .CI(n_29));
  ADDFX1 g5005(.CO(n_67), .S(n_68), .A(n_44), .B(n_24), .CI(n_26));
  ADDFX1 g5006(.CO(n_65), .S(n_66), .A(n_40), .B(n_36), .CI(n_38));
  ADDFX1 g5007(.CO(n_63), .S(n_64), .A(n_39), .B(n_35), .CI(n_21));
  ADDFX1 g5008(.CO(n_61), .S(n_62), .A(in_10[0]), .B(n_20), .CI(n_50));
  ADDFX1 g5009(.CO(n_59), .S(n_60), .A(in_12[0]), .B(in_20[1]), .CI(n_9));
  ADDFX1 g5010(.CO(n_57), .S(n_58), .A(in_34[0]), .B(n_1), .CI(n_19));
  ADDFX1 g5011(.CO(n_55), .S(n_56), .A(in_13[0]), .B(in_19[0]), .CI(in_11[0]));
  INVX1 g5012(.Y(n_54), .A(n_52));
  INVX1 g5013(.Y(n_53), .A(n_51));
  ADDFX1 g5014(.CO(n_51), .S(n_52), .A(in_10[1]), .B(in_11[1]), .CI(in_19[1]));
  ADDFX1 g5015(.CO(n_49), .S(n_50), .A(in_29[0]), .B(n_5), .CI(in_31[0]));
  ADDFX1 g5016(.CO(n_47), .S(n_48), .A(in_28[0]), .B(in_34[0]), .CI(in_37[0]));
  ADDFX1 g5017(.CO(n_45), .S(n_46), .A(n_12), .B(n_10), .CI(in_38[0]));
  INVX1 g5018(.Y(n_44), .A(n_42));
  INVX1 g5019(.Y(n_43), .A(n_41));
  ADDFX1 g5020(.CO(n_41), .S(n_42), .A(in_35[0]), .B(in_14[0]), .CI(in_40[0]));
  ADDFX1 g5021(.CO(n_39), .S(n_40), .A(in_3[1]), .B(in_0[1]), .CI(in_39[1]));
  ADDFX1 g5022(.CO(n_37), .S(n_38), .A(in_5[1]), .B(n_14), .CI(n_15));
  ADDFX1 g5023(.CO(n_35), .S(n_36), .A(in_17[1]), .B(n_2), .CI(in_32[1]));
  ADDFX1 g5024(.CO(n_33), .S(n_34), .A(in_15[0]), .B(in_27), .CI(n_16));
  ADDFX1 g5025(.CO(n_31), .S(n_32), .A(n_0), .B(n_13), .CI(in_13[1]));
  ADDFX1 g5026(.CO(n_29), .S(n_30), .A(in_12[0]), .B(n_8), .CI(in_44[0]));
  ADDFX1 g5027(.CO(n_27), .S(n_28), .A(in_9[0]), .B(in_16[0]), .CI(in_20[0]));
  ADDFX1 g5028(.CO(n_25), .S(n_26), .A(n_3), .B(n_4), .CI(in_22));
  ADDFX1 g5029(.CO(n_23), .S(n_24), .A(in_23), .B(n_7), .CI(in_41[0]));
  ADDFX1 g5030(.CO(n_21), .S(n_22), .A(in_41[0]), .B(in_28[0]), .CI(in_42[1]));
  OAI2BB1X1 g5031(.Y(n_20), .A0N(in_24[0]), .A1N(n_6), .B0(n_17));
  XOR2XL g5032(.Y(n_19), .A(in_38[0]), .B(in_44[0]));
  NOR2X1 g5033(.Y(n_18), .A(in_44[0]), .B(in_38[0]));
  OR2X1 g5034(.Y(n_17), .A(in_24[0]), .B(n_6));
  INVX1 g5035(.Y(n_16), .A(in_36[0]));
  INVX1 g5036(.Y(n_15), .A(in_43[1]));
  INVX1 g5037(.Y(n_14), .A(in_21[1]));
  INVX1 g5038(.Y(n_13), .A(in_9[1]));
  INVX1 g5039(.Y(n_12), .A(in_26[0]));
  INVX1 g5040(.Y(n_11), .A(in_7[6]));
  INVX1 g5041(.Y(n_10), .A(in_25[0]));
  INVX1 g5042(.Y(n_9), .A(in_16[1]));
  INVX1 g5043(.Y(n_8), .A(in_30[0]));
  INVX1 g5044(.Y(n_7), .A(in_8[0]));
  INVX1 g5045(.Y(n_6), .A(in_33[0]));
  INVX1 g5046(.Y(n_5), .A(in_18[0]));
  INVX1 g5047(.Y(n_4), .A(in_4[0]));
  INVX1 g5048(.Y(n_3), .A(in_1[0]));
  INVX1 g5049(.Y(n_2), .A(in_2[1]));
  INVX1 g5050(.Y(n_1), .A(in_13[2]));
  INVX1 g5051(.Y(n_0), .A(in_34[0]));
endmodule

module WALLACE_CSA_DUMMY_OP150_group_109838_6295(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, out_0);
input  in_32, in_41, in_42, in_44;
input   [4:0] in_0;
input   [9:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [1:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [1:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
input   [1:0] in_43;
input   [4:0] in_45;
input   [1:0] in_46;
output  [9:0] out_0;
wire  n_164, n_162, n_160, n_158, n_156, n_155, n_154, n_153, n_152, n_151, 
    n_150, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, 
    n_139, n_138, n_137, n_136, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_44, 
    in_42, in_41, in_32;
wire   [9:0] out_0;
wire   [2:0] in_30;
wire   [1:0] in_46;
wire   [1:0] in_43;
wire   [1:0] in_40;
wire   [1:0] in_38;
wire   [1:0] in_34;
wire   [1:0] in_33;
wire   [1:0] in_22;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [9:0] in_1;
wire   [4:0] in_45;
wire   [4:0] in_39;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g5246(.Y(out_0[9]), .A(n_164));
  ADDFX1 g5247(.CO(n_164), .S(out_0[7]), .A(n_37), .B(n_144), .CI(n_162));
  ADDFX1 g5248(.CO(n_162), .S(out_0[6]), .A(n_145), .B(n_152), .CI(n_160));
  ADDFX1 g5249(.CO(n_160), .S(out_0[5]), .A(n_153), .B(n_154), .CI(n_158));
  ADDFX1 g5250(.CO(n_158), .S(out_0[4]), .A(n_150), .B(n_155), .CI(n_156));
  ADDFX1 g5251(.CO(n_156), .S(out_0[3]), .A(n_140), .B(n_148), .CI(n_151));
  ADDFX1 g5252(.CO(n_154), .S(n_155), .A(n_131), .B(n_136), .CI(n_147));
  ADDFX1 g5253(.CO(n_152), .S(n_153), .A(n_130), .B(n_133), .CI(n_146));
  ADDFX1 g5254(.CO(n_150), .S(n_151), .A(n_143), .B(n_138), .CI(n_137));
  ADDFX1 g5255(.CO(n_148), .S(out_0[2]), .A(n_139), .B(n_134), .CI(n_141));
  ADDFX1 g5256(.CO(n_146), .S(n_147), .A(n_120), .B(n_142), .CI(n_119));
  ADDFX1 g5257(.CO(n_144), .S(n_145), .A(n_106), .B(n_38), .CI(n_132));
  ADDFX1 g5258(.CO(n_142), .S(n_143), .A(n_108), .B(n_128), .CI(n_115));
  ADDFX1 g5259(.CO(n_140), .S(n_141), .A(n_117), .B(n_125), .CI(n_122));
  ADDFX1 g5260(.CO(n_138), .S(n_139), .A(n_109), .B(n_126), .CI(n_129));
  ADDFX1 g5261(.CO(n_136), .S(n_137), .A(n_116), .B(n_124), .CI(n_121));
  ADDFX1 g5262(.CO(n_134), .S(out_0[1]), .A(n_112), .B(n_127), .CI(n_123));
  ADDFX1 g5263(.CO(n_132), .S(n_133), .A(in_3[5]), .B(n_118), .CI(n_107));
  ADDFX1 g5264(.CO(n_130), .S(n_131), .A(in_2[4]), .B(in_1[4]), .CI(n_114));
  ADDFX1 g5265(.CO(n_128), .S(n_129), .A(n_102), .B(in_2[2]), .CI(in_1[2]));
  ADDFX1 g5266(.CO(n_126), .S(n_127), .A(n_103), .B(n_97), .CI(n_100));
  ADDFX1 g5267(.CO(n_124), .S(n_125), .A(in_3[2]), .B(n_98), .CI(n_110));
  ADDFX1 g5268(.CO(n_122), .S(n_123), .A(n_94), .B(n_99), .CI(n_111));
  ADDFX1 g5269(.CO(n_120), .S(n_121), .A(n_105), .B(in_2[3]), .CI(in_3[3]));
  ADDFX1 g5270(.CO(n_118), .S(n_119), .A(n_87), .B(n_104), .CI(in_3[4]));
  ADDFX1 g5271(.CO(n_116), .S(n_117), .A(n_88), .B(n_96), .CI(n_93));
  ADDFX1 g5272(.CO(n_114), .S(n_115), .A(n_85), .B(n_92), .CI(in_1[3]));
  ADDHX1 g5273(.CO(n_112), .S(out_0[0]), .A(n_95), .B(n_101));
  ADDFX1 g5274(.CO(n_110), .S(n_111), .A(n_89), .B(n_65), .CI(in_3[1]));
  ADDFX1 g5275(.CO(n_108), .S(n_109), .A(n_74), .B(n_69), .CI(n_91));
  ADDFX1 g5276(.CO(n_106), .S(n_107), .A(n_86), .B(in_2[5]), .CI(in_1[5]));
  ADDFX1 g5277(.CO(n_104), .S(n_105), .A(n_79), .B(n_73), .CI(n_90));
  ADDFX1 g5278(.CO(n_102), .S(n_103), .A(n_75), .B(n_77), .CI(n_81));
  ADDFX1 g5279(.CO(n_100), .S(n_101), .A(n_78), .B(n_82), .CI(in_2[0]));
  ADDFX1 g5280(.CO(n_98), .S(n_99), .A(n_72), .B(in_2[1]), .CI(in_1[1]));
  ADDFX1 g5281(.CO(n_96), .S(n_97), .A(n_64), .B(n_62), .CI(n_70));
  ADDFX1 g5282(.CO(n_94), .S(n_95), .A(n_76), .B(in_3[0]), .CI(n_66));
  ADDFX1 g5283(.CO(n_92), .S(n_93), .A(n_68), .B(n_80), .CI(n_71));
  ADDFX1 g5284(.CO(n_90), .S(n_91), .A(n_63), .B(n_83), .CI(n_61));
  ADDFX1 g5285(.CO(n_88), .S(n_89), .A(n_29), .B(n_56), .CI(n_84));
  INVX1 g5286(.Y(n_87), .A(n_86));
  ADDFX1 g5287(.CO(n_86), .S(n_85), .A(n_13), .B(n_20), .CI(n_67));
  ADDFX1 g5288(.CO(n_83), .S(n_84), .A(n_43), .B(n_57), .CI(n_59));
  ADDFX1 g5289(.CO(n_81), .S(n_82), .A(n_16), .B(n_24), .CI(n_50));
  ADDFX1 g5290(.CO(n_79), .S(n_80), .A(n_15), .B(n_53), .CI(n_45));
  ADDFX1 g5291(.CO(n_77), .S(n_78), .A(n_40), .B(n_58), .CI(n_60));
  ADDFX1 g5292(.CO(n_75), .S(n_76), .A(in_9[0]), .B(n_28), .CI(n_44));
  ADDFX1 g5293(.CO(n_73), .S(n_74), .A(n_21), .B(n_25), .CI(n_55));
  ADDFX1 g5294(.CO(n_71), .S(n_72), .A(n_48), .B(n_46), .CI(n_54));
  ADDFX1 g5295(.CO(n_69), .S(n_70), .A(n_17), .B(n_34), .CI(n_26));
  ADDFX1 g5296(.CO(n_67), .S(n_68), .A(n_12), .B(n_47), .CI(n_33));
  ADDFX1 g5297(.CO(n_65), .S(n_66), .A(n_22), .B(n_30), .CI(in_1[0]));
  ADDFX1 g5298(.CO(n_63), .S(n_64), .A(n_10), .B(n_23), .CI(n_27));
  ADDFX1 g5299(.CO(n_61), .S(n_62), .A(n_19), .B(n_49), .CI(n_39));
  ADDFX1 g5300(.CO(n_59), .S(n_60), .A(in_44), .B(in_40[0]), .CI(in_46[0]));
  ADDFX1 g5301(.CO(n_57), .S(n_58), .A(in_42), .B(n_6), .CI(in_43[0]));
  ADDFX1 g5302(.CO(n_55), .S(n_56), .A(in_12[1]), .B(n_5), .CI(in_16[1]));
  INVX1 g5303(.Y(n_54), .A(n_52));
  INVX1 g5304(.Y(n_53), .A(n_51));
  ADDFX1 g5305(.CO(n_51), .S(n_52), .A(in_27[1]), .B(in_15[1]), .CI(in_31[1]));
  ADDFX1 g5306(.CO(n_49), .S(n_50), .A(in_4[0]), .B(in_38[0]), .CI(n_0));
  ADDFX1 g5307(.CO(n_47), .S(n_48), .A(in_33[0]), .B(in_13[1]), .CI(n_9));
  ADDFX1 g5308(.CO(n_45), .S(n_46), .A(in_30[1]), .B(n_3), .CI(n_1));
  INVX1 g5309(.Y(n_44), .A(n_42));
  INVX1 g5310(.Y(n_43), .A(n_41));
  ADDFX1 g5311(.CO(n_41), .S(n_42), .A(in_6[0]), .B(in_21[0]), .CI(in_23[0]));
  ADDFX1 g5312(.CO(n_39), .S(n_40), .A(in_16[0]), .B(in_19[0]), .CI(n_4));
  INVX1 g5313(.Y(n_38), .A(n_36));
  INVX1 g5314(.Y(n_37), .A(n_35));
  ADDFX1 g5315(.CO(n_35), .S(n_36), .A(in_2[6]), .B(in_1[6]), .CI(in_3[6]));
  INVX1 g5316(.Y(n_34), .A(n_32));
  INVX1 g5317(.Y(n_33), .A(n_31));
  ADDFX1 g5318(.CO(n_31), .S(n_32), .A(in_17[1]), .B(in_24[1]), .CI(in_37[1]));
  ADDFX1 g5319(.CO(n_29), .S(n_30), .A(in_5[0]), .B(in_12[0]), .CI(in_11[0]));
  ADDFX1 g5320(.CO(n_27), .S(n_28), .A(n_7), .B(n_2), .CI(in_34[0]));
  ADDFX1 g5321(.CO(n_25), .S(n_26), .A(in_43[0]), .B(in_5[1]), .CI(n_8));
  ADDFX1 g5322(.CO(n_23), .S(n_24), .A(in_22[0]), .B(in_41), .CI(in_33[0]));
  XNOR2X1 g5323(.Y(n_22), .A(in_18[0]), .B(n_14));
  XOR2XL g5324(.Y(n_21), .A(in_16[2]), .B(n_14));
  OAI22X1 g5325(.Y(n_20), .A0(in_29[0]), .A1(n_11), .B0(in_26[0]), .B1(in_16[2]));
  OAI2BB1X1 g5326(.Y(n_19), .A0N(in_18[0]), .A1N(in_26[0]), .B0(n_18));
  OAI21XL g5327(.Y(n_18), .A0(in_18[0]), .A1(in_26[0]), .B0(in_29[0]));
  OAI21X1 g5328(.Y(n_17), .A0(in_28[1]), .A1(in_25[1]), .B0(n_12));
  OAI2BB1X1 g5329(.Y(n_16), .A0N(in_32), .A1N(in_7[0]), .B0(n_10));
  XNOR2X1 g5330(.Y(n_15), .A(in_14[2]), .B(in_45[2]));
  XNOR2X1 g5331(.Y(n_14), .A(in_26[0]), .B(in_29[0]));
  NOR2BX1 g5332(.Y(n_13), .AN(in_14[2]), .B(in_45[2]));
  NAND2X1 g5333(.Y(n_12), .A(in_28[1]), .B(in_25[1]));
  AND2XL g5334(.Y(n_11), .A(in_26[0]), .B(in_16[2]));
  OR2X1 g5335(.Y(n_10), .A(in_32), .B(in_7[0]));
  INVX1 g5336(.Y(n_9), .A(in_35[1]));
  INVX1 g5337(.Y(n_8), .A(in_11[1]));
  INVX1 g5338(.Y(n_7), .A(in_20[0]));
  INVX1 g5339(.Y(n_6), .A(in_0[0]));
  INVX1 g5340(.Y(n_5), .A(in_9[1]));
  INVX1 g5341(.Y(n_4), .A(in_39[0]));
  INVX1 g5342(.Y(n_3), .A(in_36[1]));
  INVX1 g5343(.Y(n_2), .A(in_10[0]));
  INVX1 g5344(.Y(n_1), .A(in_18[1]));
  INVX1 g5345(.Y(n_0), .A(in_8[0]));
endmodule

module WALLACE_CSA_DUMMY_OP150_group_109838(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, out_0);
input  in_22;
input   [4:0] in_0;
input   [2:0] in_1;
input   [4:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [1:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [2:0] in_19;
input   [1:0] in_20;
input   [4:0] in_21;
input   [1:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [1:0] in_30;
input   [1:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [1:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
output  [9:0] out_0;
wire  n_113, n_111, n_109, n_107, n_106, n_105, n_104, n_103, n_101, n_100, n_99, 
    n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_0, in_22;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_38;
wire   [1:0] in_32;
wire   [1:0] in_31;
wire   [1:0] in_30;
wire   [1:0] in_25;
wire   [1:0] in_23;
wire   [1:0] in_20;
wire   [1:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [2:0] in_34;
wire   [2:0] in_19;
wire   [2:0] in_1;
wire   [4:0] in_39;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_21;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_2;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1281(.Y(out_0[9]), .A(n_113));
  ADDFX1 g1282(.CO(n_113), .S(out_0[5]), .A(n_74), .B(n_99), .CI(n_111));
  ADDFX1 g1283(.CO(n_111), .S(out_0[4]), .A(n_100), .B(n_105), .CI(n_109));
  ADDFX1 g1284(.CO(n_109), .S(out_0[3]), .A(n_103), .B(n_106), .CI(n_107));
  ADDFX1 g1285(.CO(n_107), .S(out_0[2]), .A(n_93), .B(n_101), .CI(n_104));
  ADDFX1 g1286(.CO(n_105), .S(n_106), .A(n_91), .B(n_97), .CI(n_96));
  ADDFX1 g1287(.CO(n_103), .S(n_104), .A(n_71), .B(n_98), .CI(n_92));
  ADDFX1 g1288(.CO(n_101), .S(out_0[1]), .A(n_72), .B(n_83), .CI(n_94));
  ADDFX1 g1289(.CO(n_99), .S(n_100), .A(n_0), .B(n_89), .CI(n_95));
  ADDFX1 g1290(.CO(n_97), .S(n_98), .A(n_80), .B(n_85), .CI(n_88));
  ADDFX1 g1291(.CO(n_95), .S(n_96), .A(n_79), .B(n_87), .CI(n_90));
  ADDFX1 g1292(.CO(n_93), .S(n_94), .A(n_61), .B(n_86), .CI(n_78));
  ADDFX1 g1293(.CO(n_91), .S(n_92), .A(n_51), .B(n_77), .CI(n_82));
  ADDFX1 g1294(.CO(n_89), .S(n_90), .A(n_73), .B(n_75), .CI(n_81));
  ADDFX1 g1295(.CO(n_87), .S(n_88), .A(n_36), .B(n_26), .CI(n_76));
  ADDFX1 g1296(.CO(n_85), .S(n_86), .A(n_50), .B(n_69), .CI(n_66));
  ADDFX1 g1297(.CO(n_83), .S(out_0[0]), .A(n_54), .B(n_62), .CI(n_70));
  ADDFX1 g1298(.CO(n_81), .S(n_82), .A(n_32), .B(n_28), .CI(n_67));
  ADDFX1 g1299(.CO(n_79), .S(n_80), .A(n_49), .B(n_57), .CI(n_65));
  ADDFX1 g1300(.CO(n_77), .S(n_78), .A(n_34), .B(n_27), .CI(n_64));
  ADDFX1 g1301(.CO(n_75), .S(n_76), .A(n_12), .B(in_4[2]), .CI(n_63));
  INVX1 g1302(.Y(n_74), .A(n_0));
  XNOR2X1 g1303(.Y(n_73), .A(n_39), .B(n_68));
  ADDFX1 g1304(.CO(n_71), .S(n_72), .A(n_58), .B(n_53), .CI(n_52));
  ADDFX1 g1306(.CO(n_69), .S(n_70), .A(in_13[0]), .B(n_44), .CI(n_60));
  ADDFX1 g1307(.CO(n_68), .S(n_67), .A(n_2), .B(n_39), .CI(n_55));
  ADDFX1 g1308(.CO(n_65), .S(n_66), .A(n_22), .B(n_47), .CI(n_59));
  ADDFX1 g1309(.CO(n_63), .S(n_64), .A(n_7), .B(in_31[1]), .CI(n_56));
  ADDFX1 g1310(.CO(n_61), .S(n_62), .A(n_48), .B(n_25), .CI(n_35));
  ADDFX1 g1311(.CO(n_59), .S(n_60), .A(n_16), .B(in_8[0]), .CI(n_21));
  ADDFX1 g1312(.CO(n_57), .S(n_58), .A(n_45), .B(n_24), .CI(n_43));
  ADDFX1 g1313(.CO(n_55), .S(n_56), .A(n_18), .B(n_20), .CI(n_40));
  ADDFX1 g1314(.CO(n_53), .S(n_54), .A(n_23), .B(n_42), .CI(n_46));
  ADDFX1 g1315(.CO(n_51), .S(n_52), .A(n_37), .B(n_29), .CI(n_33));
  ADDFX1 g1316(.CO(n_49), .S(n_50), .A(n_8), .B(in_4[1]), .CI(n_41));
  ADDFX1 g1317(.CO(n_47), .S(n_48), .A(in_15[0]), .B(in_38[0]), .CI(n_3));
  ADDFX1 g1318(.CO(n_45), .S(n_46), .A(n_10), .B(in_40[0]), .CI(n_14));
  ADDFX1 g1319(.CO(n_43), .S(n_44), .A(in_25[0]), .B(in_32[0]), .CI(in_36[0]));
  ADDFX1 g1320(.CO(n_41), .S(n_42), .A(n_9), .B(n_15), .CI(in_30[0]));
  INVX1 g1321(.Y(n_40), .A(n_38));
  ADDFX1 g1323(.CO(n_39), .S(n_38), .A(in_9[1]), .B(in_10[1]), .CI(in_11[1]));
  ADDFX1 g1324(.CO(n_36), .S(n_37), .A(in_23[1]), .B(n_4), .CI(in_32[0]));
  ADDFX1 g1325(.CO(n_34), .S(n_35), .A(in_4[0]), .B(in_7[0]), .CI(in_6[0]));
  INVX1 g1326(.Y(n_33), .A(n_31));
  INVX1 g1327(.Y(n_32), .A(n_30));
  ADDFX1 g1328(.CO(n_30), .S(n_31), .A(in_21[1]), .B(in_29[1]), .CI(in_39[1]));
  ADDFX1 g1329(.CO(n_28), .S(n_29), .A(in_1[1]), .B(in_19[1]), .CI(n_11));
  ADDFX1 g1330(.CO(n_26), .S(n_27), .A(in_34[1]), .B(n_6), .CI(n_13));
  ADDFX1 g1331(.CO(n_24), .S(n_25), .A(in_16[0]), .B(n_5), .CI(n_17));
  ADDFX1 g1332(.CO(n_22), .S(n_23), .A(in_3[0]), .B(in_20[0]), .CI(in_22));
  OAI21X1 g1333(.Y(n_21), .A0(in_12[0]), .A1(n_19), .B0(n_20));
  NAND2X1 g1334(.Y(n_20), .A(in_12[0]), .B(n_19));
  XNOR2X1 g1335(.Y(n_19), .A(in_5[0]), .B(in_14[0]));
  NOR2X1 g1336(.Y(n_18), .A(in_14[0]), .B(in_5[0]));
  INVX1 g1337(.Y(n_17), .A(in_37[0]));
  INVX1 g1338(.Y(n_16), .A(in_27[0]));
  INVX1 g1339(.Y(n_15), .A(in_24[0]));
  INVX1 g1340(.Y(n_14), .A(in_18[0]));
  INVX1 g1341(.Y(n_13), .A(in_6[1]));
  INVX1 g1342(.Y(n_12), .A(in_36[0]));
  INVX1 g1343(.Y(n_11), .A(in_35[1]));
  INVX1 g1344(.Y(n_10), .A(in_17[0]));
  INVX1 g1345(.Y(n_9), .A(in_0[0]));
  INVX1 g1346(.Y(n_8), .A(in_7[1]));
  INVX1 g1347(.Y(n_7), .A(in_26[1]));
  INVX1 g1348(.Y(n_6), .A(in_13[1]));
  INVX1 g1349(.Y(n_5), .A(in_33[0]));
  INVX1 g1350(.Y(n_4), .A(in_2[1]));
  INVX1 g1351(.Y(n_3), .A(in_28[0]));
  INVX1 g1352(.Y(n_2), .A(in_16[0]));
  NAND2BX1 g2(.Y(n_0), .AN(n_39), .B(n_68));
endmodule

module WALLACE_CSA_DUMMY_OP154_group_109832(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, out_0);
input  in_37, in_39;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [6:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [1:0] in_20;
input   [4:0] in_21;
input   [2:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [2:0] in_26;
input   [1:0] in_27;
input   [1:0] in_28;
input   [2:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [2:0] in_35;
input   [4:0] in_36;
input   [1:0] in_38;
input   [1:0] in_40;
input   [2:0] in_41;
input   [4:0] in_42;
output  [9:0] out_0;
wire  n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, 
    n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_39, in_37;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_38;
wire   [1:0] in_28;
wire   [1:0] in_27;
wire   [1:0] in_20;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_5;
wire   [2:0] in_41;
wire   [2:0] in_35;
wire   [2:0] in_34;
wire   [2:0] in_29;
wire   [2:0] in_26;
wire   [2:0] in_22;
wire   [2:0] in_3;
wire   [4:0] in_42;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_110), .S(n_109), .A(n_3), .B(in_34[0]), .CI(n_9));
  ADDFX1 cdnfadd_000_1(.CO(n_108), .S(n_107), .A(n_15), .B(in_10[0]), .CI(
    in_41[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_106), .S(n_105), .A(in_39), .B(n_16), .CI(n_19));
  ADDFX1 cdnfadd_000_3(.CO(n_104), .S(n_103), .A(n_6), .B(in_17[0]), .CI(n_4));
  ADDFX1 cdnfadd_000_4(.CO(n_102), .S(n_101), .A(in_12[0]), .B(n_18), .CI(in_37));
  ADDFX1 cdnfadd_000_5(.CO(n_100), .S(n_99), .A(in_8[0]), .B(n_8), .CI(in_20[0]));
  ADDFX1 cdnfadd_000_6(.CO(n_98), .S(n_97), .A(in_28[0]), .B(n_2), .CI(in_26[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_96), .S(n_95), .A(n_12), .B(n_20), .CI(in_38[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_94), .S(n_93), .A(in_6[0]), .B(in_5[0]), .CI(
    in_16[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_76), .S(n_56), .A(in_2[0]), .B(in_7[0]), .CI(n_103));
  ADDFX1 cdnfadd_000_10(.CO(n_75), .S(n_111), .A(n_107), .B(n_109), .CI(n_95));
  ADDFX1 cdnfadd_000_11(.CO(n_74), .S(n_118), .A(n_97), .B(n_101), .CI(n_105));
  ADDFX1 cdnfadd_000_12(.CO(n_73), .S(n_112), .A(n_99), .B(n_93), .CI(n_56));
  ADDFX1 cdnfadd_001_0(.CO(n_77), .S(n_92), .A(in_38[0]), .B(in_12[0]), .CI(n_13));
  ADDFX1 cdnfadd_001_1(.CO(n_91), .S(n_90), .A(in_28[0]), .B(in_15[1]), .CI(
    in_40[1]));
  ADDFX1 cdnfadd_001_2(.CO(n_89), .S(n_88), .A(in_26[0]), .B(in_8[1]), .CI(n_17));
  ADDFX1 cdnfadd_001_3(.CO(n_87), .S(n_86), .A(in_35[1]), .B(in_22[1]), .CI(
    in_29[1]));
  ADDFX1 cdnfadd_001_4(.CO(n_85), .S(n_84), .A(in_14[1]), .B(in_27[1]), .CI(n_11));
  ADDFX1 cdnfadd_001_5(.CO(n_83), .S(n_82), .A(n_5), .B(in_41[0]), .CI(in_34[0]));
  ADDFX1 cdnfadd_001_6(.CO(n_81), .S(n_80), .A(in_3[1]), .B(n_1), .CI(n_7));
  ADDFX1 cdnfadd_001_7(.CO(n_79), .S(n_78), .A(n_14), .B(in_5[1]), .CI(in_7[1]));
  ADDFX1 cdnfadd_001_8(.CO(n_55), .S(n_72), .A(n_10), .B(n_108), .CI(n_100));
  ADDFX1 cdnfadd_001_9(.CO(n_71), .S(n_70), .A(n_102), .B(n_110), .CI(n_104));
  ADDFX1 cdnfadd_001_10(.CO(n_69), .S(n_68), .A(n_96), .B(n_98), .CI(n_106));
  ADDFX1 cdnfadd_001_11(.CO(n_67), .S(n_66), .A(n_80), .B(n_88), .CI(n_90));
  ADDFX1 cdnfadd_001_12(.CO(n_65), .S(n_64), .A(n_92), .B(n_84), .CI(n_86));
  ADDFX1 cdnfadd_001_13(.CO(n_63), .S(n_62), .A(n_82), .B(n_78), .CI(n_94));
  ADDFX1 cdnfadd_001_14(.CO(n_53), .S(n_52), .A(n_70), .B(n_75), .CI(n_68));
  ADDFX1 cdnfadd_001_15(.CO(n_51), .S(n_50), .A(n_74), .B(n_76), .CI(n_72));
  ADDFX1 cdnfadd_001_16(.CO(n_49), .S(n_119), .A(n_64), .B(n_66), .CI(n_62));
  ADDFX1 cdnfadd_001_17(.CO(n_120), .S(n_113), .A(n_73), .B(n_52), .CI(n_50));
  ADDFX1 cdnfadd_002_0(.CO(n_54), .S(n_61), .A(n_89), .B(n_87), .CI(n_91));
  ADDFX1 cdnfadd_002_1(.CO(n_60), .S(n_59), .A(n_81), .B(n_85), .CI(n_83));
  ADDFX1 cdnfadd_002_2(.CO(n_58), .S(n_57), .A(n_79), .B(n_21), .CI(n_55));
  ADDFX1 cdnfadd_002_3(.CO(n_48), .S(n_47), .A(n_71), .B(n_69), .CI(n_61));
  ADDFX1 cdnfadd_002_4(.CO(n_46), .S(n_45), .A(n_67), .B(n_65), .CI(n_59));
  ADDFX1 cdnfadd_002_5(.CO(n_42), .S(n_38), .A(n_63), .B(n_57), .CI(n_53));
  ADDFX1 cdnfadd_002_6(.CO(n_41), .S(n_37), .A(n_51), .B(n_47), .CI(n_45));
  ADDFX1 cdnfadd_002_7(.CO(n_121), .S(n_114), .A(n_49), .B(n_38), .CI(n_37));
  ADDFX1 cdnfadd_003_0(.CO(n_44), .S(n_43), .A(n_60), .B(n_24), .CI(n_58));
  ADDFX1 cdnfadd_003_1(.CO(n_40), .S(n_39), .A(n_48), .B(n_46), .CI(n_43));
  ADDFX1 cdnfadd_003_2(.CO(n_122), .S(n_115), .A(n_42), .B(n_41), .CI(n_39));
  ADDFX1 cdnfadd_004_0(.CO(n_117), .S(n_116), .A(n_23), .B(n_44), .CI(n_40));
  AO21XL g233(.Y(out_0[5]), .A0(n_117), .A1(n_34), .B0(out_0[9]));
  NOR2X1 g234(.Y(out_0[9]), .A(n_117), .B(n_34));
  ADDFX1 g235(.CO(n_34), .S(out_0[4]), .A(n_116), .B(n_122), .CI(n_31));
  ADDFX1 g236(.CO(n_31), .S(out_0[3]), .A(n_121), .B(n_115), .CI(n_29));
  ADDFX1 g237(.CO(n_29), .S(out_0[2]), .A(n_120), .B(n_27), .CI(n_114));
  ADDFX1 g238(.CO(n_27), .S(out_0[1]), .A(n_25), .B(n_119), .CI(n_113));
  ADDFX1 g239(.CO(n_25), .S(out_0[0]), .A(n_118), .B(n_111), .CI(n_112));
  AOI21X1 g240(.Y(n_24), .A0(n_21), .A1(n_22), .B0(n_23));
  NOR2X1 g241(.Y(n_23), .A(n_21), .B(n_22));
  INVX1 g242(.Y(n_22), .A(n_54));
  INVX1 g243(.Y(n_21), .A(n_77));
  INVX1 g244(.Y(n_20), .A(in_0[0]));
  INVX1 g245(.Y(n_19), .A(in_1[0]));
  INVX1 g246(.Y(n_18), .A(in_21[0]));
  INVX1 g247(.Y(n_17), .A(in_42[1]));
  INVX1 g248(.Y(n_16), .A(in_32[0]));
  INVX1 g249(.Y(n_15), .A(in_30[0]));
  INVX1 g250(.Y(n_14), .A(in_16[1]));
  INVX1 g251(.Y(n_13), .A(in_23[1]));
  INVX1 g252(.Y(n_12), .A(in_31[0]));
  INVX1 g253(.Y(n_11), .A(in_4[1]));
  INVX1 g254(.Y(n_10), .A(in_2[0]));
  INVX1 g255(.Y(n_9), .A(in_36[0]));
  INVX1 g256(.Y(n_8), .A(in_13[0]));
  INVX1 g257(.Y(n_7), .A(in_11[1]));
  INVX1 g258(.Y(n_6), .A(in_25[0]));
  INVX1 g259(.Y(n_5), .A(in_18[1]));
  INVX1 g260(.Y(n_4), .A(in_24[0]));
  INVX1 g261(.Y(n_3), .A(in_33[0]));
  INVX1 g262(.Y(n_2), .A(in_19[0]));
  INVX1 g263(.Y(n_1), .A(in_9[1]));
endmodule

module WALLACE_CSA_DUMMY_OP155_group_106213(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, out_0);
input  in_22, in_29, in_32, in_33, in_37, in_38, in_41, in_42, in_43, in_50, 
    in_51, in_63, in_65;
input   [4:0] in_0;
input   [4:0] in_1;
input   [2:0] in_2;
input   [9:0] in_3;
input   [9:0] in_4;
input   [5:0] in_5;
input   [4:0] in_6;
input   [4:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [4:0] in_20;
input   [5:0] in_21;
input   [1:0] in_23;
input   [2:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [1:0] in_27;
input   [1:0] in_28;
input   [2:0] in_30;
input   [3:0] in_31;
input   [2:0] in_34;
input   [1:0] in_35;
input   [1:0] in_36;
input   [1:0] in_39;
input   [1:0] in_40;
input   [2:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [1:0] in_47;
input   [1:0] in_48;
input   [4:0] in_49;
input   [4:0] in_52;
input   [1:0] in_53;
input   [1:0] in_54;
input   [4:0] in_55;
input   [4:0] in_56;
input   [4:0] in_57;
input   [2:0] in_58;
input   [4:0] in_59;
input   [1:0] in_60;
input   [1:0] in_61;
input   [1:0] in_62;
input   [1:0] in_64;
output  [9:0] out_0;
wire  n_213, n_210, n_208, n_206, n_204, n_203, n_202, n_201, n_200, n_199, 
    n_198, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, 
    n_187, n_186, n_185, n_184, n_183, n_182, n_180, n_179, n_178, n_177, 
    n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
    n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, 
    n_156, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, 
    n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, 
    n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, 
    n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, 
    n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, 
    n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, 
    n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, 
    n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, 
    n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, 
    n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, 
    n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, 
    n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, 
    n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_65, in_63, 
    in_51, in_50, in_43, in_42, in_41, in_38, in_37, in_33, in_32, in_29, 
    in_22;
wire   [9:0] out_0;
wire   [3:0] in_31;
wire   [1:0] in_64;
wire   [1:0] in_62;
wire   [1:0] in_61;
wire   [1:0] in_60;
wire   [1:0] in_54;
wire   [1:0] in_53;
wire   [1:0] in_48;
wire   [1:0] in_47;
wire   [1:0] in_40;
wire   [1:0] in_39;
wire   [1:0] in_36;
wire   [1:0] in_35;
wire   [1:0] in_28;
wire   [1:0] in_27;
wire   [1:0] in_26;
wire   [1:0] in_23;
wire   [5:0] in_21;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_5;
wire   [9:0] in_4;
wire   [9:0] in_3;
wire   [2:0] in_58;
wire   [2:0] in_44;
wire   [2:0] in_34;
wire   [2:0] in_30;
wire   [2:0] in_24;
wire   [2:0] in_2;
wire   [4:0] in_59;
wire   [4:0] in_57;
wire   [4:0] in_56;
wire   [4:0] in_55;
wire   [4:0] in_52;
wire   [4:0] in_49;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_25;
wire   [4:0] in_20;
wire   [4:0] in_7;
wire   [4:0] in_6;
wire   [4:0] in_1;
wire   [4:0] in_0;
  AO21X1 g7007(.Y(out_0[8]), .A0(n_170), .A1(n_213), .B0(out_0[9]));
  NOR2X1 g7008(.Y(out_0[9]), .A(n_170), .B(n_213));
  ADDFX1 g7009(.CO(n_213), .S(out_0[7]), .A(n_171), .B(n_194), .CI(n_210));
  ADDFX1 g7010(.CO(n_210), .S(out_0[6]), .A(n_198), .B(n_195), .CI(n_208));
  ADDFX1 g7011(.CO(n_208), .S(out_0[5]), .A(n_202), .B(n_199), .CI(n_206));
  ADDFX1 g7012(.CO(n_206), .S(out_0[4]), .A(n_200), .B(n_203), .CI(n_204));
  ADDFX1 g7013(.CO(n_204), .S(out_0[3]), .A(n_186), .B(n_196), .CI(n_201));
  ADDFX1 g7014(.CO(n_202), .S(n_203), .A(n_185), .B(n_190), .CI(n_193));
  ADDFX1 g7015(.CO(n_200), .S(n_201), .A(n_191), .B(n_178), .CI(n_183));
  ADDFX1 g7016(.CO(n_198), .S(n_199), .A(n_184), .B(n_189), .CI(n_192));
  ADDFX1 g7017(.CO(n_196), .S(out_0[2]), .A(n_180), .B(n_187), .CI(n_179));
  ADDFX1 g7018(.CO(n_194), .S(n_195), .A(n_161), .B(in_3[6]), .CI(n_188));
  ADDFX1 g7019(.CO(n_192), .S(n_193), .A(n_176), .B(in_3[4]), .CI(n_182));
  ADDFX1 g7020(.CO(n_190), .S(n_191), .A(n_157), .B(n_177), .CI(n_172));
  ADDFX1 g7021(.CO(n_188), .S(n_189), .A(n_174), .B(n_147), .CI(in_3[5]));
  ADDFX1 g7022(.CO(n_186), .S(n_187), .A(n_173), .B(n_168), .CI(n_152));
  ADDFX1 g7023(.CO(n_184), .S(n_185), .A(n_166), .B(n_164), .CI(n_175));
  ADDFX1 g7024(.CO(n_182), .S(n_183), .A(n_159), .B(n_167), .CI(in_3[3]));
  ADDFX1 g7025(.CO(n_180), .S(out_0[1]), .A(n_154), .B(n_169), .CI(n_153));
  ADDFX1 g7026(.CO(n_178), .S(n_179), .A(n_163), .B(n_158), .CI(in_3[2]));
  ADDFX1 g7027(.CO(n_176), .S(n_177), .A(n_162), .B(n_138), .CI(n_165));
  ADDFX1 g7028(.CO(n_174), .S(n_175), .A(n_137), .B(n_150), .CI(in_4[4]));
  ADDFX1 g7029(.CO(n_172), .S(n_173), .A(n_160), .B(n_148), .CI(n_139));
  XNOR2X1 g7030(.Y(n_171), .A(n_156), .B(in_3[7]));
  NOR2BX1 g7031(.Y(n_170), .AN(n_156), .B(in_3[7]));
  ADDFX1 g7032(.CO(n_168), .S(n_169), .A(n_149), .B(n_145), .CI(n_135));
  ADDFX1 g7033(.CO(n_166), .S(n_167), .A(n_122), .B(n_133), .CI(n_151));
  ADDFX1 g7034(.CO(n_164), .S(n_165), .A(n_142), .B(n_120), .CI(in_4[3]));
  ADDFX1 g7035(.CO(n_162), .S(n_163), .A(n_143), .B(n_141), .CI(n_131));
  XNOR2X1 g7036(.Y(n_161), .A(in_4[6]), .B(n_146));
  ADDFX1 g7037(.CO(n_159), .S(n_160), .A(n_129), .B(n_124), .CI(n_134));
  ADDFX1 g7038(.CO(n_157), .S(n_158), .A(n_123), .B(n_144), .CI(n_118));
  NOR2BX1 g7039(.Y(n_156), .AN(n_146), .B(in_4[6]));
  ADDFX1 g7040(.CO(n_154), .S(out_0[0]), .A(n_127), .B(n_91), .CI(n_136));
  ADDFX1 g7041(.CO(n_152), .S(n_153), .A(n_130), .B(n_119), .CI(in_3[1]));
  ADDFX1 g7042(.CO(n_150), .S(n_151), .A(n_104), .B(n_80), .CI(n_140));
  ADDFX1 g7043(.CO(n_148), .S(n_149), .A(n_125), .B(n_132), .CI(n_126));
  XNOR2X1 g7044(.Y(n_147), .A(n_128), .B(in_4[5]));
  NOR2BX1 g7045(.Y(n_146), .AN(in_4[5]), .B(n_128));
  ADDFX1 g7046(.CO(n_144), .S(n_145), .A(n_113), .B(n_117), .CI(n_90));
  ADDFX1 g7047(.CO(n_142), .S(n_143), .A(n_44), .B(n_114), .CI(n_84));
  ADDFX1 g7048(.CO(n_140), .S(n_141), .A(n_86), .B(n_108), .CI(n_94));
  ADDFX1 g7049(.CO(n_138), .S(n_139), .A(n_82), .B(n_116), .CI(in_4[2]));
  AO21X1 g7050(.Y(n_137), .A0(n_105), .A1(n_121), .B0(n_128));
  ADDFX1 g7051(.CO(n_135), .S(n_136), .A(n_111), .B(n_93), .CI(in_3[0]));
  ADDFX1 g7052(.CO(n_133), .S(n_134), .A(n_89), .B(n_107), .CI(n_81));
  ADDFX1 g7053(.CO(n_131), .S(n_132), .A(n_87), .B(n_109), .CI(n_102));
  ADDFX1 g7054(.CO(n_129), .S(n_130), .A(n_78), .B(n_92), .CI(n_110));
  NOR2X1 g7055(.Y(n_128), .A(n_105), .B(n_121));
  ADDFX1 g7056(.CO(n_126), .S(n_127), .A(n_79), .B(n_101), .CI(n_103));
  ADDFX1 g7057(.CO(n_124), .S(n_125), .A(n_95), .B(n_85), .CI(n_100));
  ADDFX1 g7058(.CO(n_122), .S(n_123), .A(n_99), .B(n_112), .CI(n_96));
  ADDFX1 g7059(.CO(n_121), .S(n_120), .A(n_98), .B(n_106), .CI(n_88));
  ADDFX1 g7060(.CO(n_118), .S(n_119), .A(n_97), .B(n_83), .CI(in_4[1]));
  ADDFX1 g7061(.CO(n_116), .S(n_117), .A(n_45), .B(n_28), .CI(n_115));
  ADDFX1 g7062(.CO(n_114), .S(n_115), .A(n_70), .B(n_18), .CI(n_50));
  ADDFX1 g7063(.CO(n_112), .S(n_113), .A(n_61), .B(n_75), .CI(n_77));
  ADDFX1 g7064(.CO(n_110), .S(n_111), .A(n_71), .B(n_41), .CI(n_33));
  ADDFX1 g7065(.CO(n_108), .S(n_109), .A(n_52), .B(n_68), .CI(n_32));
  ADDFX1 g7066(.CO(n_106), .S(n_107), .A(n_56), .B(n_24), .CI(n_76));
  ADDFX1 g7067(.CO(n_105), .S(n_104), .A(n_22), .B(n_26), .CI(n_66));
  ADDFX1 g7068(.CO(n_102), .S(n_103), .A(n_65), .B(n_63), .CI(n_43));
  ADDFX1 g7069(.CO(n_100), .S(n_101), .A(n_51), .B(n_35), .CI(n_69));
  ADDFX1 g7070(.CO(n_98), .S(n_99), .A(n_23), .B(n_46), .CI(n_72));
  ADDFX1 g7071(.CO(n_96), .S(n_97), .A(n_47), .B(n_55), .CI(n_73));
  ADDFX1 g7072(.CO(n_94), .S(n_95), .A(n_64), .B(n_58), .CI(n_62));
  ADDFX1 g7073(.CO(n_92), .S(n_93), .A(n_53), .B(n_49), .CI(n_31));
  ADDFX1 g7074(.CO(n_90), .S(n_91), .A(n_59), .B(n_29), .CI(in_4[0]));
  ADDFX1 g7075(.CO(n_88), .S(n_89), .A(n_74), .B(n_60), .CI(n_54));
  ADDFX1 g7076(.CO(n_86), .S(n_87), .A(n_48), .B(n_36), .CI(n_42));
  ADDFX1 g7077(.CO(n_84), .S(n_85), .A(n_40), .B(n_30), .CI(n_34));
  ADDFX1 g7078(.CO(n_82), .S(n_83), .A(n_25), .B(n_57), .CI(n_39));
  ADDFX1 g7079(.CO(n_80), .S(n_81), .A(n_27), .B(n_38), .CI(n_67));
  ADDFX1 g7080(.CO(n_78), .S(n_79), .A(in_13[0]), .B(in_10[0]), .CI(n_37));
  ADDFX1 g7081(.CO(n_76), .S(n_77), .A(in_27[0]), .B(in_61[0]), .CI(in_36[0]));
  ADDFX1 g7082(.CO(n_74), .S(n_75), .A(in_28[1]), .B(in_30[0]), .CI(in_60[0]));
  ADDFX1 g7083(.CO(n_72), .S(n_73), .A(in_24[0]), .B(n_10), .CI(n_21));
  ADDFX1 g7084(.CO(n_70), .S(n_71), .A(in_41), .B(in_44[0]), .CI(in_63));
  ADDFX1 g7085(.CO(n_68), .S(n_69), .A(in_51), .B(in_53[0]), .CI(in_54[0]));
  ADDFX1 g7086(.CO(n_66), .S(n_67), .A(n_8), .B(in_64[1]), .CI(n_16));
  ADDFX1 g7087(.CO(n_64), .S(n_65), .A(in_37), .B(n_11), .CI(n_15));
  ADDFX1 g7088(.CO(n_62), .S(n_63), .A(in_24[0]), .B(n_14), .CI(in_40[0]));
  ADDFX1 g7089(.CO(n_60), .S(n_61), .A(in_9[1]), .B(in_34[0]), .CI(in_44[0]));
  ADDFX1 g7090(.CO(n_58), .S(n_59), .A(in_32), .B(in_15[0]), .CI(in_42));
  ADDFX1 g7091(.CO(n_56), .S(n_57), .A(in_23[1]), .B(in_26[1]), .CI(in_58[1]));
  ADDFX1 g7092(.CO(n_54), .S(n_55), .A(in_39[0]), .B(in_2[1]), .CI(in_62[0]));
  ADDFX1 g7093(.CO(n_52), .S(n_53), .A(in_8[0]), .B(in_50), .CI(in_22));
  ADDFX1 g7094(.CO(n_50), .S(n_51), .A(in_34[0]), .B(in_38), .CI(n_20));
  ADDFX1 g7095(.CO(n_48), .S(n_49), .A(in_35[0]), .B(n_17), .CI(in_62[0]));
  ADDFX1 g7096(.CO(n_46), .S(n_47), .A(in_40[0]), .B(n_3), .CI(n_19));
  ADDFX1 g7097(.CO(n_44), .S(n_45), .A(in_39[0]), .B(n_2), .CI(n_4));
  ADDFX1 g7098(.CO(n_42), .S(n_43), .A(in_18[0]), .B(in_30[0]), .CI(in_47[0]));
  ADDFX1 g7099(.CO(n_40), .S(n_41), .A(in_43), .B(n_13), .CI(in_65));
  ADDFX1 g7100(.CO(n_38), .S(n_39), .A(n_7), .B(n_12), .CI(in_13[1]));
  ADDFX1 g7101(.CO(n_36), .S(n_37), .A(in_14[0]), .B(in_48[0]), .CI(in_20[0]));
  ADDFX1 g7102(.CO(n_34), .S(n_35), .A(in_36[0]), .B(in_61[0]), .CI(n_5));
  ADDFX1 g7103(.CO(n_32), .S(n_33), .A(in_29), .B(in_33), .CI(in_60[0]));
  ADDFX1 g7104(.CO(n_30), .S(n_31), .A(in_7[0]), .B(in_27[0]), .CI(in_49[0]));
  ADDFX1 g7105(.CO(n_28), .S(n_29), .A(n_0), .B(in_11[0]), .CI(in_19[0]));
  ADDFX1 g7106(.CO(n_26), .S(n_27), .A(in_16[2]), .B(n_1), .CI(n_9));
  ADDFX1 g7107(.CO(n_24), .S(n_25), .A(in_17[1]), .B(in_12[1]), .CI(n_6));
  XNOR2X1 g7108(.Y(n_23), .A(in_31[2]), .B(in_49[0]));
  NOR2BX1 g7109(.Y(n_22), .AN(in_31[2]), .B(in_49[0]));
  INVX1 g7110(.Y(n_21), .A(in_59[1]));
  INVX1 g7111(.Y(n_20), .A(in_52[0]));
  INVX1 g7112(.Y(n_19), .A(in_55[1]));
  INVX1 g7113(.Y(n_18), .A(in_11[1]));
  INVX1 g7114(.Y(n_17), .A(in_45[0]));
  INVX1 g7115(.Y(n_16), .A(in_13[2]));
  INVX1 g7116(.Y(n_15), .A(in_5[0]));
  INVX1 g7117(.Y(n_14), .A(in_0[0]));
  INVX1 g7118(.Y(n_13), .A(in_46[0]));
  INVX1 g7119(.Y(n_12), .A(in_19[1]));
  INVX1 g7120(.Y(n_11), .A(in_1[0]));
  INVX1 g7121(.Y(n_10), .A(in_6[1]));
  INVX1 g7122(.Y(n_9), .A(in_20[0]));
  INVX1 g7123(.Y(n_8), .A(in_15[0]));
  INVX1 g7124(.Y(n_7), .A(in_57[1]));
  INVX1 g7125(.Y(n_6), .A(in_56[1]));
  INVX1 g7126(.Y(n_5), .A(in_21[0]));
  INVX1 g7127(.Y(n_4), .A(in_10[1]));
  INVX1 g7128(.Y(n_3), .A(in_25[1]));
  INVX1 g7129(.Y(n_2), .A(in_64[1]));
  INVX1 g7130(.Y(n_1), .A(in_7[0]));
  INVX1 g7131(.Y(n_0), .A(in_39[0]));
endmodule

module WALLACE_CSA_DUMMY_OP157_group_109824(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, out_0);
input  in_29, in_30, in_39, in_40;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [2:0] in_19;
input   [4:0] in_20;
input   [2:0] in_21;
input   [2:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [1:0] in_28;
input   [2:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
output  [9:0] out_0;
wire  n_111, n_108, n_106, n_105, n_104, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_40, in_39, 
    in_30, in_29;
wire   [9:0] out_0;
wire   [1:0] in_28;
wire   [2:0] in_31;
wire   [2:0] in_22;
wire   [2:0] in_21;
wire   [2:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_20;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  OA21X1 g3106(.Y(out_0[5]), .A0(n_98), .A1(n_111), .B0(out_0[9]));
  NAND2X1 g3107(.Y(out_0[9]), .A(n_98), .B(n_111));
  ADDFX1 g3108(.CO(n_111), .S(out_0[4]), .A(n_99), .B(n_104), .CI(n_108));
  ADDFX1 g3109(.CO(n_108), .S(out_0[3]), .A(n_100), .B(n_105), .CI(n_106));
  ADDFX1 g3110(.CO(n_106), .S(out_0[2]), .A(n_92), .B(n_101), .CI(n_102));
  ADDFX1 g3111(.CO(n_104), .S(n_105), .A(n_84), .B(n_94), .CI(n_96));
  ADDFX1 g3112(.CO(n_102), .S(out_0[1]), .A(n_87), .B(n_90), .CI(n_93));
  ADDFX1 g3113(.CO(n_100), .S(n_101), .A(n_86), .B(n_85), .CI(n_95));
  OAI2BB1X1 g3114(.Y(n_99), .A0N(n_72), .A1N(n_97), .B0(n_98));
  OR2X1 g3115(.Y(n_98), .A(n_72), .B(n_97));
  ADDFX1 g3116(.CO(n_97), .S(n_96), .A(n_75), .B(n_76), .CI(n_88));
  ADDFX1 g3117(.CO(n_94), .S(n_95), .A(n_77), .B(n_89), .CI(n_82));
  ADDFX1 g3118(.CO(n_92), .S(n_93), .A(n_78), .B(n_83), .CI(n_81));
  ADDFX1 g3119(.CO(n_90), .S(out_0[0]), .A(n_69), .B(n_57), .CI(n_79));
  ADDFX1 g3120(.CO(n_88), .S(n_89), .A(n_62), .B(n_73), .CI(n_60));
  ADDFX1 g3121(.CO(n_86), .S(n_87), .A(n_74), .B(n_65), .CI(n_61));
  ADDFX1 g3122(.CO(n_84), .S(n_85), .A(n_64), .B(n_70), .CI(n_80));
  ADDFX1 g3123(.CO(n_82), .S(n_83), .A(n_37), .B(n_63), .CI(n_66));
  ADDFX1 g3124(.CO(n_80), .S(n_81), .A(n_68), .B(n_59), .CI(n_56));
  ADDFX1 g3125(.CO(n_78), .S(n_79), .A(n_33), .B(n_38), .CI(n_67));
  ADDFX1 g3126(.CO(n_76), .S(n_77), .A(n_41), .B(n_55), .CI(n_58));
  OAI2BB1X1 g3127(.Y(n_75), .A0N(n_52), .A1N(n_71), .B0(n_72));
  ADDFX1 g3128(.CO(n_73), .S(n_74), .A(n_4), .B(n_53), .CI(n_28));
  OR2X1 g3129(.Y(n_72), .A(n_52), .B(n_71));
  ADDFX1 g3130(.CO(n_71), .S(n_70), .A(n_22), .B(n_39), .CI(n_26));
  ADDFX1 g3131(.CO(n_68), .S(n_69), .A(in_12[0]), .B(n_31), .CI(n_35));
  ADDFX1 g3132(.CO(n_66), .S(n_67), .A(n_48), .B(n_46), .CI(n_54));
  ADDFX1 g3133(.CO(n_64), .S(n_65), .A(n_23), .B(n_47), .CI(n_36));
  ADDFX1 g3134(.CO(n_62), .S(n_63), .A(n_34), .B(n_32), .CI(n_30));
  ADDFX1 g3135(.CO(n_60), .S(n_61), .A(n_40), .B(n_27), .CI(n_42));
  ADDFX1 g3136(.CO(n_58), .S(n_59), .A(n_50), .B(n_45), .CI(n_24));
  ADDFX1 g3137(.CO(n_56), .S(n_57), .A(n_51), .B(n_29), .CI(n_25));
  OAI2BB1X1 g3138(.Y(n_55), .A0N(n_13), .A1N(n_49), .B0(n_52));
  ADDFX1 g3139(.CO(n_53), .S(n_54), .A(in_30), .B(n_18), .CI(n_6));
  OR2X1 g3140(.Y(n_52), .A(n_13), .B(n_49));
  INVX1 g3141(.Y(n_51), .A(n_44));
  INVX1 g3142(.Y(n_50), .A(n_43));
  ADDFX1 g3143(.CO(n_47), .S(n_48), .A(in_8[0]), .B(in_5[0]), .CI(in_22[0]));
  ADDFX1 g3144(.CO(n_45), .S(n_46), .A(in_28[0]), .B(n_16), .CI(in_39));
  ADDFX1 g3145(.CO(n_43), .S(n_44), .A(in_1[0]), .B(in_0[0]), .CI(in_27[0]));
  ADDFX1 g3146(.CO(n_41), .S(n_42), .A(in_16[1]), .B(in_31[1]), .CI(n_15));
  ADDFX1 g3147(.CO(n_39), .S(n_40), .A(in_8[1]), .B(in_19[1]), .CI(in_21[1]));
  ADDFX1 g3148(.CO(n_37), .S(n_38), .A(n_14), .B(in_29), .CI(in_3[0]));
  ADDFX1 g3149(.CO(n_49), .S(n_36), .A(in_10[1]), .B(n_17), .CI(n_19));
  ADDFX1 g3150(.CO(n_34), .S(n_35), .A(n_1), .B(n_2), .CI(in_40));
  ADDFX1 g3151(.CO(n_32), .S(n_33), .A(in_14[0]), .B(n_7), .CI(n_12));
  ADDFX1 g3152(.CO(n_30), .S(n_31), .A(in_7[0]), .B(n_8), .CI(n_11));
  ADDFX1 g3153(.CO(n_28), .S(n_29), .A(in_4[0]), .B(n_5), .CI(n_20));
  ADDFX1 g3154(.CO(n_26), .S(n_27), .A(in_22[0]), .B(n_3), .CI(n_10));
  ADDFX1 g3155(.CO(n_24), .S(n_25), .A(in_6[0]), .B(in_13[0]), .CI(n_9));
  OAI2BB1X1 g3156(.Y(n_23), .A0N(in_5[1]), .A1N(n_21), .B0(n_22));
  OR2X1 g3157(.Y(n_22), .A(in_5[1]), .B(n_21));
  INVX1 g3158(.Y(n_21), .A(in_25[1]));
  INVX1 g3159(.Y(n_20), .A(in_32[0]));
  INVX1 g3160(.Y(n_19), .A(in_34[1]));
  INVX1 g3161(.Y(n_18), .A(in_33[0]));
  INVX1 g3162(.Y(n_17), .A(in_23[1]));
  INVX1 g3163(.Y(n_16), .A(in_2[0]));
  INVX1 g3164(.Y(n_15), .A(in_12[1]));
  INVX1 g3165(.Y(n_14), .A(in_18[0]));
  INVX1 g3166(.Y(n_13), .A(in_6[0]));
  INVX1 g3167(.Y(n_12), .A(in_24[0]));
  INVX1 g3168(.Y(n_11), .A(in_36[0]));
  INVX1 g3169(.Y(n_10), .A(in_37[1]));
  INVX1 g3170(.Y(n_9), .A(in_38[0]));
  INVX1 g3171(.Y(n_8), .A(in_17[0]));
  INVX1 g3172(.Y(n_7), .A(in_15[0]));
  INVX1 g3173(.Y(n_6), .A(in_9[0]));
  INVX1 g3174(.Y(n_5), .A(in_26[0]));
  INVX1 g3175(.Y(n_4), .A(in_3[1]));
  INVX1 g3176(.Y(n_3), .A(in_20[1]));
  INVX1 g3177(.Y(n_2), .A(in_35[0]));
  INVX1 g3178(.Y(n_1), .A(in_11[0]));
endmodule

module WALLACE_CSA_DUMMY_OP162_group_109829_6307(in_0, in_1, in_2, in_3, in_4, 
    in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, in_39, in_40, in_41, out_0);
input  in_24, in_25, in_31, in_32, in_35, in_41;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [2:0] in_4;
input   [4:0] in_5;
input   [9:0] in_6;
input   [6:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [2:0] in_26;
input   [4:0] in_27;
input   [2:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_33;
input   [2:0] in_34;
input   [1:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
output  [9:0] out_0;
wire  n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, 
    n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, 
    n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, 
    n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, 
    n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, 
    n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, 
    n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_39, n_37, n_35, 
    n_33, n_31, n_29, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1, in_41, in_35, in_32, in_31, in_25, in_24;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_36;
wire   [1:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_7;
wire   [9:0] in_6;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_33;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_23;
wire   [4:0] in_5;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_34;
wire   [2:0] in_30;
wire   [2:0] in_28;
wire   [2:0] in_26;
wire   [2:0] in_4;
wire   [2:0] in_3;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_113), .S(n_112), .A(in_18[0]), .B(n_7), .CI(
    in_13[0]));
  ADDFX1 cdnfadd_000_1(.CO(n_111), .S(n_110), .A(n_19), .B(n_21), .CI(in_25));
  ADDFX1 cdnfadd_000_2(.CO(n_109), .S(n_108), .A(in_39[0]), .B(in_41), .CI(in_24));
  ADDFX1 cdnfadd_000_3(.CO(n_107), .S(n_106), .A(n_4), .B(in_9[0]), .CI(in_28[0]));
  ADDFX1 cdnfadd_000_4(.CO(n_105), .S(n_104), .A(in_32), .B(in_19[0]), .CI(
    in_30[0]));
  ADDFX1 cdnfadd_000_5(.CO(n_103), .S(n_102), .A(in_22[0]), .B(n_16), .CI(n_6));
  ADDFX1 cdnfadd_000_6(.CO(n_101), .S(n_100), .A(n_8), .B(in_11[0]), .CI(in_31));
  ADDFX1 cdnfadd_000_7(.CO(n_99), .S(n_98), .A(in_10[0]), .B(n_24), .CI(in_14[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_76), .S(n_116), .A(n_110), .B(n_112), .CI(n_100));
  ADDFX1 cdnfadd_000_9(.CO(n_75), .S(n_124), .A(n_104), .B(n_106), .CI(n_102));
  ADDFX1 cdnfadd_000_10(.CO(n_74), .S(n_117), .A(n_108), .B(n_98), .CI(in_6[0]));
  ADDFX1 cdnfadd_001_0(.CO(n_97), .S(n_96), .A(in_28[0]), .B(n_9), .CI(n_17));
  ADDFX1 cdnfadd_001_1(.CO(n_95), .S(n_94), .A(n_20), .B(n_14), .CI(in_7[1]));
  ADDFX1 cdnfadd_001_2(.CO(n_93), .S(n_92), .A(in_30[0]), .B(in_40[1]), .CI(n_15));
  ADDFX1 cdnfadd_001_3(.CO(n_91), .S(n_90), .A(n_10), .B(in_36[1]), .CI(in_34[1]));
  ADDFX1 cdnfadd_001_4(.CO(n_89), .S(n_88), .A(n_5), .B(in_0[1]), .CI(in_4[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_87), .S(n_86), .A(in_26[1]), .B(in_14[1]), .CI(n_2));
  ADDFX1 cdnfadd_001_6(.CO(n_73), .S(n_72), .A(in_18[1]), .B(n_23), .CI(n_101));
  ADDFX1 cdnfadd_001_7(.CO(n_71), .S(n_70), .A(n_107), .B(n_111), .CI(n_103));
  ADDFX1 cdnfadd_001_8(.CO(n_69), .S(n_68), .A(n_113), .B(n_105), .CI(n_109));
  ADDFX1 cdnfadd_001_9(.CO(n_67), .S(n_66), .A(n_94), .B(n_88), .CI(n_96));
  ADDFX1 cdnfadd_001_10(.CO(n_65), .S(n_64), .A(n_92), .B(n_90), .CI(n_86));
  ADDFX1 cdnfadd_001_11(.CO(n_57), .S(n_56), .A(n_99), .B(n_72), .CI(n_75));
  ADDFX1 cdnfadd_001_12(.CO(n_55), .S(n_54), .A(n_76), .B(n_68), .CI(n_70));
  ADDFX1 cdnfadd_001_13(.CO(n_53), .S(n_125), .A(n_64), .B(n_66), .CI(n_74));
  ADDFX1 cdnfadd_001_14(.CO(n_44), .S(n_118), .A(n_56), .B(in_6[1]), .CI(n_54));
  ADDFX1 cdnfadd_002_0(.CO(n_85), .S(n_84), .A(n_12), .B(n_1), .CI(n_11));
  ADDFX1 cdnfadd_002_1(.CO(n_83), .S(n_82), .A(n_18), .B(n_25), .CI(in_3[1]));
  ADDFX1 cdnfadd_002_2(.CO(n_63), .S(n_62), .A(n_97), .B(n_95), .CI(n_91));
  ADDFX1 cdnfadd_002_3(.CO(n_61), .S(n_60), .A(n_93), .B(n_89), .CI(n_84));
  ADDFX1 cdnfadd_002_4(.CO(n_52), .S(n_51), .A(n_87), .B(n_71), .CI(n_69));
  ADDFX1 cdnfadd_002_5(.CO(n_50), .S(n_49), .A(n_82), .B(n_73), .CI(n_67));
  ADDFX1 cdnfadd_002_6(.CO(n_48), .S(n_47), .A(n_62), .B(n_60), .CI(n_65));
  ADDFX1 cdnfadd_002_7(.CO(n_43), .S(n_42), .A(n_55), .B(n_57), .CI(n_49));
  ADDFX1 cdnfadd_002_8(.CO(n_81), .S(n_126), .A(n_51), .B(n_47), .CI(in_6[2]));
  ADDFX1 cdnfadd_002_9(.CO(n_127), .S(n_119), .A(n_53), .B(n_42), .CI(n_44));
  ADDFX1 cdnfadd_003_0(.CO(n_59), .S(n_58), .A(n_22), .B(n_85), .CI(n_83));
  ADDFX1 cdnfadd_003_1(.CO(n_46), .S(n_45), .A(n_63), .B(n_61), .CI(n_58));
  ADDFX1 cdnfadd_003_2(.CO(n_115), .S(n_114), .A(n_52), .B(n_50), .CI(n_48));
  ADDFX1 cdnfadd_003_3(.CO(n_80), .S(n_79), .A(n_45), .B(in_6[3]), .CI(n_43));
  ADDFX1 cdnfadd_003_4(.CO(n_128), .S(n_120), .A(n_114), .B(n_81), .CI(n_79));
  ADDFX1 cdnfadd_004_0(.CO(n_77), .S(n_78), .A(n_26), .B(n_46), .CI(in_6[4]));
  ADDFX1 cdnfadd_004_1(.CO(n_129), .S(n_121), .A(n_115), .B(n_78), .CI(n_80));
  ADDFX1 cdnfadd_005_0(.CO(n_123), .S(n_122), .A(n_59), .B(in_6[5]), .CI(n_77));
  INVX1 g308(.Y(out_0[9]), .A(n_39));
  ADDFX1 g309(.CO(n_39), .S(out_0[6]), .A(n_13), .B(n_123), .CI(n_37));
  ADDFX1 g310(.CO(n_37), .S(out_0[5]), .A(n_122), .B(n_129), .CI(n_35));
  ADDFX1 g311(.CO(n_35), .S(out_0[4]), .A(n_128), .B(n_121), .CI(n_33));
  ADDFX1 g312(.CO(n_33), .S(out_0[3]), .A(n_127), .B(n_31), .CI(n_120));
  ADDFX1 g313(.CO(n_31), .S(out_0[2]), .A(n_126), .B(n_29), .CI(n_119));
  ADDFX1 g314(.CO(n_29), .S(out_0[1]), .A(n_27), .B(n_125), .CI(n_118));
  ADDFX1 g315(.CO(n_27), .S(out_0[0]), .A(n_116), .B(n_124), .CI(n_117));
  INVX1 g316(.Y(n_26), .A(n_59));
  AOI21X1 g317(.Y(n_25), .A0(in_14[2]), .A1(in_37[2]), .B0(n_22));
  AOI21X1 g318(.Y(n_24), .A0(in_33[0]), .A1(n_3), .B0(n_23));
  NOR2X1 g319(.Y(n_23), .A(in_33[0]), .B(n_3));
  NOR2X1 g320(.Y(n_22), .A(in_37[2]), .B(in_14[2]));
  INVX1 g321(.Y(n_21), .A(in_8[0]));
  INVX1 g322(.Y(n_20), .A(in_15[1]));
  INVX1 g323(.Y(n_19), .A(in_5[0]));
  INVX1 g324(.Y(n_18), .A(in_18[2]));
  INVX1 g325(.Y(n_17), .A(in_27[1]));
  INVX1 g326(.Y(n_16), .A(in_38[0]));
  INVX1 g327(.Y(n_15), .A(in_29[1]));
  INVX1 g328(.Y(n_14), .A(in_12[1]));
  INVX1 g329(.Y(n_13), .A(in_6[6]));
  INVX1 g330(.Y(n_12), .A(in_13[0]));
  INVX1 g331(.Y(n_11), .A(in_10[0]));
  INVX1 g332(.Y(n_10), .A(in_2[1]));
  INVX1 g333(.Y(n_9), .A(in_23[1]));
  INVX1 g334(.Y(n_8), .A(in_17[0]));
  INVX1 g335(.Y(n_7), .A(in_20[0]));
  INVX1 g336(.Y(n_6), .A(in_16[0]));
  INVX1 g337(.Y(n_5), .A(in_21[1]));
  INVX1 g338(.Y(n_4), .A(in_1[0]));
  INVX1 g339(.Y(n_3), .A(in_35));
  INVX1 g340(.Y(n_2), .A(in_3[1]));
  INVX1 g341(.Y(n_1), .A(in_39[0]));
endmodule

module WALLACE_CSA_DUMMY_OP162_group_109829(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, out_0);
input  in_31, in_34, in_35, in_41;
input   [2:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [4:0] in_8;
input   [4:0] in_9;
input   [1:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [1:0] in_21;
input   [2:0] in_22;
input   [4:0] in_23;
input   [1:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [2:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [2:0] in_32;
input   [4:0] in_33;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [1:0] in_40;
output  [9:0] out_0;
wire  n_133, n_130, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, 
    n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_41, 
    in_35, in_34, in_31;
wire   [9:0] out_0;
wire   [1:0] in_40;
wire   [1:0] in_29;
wire   [1:0] in_27;
wire   [1:0] in_24;
wire   [1:0] in_21;
wire   [1:0] in_10;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_30;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_23;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [4:0] in_9;
wire   [4:0] in_8;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [2:0] in_37;
wire   [2:0] in_32;
wire   [2:0] in_28;
wire   [2:0] in_22;
wire   [2:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  OAI211X1 g3968(.Y(out_0[9]), .A0(n_124), .A1(n_133), .B0(n_107), .C0(n_123));
  XNOR2X1 g3969(.Y(out_0[5]), .A(n_127), .B(n_133));
  ADDFX1 g3970(.CO(n_133), .S(out_0[4]), .A(n_121), .B(n_125), .CI(n_130));
  ADDFX1 g3971(.CO(n_130), .S(out_0[3]), .A(n_119), .B(n_126), .CI(n_128));
  ADDFX1 g3972(.CO(n_128), .S(out_0[2]), .A(n_108), .B(n_117), .CI(n_120));
  NAND2BX1 g3973(.Y(n_127), .AN(n_124), .B(n_123));
  ADDFX1 g3974(.CO(n_125), .S(n_126), .A(n_112), .B(n_115), .CI(n_114));
  NOR2BX1 g3975(.Y(n_124), .AN(n_122), .B(n_110));
  NAND2BX1 g3976(.Y(n_123), .AN(n_122), .B(n_110));
  ADDFX1 g3977(.CO(n_122), .S(n_121), .A(n_111), .B(n_102), .CI(n_113));
  ADDFX1 g3978(.CO(n_119), .S(n_120), .A(n_96), .B(n_105), .CI(n_116));
  ADDFX1 g3979(.CO(n_117), .S(out_0[1]), .A(n_97), .B(n_98), .CI(n_109));
  ADDFX1 g3980(.CO(n_115), .S(n_116), .A(n_93), .B(n_100), .CI(n_91));
  ADDFX1 g3981(.CO(n_113), .S(n_114), .A(n_95), .B(n_90), .CI(n_104));
  ADDFX1 g3982(.CO(n_111), .S(n_112), .A(n_88), .B(n_83), .CI(n_92));
  AOI21X1 g3983(.Y(n_110), .A0(n_49), .A1(n_103), .B0(n_106));
  ADDFX1 g3984(.CO(n_108), .S(n_109), .A(n_70), .B(n_87), .CI(n_101));
  INVX1 g3985(.Y(n_107), .A(n_106));
  NOR2X1 g3986(.Y(n_106), .A(n_49), .B(n_103));
  ADDFX1 g3987(.CO(n_104), .S(n_105), .A(n_79), .B(n_89), .CI(n_86));
  ADDFX1 g3988(.CO(n_103), .S(n_102), .A(n_20), .B(n_82), .CI(n_94));
  ADDFX1 g3989(.CO(n_100), .S(n_101), .A(n_77), .B(n_84), .CI(n_81));
  ADDFX1 g3990(.CO(n_98), .S(out_0[0]), .A(n_85), .B(n_75), .CI(n_71));
  ADDFX1 g3991(.CO(n_96), .S(n_97), .A(n_74), .B(n_69), .CI(n_67));
  ADDFX1 g3992(.CO(n_94), .S(n_95), .A(n_64), .B(n_72), .CI(n_78));
  ADDFX1 g3993(.CO(n_92), .S(n_93), .A(n_60), .B(n_65), .CI(n_76));
  ADDFX1 g3994(.CO(n_90), .S(n_91), .A(n_73), .B(n_68), .CI(n_66));
  ADDFX1 g3995(.CO(n_88), .S(n_89), .A(n_32), .B(n_58), .CI(n_80));
  ADDFX1 g3996(.CO(n_86), .S(n_87), .A(n_42), .B(n_59), .CI(n_61));
  ADDFX1 g3997(.CO(n_84), .S(n_85), .A(n_57), .B(n_23), .CI(n_55));
  ADDFX1 g3998(.CO(n_82), .S(n_83), .A(n_52), .B(n_21), .CI(n_30));
  ADDFX1 g3999(.CO(n_80), .S(n_81), .A(n_54), .B(n_56), .CI(n_22));
  ADDFX1 g4000(.CO(n_78), .S(n_79), .A(n_19), .B(n_53), .CI(n_31));
  ADDFX1 g4001(.CO(n_76), .S(n_77), .A(n_44), .B(n_28), .CI(n_40));
  ADDFX1 g4002(.CO(n_74), .S(n_75), .A(n_29), .B(n_35), .CI(n_41));
  ADDFX1 g4003(.CO(n_72), .S(n_73), .A(n_46), .B(n_26), .CI(n_24));
  ADDFX1 g4004(.CO(n_70), .S(n_71), .A(n_45), .B(n_43), .CI(n_37));
  ADDFX1 g4005(.CO(n_68), .S(n_69), .A(n_27), .B(n_47), .CI(n_25));
  ADDFX1 g4006(.CO(n_66), .S(n_67), .A(n_48), .B(n_36), .CI(n_33));
  INVX1 g4007(.Y(n_65), .A(n_63));
  INVX1 g4008(.Y(n_64), .A(n_62));
  ADDFX1 g4009(.CO(n_62), .S(n_63), .A(n_17), .B(in_7[2]), .CI(n_38));
  ADDFX1 g4010(.CO(n_60), .S(n_61), .A(in_11[0]), .B(in_6[1]), .CI(n_34));
  ADDFX1 g4011(.CO(n_58), .S(n_59), .A(n_12), .B(n_18), .CI(in_7[1]));
  ADDFX1 g4012(.CO(n_56), .S(n_57), .A(in_10[0]), .B(in_35), .CI(n_3));
  ADDFX1 g4013(.CO(n_54), .S(n_55), .A(in_2[0]), .B(in_27[0]), .CI(in_4[0]));
  INVX1 g4014(.Y(n_53), .A(n_51));
  INVX1 g4015(.Y(n_52), .A(n_50));
  ADDFX1 g4016(.CO(n_50), .S(n_51), .A(in_9[0]), .B(in_20[2]), .CI(in_30[0]));
  INVX1 g4017(.Y(n_49), .A(n_20));
  INVX1 g4018(.Y(n_48), .A(n_39));
  ADDFX1 g4019(.CO(n_46), .S(n_47), .A(in_17[0]), .B(n_4), .CI(n_7));
  ADDFX1 g4020(.CO(n_44), .S(n_45), .A(in_31), .B(n_5), .CI(n_6));
  ADDFX1 g4021(.CO(n_42), .S(n_43), .A(in_23[0]), .B(in_12[0]), .CI(in_16[0]));
  ADDFX1 g4022(.CO(n_40), .S(n_41), .A(in_7[0]), .B(n_10), .CI(in_17[0]));
  ADDFX1 g4023(.CO(n_38), .S(n_39), .A(in_3[1]), .B(in_8[1]), .CI(in_13[1]));
  ADDFX1 g4024(.CO(n_36), .S(n_37), .A(n_9), .B(in_5[0]), .CI(in_14[0]));
  ADDFX1 g4025(.CO(n_34), .S(n_35), .A(in_6[0]), .B(in_34), .CI(in_41));
  ADDFX1 g4026(.CO(n_32), .S(n_33), .A(in_5[1]), .B(n_2), .CI(n_14));
  ADDFX1 g4027(.CO(n_30), .S(n_31), .A(in_32[2]), .B(n_9), .CI(n_13));
  ADDFX1 g4028(.CO(n_28), .S(n_29), .A(in_21[0]), .B(in_29[0]), .CI(in_30[0]));
  ADDFX1 g4029(.CO(n_26), .S(n_27), .A(in_22[1]), .B(n_11), .CI(n_15));
  ADDFX1 g4030(.CO(n_24), .S(n_25), .A(in_28[1]), .B(in_0[1]), .CI(in_40[1]));
  ADDFX1 g4031(.CO(n_22), .S(n_23), .A(in_9[0]), .B(in_24[0]), .CI(n_8));
  OAI2BB1X1 g4032(.Y(n_21), .A0N(n_1), .A1N(n_16), .B0(n_49));
  NOR2X1 g4034(.Y(n_20), .A(n_1), .B(n_16));
  OAI21X1 g4035(.Y(n_19), .A0(in_2[0]), .A1(in_23[0]), .B0(n_16));
  XNOR2X1 g4036(.Y(n_18), .A(in_25[1]), .B(in_37[1]));
  NAND2BX1 g4037(.Y(n_17), .AN(in_25[1]), .B(in_37[1]));
  NAND2X1 g4038(.Y(n_16), .A(in_23[0]), .B(in_2[0]));
  INVX1 g4039(.Y(n_15), .A(in_38[1]));
  INVX1 g4040(.Y(n_14), .A(in_14[1]));
  INVX1 g4041(.Y(n_13), .A(in_6[2]));
  INVX1 g4042(.Y(n_12), .A(in_16[1]));
  INVX1 g4043(.Y(n_11), .A(in_18[1]));
  INVX1 g4044(.Y(n_10), .A(in_1[0]));
  INVX1 g4045(.Y(n_9), .A(in_11[0]));
  INVX1 g4046(.Y(n_8), .A(in_39[0]));
  INVX1 g4047(.Y(n_7), .A(in_33[1]));
  INVX1 g4048(.Y(n_6), .A(in_36[0]));
  INVX1 g4049(.Y(n_5), .A(in_19[0]));
  INVX1 g4050(.Y(n_4), .A(in_15[1]));
  INVX1 g4051(.Y(n_3), .A(in_26[0]));
  INVX1 g4052(.Y(n_2), .A(in_12[1]));
  INVX1 g4053(.Y(n_1), .A(in_17[0]));
endmodule

module WALLACE_CSA_DUMMY_OP258_group_359288(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, out_0);
input  in_19, in_27, in_35;
input   [4:0] in_0;
input   [4:0] in_1;
input   [1:0] in_2;
input   [1:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [1:0] in_18;
input   [4:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [1:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [1:0] in_32;
input   [4:0] in_33;
input   [1:0] in_34;
input   [1:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [2:0] in_43;
input   [2:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
output  [9:0] out_0;
wire  n_131, n_129, n_127, n_125, n_124, n_123, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_0, in_35, in_27, 
    in_19;
wire   [9:0] out_0;
wire   [2:0] in_44;
wire   [2:0] in_43;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [1:0] in_36;
wire   [1:0] in_34;
wire   [1:0] in_32;
wire   [1:0] in_28;
wire   [1:0] in_23;
wire   [1:0] in_21;
wire   [1:0] in_18;
wire   [1:0] in_3;
wire   [1:0] in_2;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3948(.Y(out_0[9]), .A(n_131));
  ADDFX1 g3949(.CO(n_131), .S(out_0[5]), .A(n_93), .B(n_117), .CI(n_129));
  ADDFX1 g3950(.CO(n_129), .S(out_0[4]), .A(n_118), .B(n_119), .CI(n_127));
  ADDFX1 g3951(.CO(n_127), .S(out_0[3]), .A(n_123), .B(n_120), .CI(n_125));
  ADDFX1 g3952(.CO(n_125), .S(out_0[2]), .A(n_111), .B(n_121), .CI(n_124));
  ADDFX1 g3953(.CO(n_123), .S(n_124), .A(n_96), .B(n_114), .CI(n_108));
  ADDFX1 g3954(.CO(n_121), .S(out_0[1]), .A(n_97), .B(n_105), .CI(n_112));
  ADDFX1 g3955(.CO(n_119), .S(n_120), .A(n_110), .B(n_113), .CI(n_116));
  ADDFX1 g3956(.CO(n_117), .S(n_118), .A(n_100), .B(n_109), .CI(n_115));
  ADDFX1 g3957(.CO(n_115), .S(n_116), .A(n_89), .B(n_94), .CI(n_107));
  ADDFX1 g3958(.CO(n_113), .S(n_114), .A(n_92), .B(n_102), .CI(n_95));
  ADDFX1 g3959(.CO(n_111), .S(n_112), .A(n_87), .B(n_104), .CI(n_99));
  ADDFX1 g3960(.CO(n_109), .S(n_110), .A(n_81), .B(n_91), .CI(n_101));
  ADDFX1 g3961(.CO(n_107), .S(n_108), .A(n_65), .B(n_103), .CI(n_98));
  ADDFX1 g3962(.CO(n_105), .S(out_0[0]), .A(n_76), .B(n_84), .CI(n_88));
  ADDFX1 g3963(.CO(n_103), .S(n_104), .A(n_70), .B(n_86), .CI(n_75));
  ADDFX1 g3964(.CO(n_101), .S(n_102), .A(n_69), .B(n_85), .CI(n_82));
  XNOR2X1 g3965(.Y(n_100), .A(n_0), .B(n_90));
  ADDFX1 g3966(.CO(n_98), .S(n_99), .A(n_73), .B(n_72), .CI(n_83));
  ADDFX1 g3967(.CO(n_96), .S(n_97), .A(n_78), .B(n_80), .CI(n_66));
  ADDFX1 g3968(.CO(n_94), .S(n_95), .A(n_79), .B(n_68), .CI(n_77));
  NOR2BX1 g3969(.Y(n_93), .AN(n_90), .B(n_0));
  ADDFX1 g3970(.CO(n_91), .S(n_92), .A(n_47), .B(n_64), .CI(n_71));
  ADDFX1 g3971(.CO(n_90), .S(n_89), .A(n_24), .B(n_63), .CI(n_67));
  ADDFX1 g3972(.CO(n_87), .S(n_88), .A(n_30), .B(n_40), .CI(n_74));
  ADDFX1 g3973(.CO(n_85), .S(n_86), .A(n_11), .B(n_49), .CI(n_55));
  ADDFX1 g3974(.CO(n_83), .S(n_84), .A(n_46), .B(n_34), .CI(n_62));
  ADDFX1 g3975(.CO(n_81), .S(n_82), .A(n_23), .B(n_59), .CI(n_35));
  ADDFX1 g3976(.CO(n_79), .S(n_80), .A(n_43), .B(n_42), .CI(n_52));
  ADDFX1 g3977(.CO(n_77), .S(n_78), .A(n_58), .B(n_60), .CI(n_54));
  ADDFX1 g3978(.CO(n_75), .S(n_76), .A(in_1[0]), .B(n_56), .CI(n_44));
  ADDFX1 g3979(.CO(n_73), .S(n_74), .A(n_38), .B(n_50), .CI(n_32));
  ADDFX1 g3980(.CO(n_71), .S(n_72), .A(n_37), .B(n_33), .CI(n_45));
  ADDFX1 g3981(.CO(n_69), .S(n_70), .A(n_31), .B(n_29), .CI(n_61));
  ADDFX1 g3982(.CO(n_67), .S(n_68), .A(n_51), .B(n_53), .CI(n_41));
  ADDFX1 g3983(.CO(n_65), .S(n_66), .A(n_36), .B(n_48), .CI(n_39));
  ADDFX1 g3984(.CO(n_63), .S(n_64), .A(n_4), .B(n_12), .CI(n_57));
  ADDFX1 g3985(.CO(n_61), .S(n_62), .A(in_5[0]), .B(n_8), .CI(n_18));
  ADDFX1 g3986(.CO(n_59), .S(n_60), .A(n_20), .B(in_28[1]), .CI(n_5));
  ADDFX1 g3987(.CO(n_57), .S(n_58), .A(in_2[1]), .B(in_44[1]), .CI(in_18[0]));
  ADDFX1 g3988(.CO(n_55), .S(n_56), .A(in_16[0]), .B(n_17), .CI(n_9));
  INVX1 g3989(.Y(n_54), .A(n_28));
  INVX1 g3990(.Y(n_53), .A(n_27));
  INVX1 g3991(.Y(n_52), .A(n_26));
  INVX1 g3992(.Y(n_51), .A(n_25));
  ADDFX1 g3993(.CO(n_49), .S(n_50), .A(n_2), .B(n_16), .CI(in_23[0]));
  ADDFX1 g3994(.CO(n_47), .S(n_48), .A(in_36[1]), .B(n_15), .CI(in_15[1]));
  ADDFX1 g3995(.CO(n_45), .S(n_46), .A(in_6[0]), .B(in_10[0]), .CI(in_22[0]));
  ADDFX1 g3996(.CO(n_43), .S(n_44), .A(in_19), .B(n_6), .CI(n_21));
  ADDFX1 g3997(.CO(n_41), .S(n_42), .A(n_19), .B(n_3), .CI(in_37[0]));
  ADDFX1 g3998(.CO(n_39), .S(n_40), .A(in_35), .B(in_15[0]), .CI(in_7[0]));
  ADDFX1 g3999(.CO(n_37), .S(n_38), .A(in_18[0]), .B(in_3[0]), .CI(in_34[0]));
  ADDFX1 g4000(.CO(n_35), .S(n_36), .A(in_3[0]), .B(in_4[1]), .CI(in_43[1]));
  ADDFX1 g4001(.CO(n_33), .S(n_34), .A(in_13[0]), .B(in_27), .CI(n_7));
  ADDFX1 g4002(.CO(n_31), .S(n_32), .A(n_13), .B(n_14), .CI(in_37[0]));
  ADDFX1 g4003(.CO(n_29), .S(n_30), .A(in_21[0]), .B(in_32[0]), .CI(n_10));
  ADDFX1 g4004(.CO(n_27), .S(n_28), .A(in_33[1]), .B(in_39[1]), .CI(in_45[1]));
  ADDFX1 g4005(.CO(n_25), .S(n_26), .A(in_29[1]), .B(in_41[1]), .CI(in_46[1]));
  XNOR2X1 g4006(.Y(n_24), .A(in_37[0]), .B(n_22));
  OAI21X1 g4008(.Y(n_23), .A0(in_16[0]), .A1(in_22[0]), .B0(n_22));
  NAND2X1 g4009(.Y(n_22), .A(in_22[0]), .B(in_16[0]));
  INVX1 g4010(.Y(n_21), .A(in_26[0]));
  INVX1 g4011(.Y(n_20), .A(in_5[1]));
  INVX1 g4012(.Y(n_19), .A(in_0[1]));
  INVX1 g4013(.Y(n_18), .A(in_12[0]));
  INVX1 g4014(.Y(n_17), .A(in_40[0]));
  INVX1 g4015(.Y(n_16), .A(in_14[0]));
  INVX1 g4016(.Y(n_15), .A(in_7[1]));
  INVX1 g4017(.Y(n_14), .A(in_17[0]));
  INVX1 g4018(.Y(n_13), .A(in_11[0]));
  INVX1 g4019(.Y(n_12), .A(in_31[2]));
  INVX1 g4020(.Y(n_11), .A(in_1[0]));
  INVX1 g4021(.Y(n_10), .A(in_38[0]));
  INVX1 g4022(.Y(n_9), .A(in_47[0]));
  INVX1 g4023(.Y(n_8), .A(in_42[0]));
  INVX1 g4024(.Y(n_7), .A(in_30[0]));
  INVX1 g4025(.Y(n_6), .A(in_20[0]));
  INVX1 g4026(.Y(n_5), .A(in_25[1]));
  INVX1 g4027(.Y(n_4), .A(in_24[2]));
  INVX1 g4028(.Y(n_3), .A(in_8[1]));
  INVX1 g4029(.Y(n_2), .A(in_9[0]));
  NAND2BX1 g2(.Y(n_0), .AN(in_37[0]), .B(n_22));
endmodule

module WALLACE_CSA_DUMMY_OP752_group_359251(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, out_0);
input  in_20, in_25;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [4:0] in_4;
input   [2:0] in_5;
input   [4:0] in_6;
input   [6:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [1:0] in_18;
input   [4:0] in_19;
input   [1:0] in_21;
input   [4:0] in_22;
input   [1:0] in_23;
input   [1:0] in_24;
input   [4:0] in_26;
input   [2:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [1:0] in_38;
input   [1:0] in_39;
input   [2:0] in_40;
input   [4:0] in_41;
input   [1:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
output  [9:0] out_0;
wire  n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_45, n_43, n_41, n_39, 
    n_37, n_36, n_35, n_34, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_25, 
    in_20;
wire   [9:0] out_0;
wire   [1:0] in_42;
wire   [1:0] in_39;
wire   [1:0] in_38;
wire   [1:0] in_24;
wire   [1:0] in_23;
wire   [1:0] in_21;
wire   [1:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_7;
wire   [2:0] in_40;
wire   [2:0] in_30;
wire   [2:0] in_27;
wire   [2:0] in_5;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_41;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_22;
wire   [4:0] in_19;
wire   [4:0] in_6;
wire   [4:0] in_4;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  ADDFX1 cdnfadd_000_1(.CO(n_131), .S(n_130), .A(in_10[0]), .B(in_30[0]), .CI(
    in_38[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_129), .S(n_128), .A(in_35[0]), .B(n_22), .CI(in_25));
  ADDFX1 cdnfadd_000_3(.CO(n_127), .S(n_126), .A(in_18[0]), .B(in_37[0]), .CI(
    n_15));
  ADDFX1 cdnfadd_000_4(.CO(n_125), .S(n_124), .A(n_19), .B(n_16), .CI(in_42[0]));
  ADDFX1 cdnfadd_000_5(.CO(n_123), .S(n_122), .A(in_23[0]), .B(n_21), .CI(n_11));
  ADDFX1 cdnfadd_000_6(.CO(n_121), .S(n_120), .A(in_20), .B(in_11[0]), .CI(
    in_39[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_119), .S(n_118), .A(in_43[0]), .B(n_10), .CI(
    in_13[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_117), .S(n_116), .A(in_14[0]), .B(in_17[0]), .CI(
    in_9[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_97), .S(n_96), .A(in_12[0]), .B(in_7[0]), .CI(n_126));
  ADDFX1 cdnfadd_000_10(.CO(n_95), .S(n_132), .A(n_29), .B(n_128), .CI(n_118));
  ADDFX1 cdnfadd_000_11(.CO(n_94), .S(n_139), .A(n_120), .B(n_130), .CI(n_122));
  ADDFX1 cdnfadd_000_12(.CO(n_73), .S(n_133), .A(n_124), .B(n_116), .CI(n_96));
  ADDFX1 cdnfadd_001_0(.CO(n_115), .S(n_114), .A(n_20), .B(in_24[1]), .CI(
    in_8[1]));
  ADDFX1 cdnfadd_001_1(.CO(n_113), .S(n_112), .A(n_24), .B(n_7), .CI(n_6));
  ADDFX1 cdnfadd_001_2(.CO(n_111), .S(n_110), .A(n_18), .B(in_30[0]), .CI(
    in_27[1]));
  ADDFX1 cdnfadd_001_3(.CO(n_109), .S(n_108), .A(in_21[1]), .B(in_40[1]), .CI(
    n_3));
  ADDFX1 cdnfadd_001_4(.CO(n_107), .S(n_106), .A(n_23), .B(n_25), .CI(in_5[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_105), .S(n_104), .A(in_16[1]), .B(in_9[1]), .CI(n_9));
  ADDFX1 cdnfadd_001_6(.CO(n_103), .S(n_102), .A(n_4), .B(in_14[1]), .CI(
    in_36[1]));
  ADDFX1 cdnfadd_001_7(.CO(n_93), .S(n_92), .A(in_10[1]), .B(n_121), .CI(n_131));
  ADDFX1 cdnfadd_001_8(.CO(n_91), .S(n_90), .A(in_7[1]), .B(n_123), .CI(n_27));
  ADDFX1 cdnfadd_001_9(.CO(n_89), .S(n_88), .A(n_127), .B(n_129), .CI(n_119));
  ADDFX1 cdnfadd_001_10(.CO(n_87), .S(n_86), .A(n_125), .B(n_106), .CI(n_112));
  ADDFX1 cdnfadd_001_11(.CO(n_85), .S(n_84), .A(n_114), .B(n_110), .CI(n_108));
  ADDFX1 cdnfadd_001_12(.CO(n_83), .S(n_82), .A(n_104), .B(n_117), .CI(n_102));
  ADDFX1 cdnfadd_001_13(.CO(n_72), .S(n_71), .A(n_88), .B(n_94), .CI(n_90));
  ADDFX1 cdnfadd_001_14(.CO(n_70), .S(n_69), .A(n_97), .B(n_92), .CI(n_95));
  ADDFX1 cdnfadd_001_15(.CO(n_68), .S(n_140), .A(n_84), .B(n_86), .CI(n_82));
  ADDFX1 cdnfadd_001_16(.CO(n_53), .S(n_134), .A(n_73), .B(n_69), .CI(n_71));
  ADDFX1 cdnfadd_002_1(.CO(n_98), .S(n_101), .A(n_12), .B(n_13), .CI(n_14));
  ADDFX1 cdnfadd_002_2(.CO(n_100), .S(n_99), .A(n_1), .B(n_8), .CI(n_5));
  ADDFX1 cdnfadd_002_3(.CO(n_81), .S(n_80), .A(n_2), .B(n_28), .CI(n_107));
  ADDFX1 cdnfadd_002_4(.CO(n_79), .S(n_78), .A(n_17), .B(n_111), .CI(n_115));
  ADDFX1 cdnfadd_002_5(.CO(n_77), .S(n_76), .A(n_113), .B(n_109), .CI(n_105));
  ADDFX1 cdnfadd_002_6(.CO(n_75), .S(n_74), .A(n_101), .B(n_103), .CI(n_99));
  ADDFX1 cdnfadd_002_7(.CO(n_67), .S(n_66), .A(n_93), .B(n_89), .CI(n_91));
  ADDFX1 cdnfadd_002_8(.CO(n_65), .S(n_64), .A(n_85), .B(n_76), .CI(n_87));
  ADDFX1 cdnfadd_002_9(.CO(n_63), .S(n_62), .A(n_80), .B(n_78), .CI(n_83));
  ADDFX1 cdnfadd_002_10(.CO(n_57), .S(n_56), .A(n_74), .B(n_72), .CI(n_70));
  ADDFX1 cdnfadd_002_11(.CO(n_52), .S(n_141), .A(n_66), .B(n_62), .CI(n_64));
  ADDFX1 cdnfadd_002_12(.CO(n_142), .S(n_135), .A(n_68), .B(n_56), .CI(n_53));
  ADDFX1 cdnfadd_003_1(.CO(n_61), .S(n_60), .A(n_100), .B(n_81), .CI(n_79));
  ADDFX1 cdnfadd_003_2(.CO(n_59), .S(n_58), .A(n_77), .B(n_31), .CI(n_75));
  ADDFX1 cdnfadd_003_3(.CO(n_51), .S(n_50), .A(n_67), .B(n_65), .CI(n_60));
  ADDFX1 cdnfadd_003_4(.CO(n_49), .S(n_48), .A(n_58), .B(n_63), .CI(n_57));
  ADDFX1 cdnfadd_003_5(.CO(n_143), .S(n_136), .A(n_52), .B(n_50), .CI(n_48));
  ADDFX1 cdnfadd_004_0(.CO(n_55), .S(n_54), .A(n_30), .B(n_61), .CI(n_59));
  ADDFX1 cdnfadd_004_1(.CO(n_138), .S(n_137), .A(n_51), .B(n_54), .CI(n_49));
  NAND2X1 g327(.Y(out_0[9]), .A(n_35), .B(n_45));
  ADDFX1 g328(.CO(n_45), .S(out_0[5]), .A(n_36), .B(n_138), .CI(n_43));
  ADDFX1 g329(.CO(n_43), .S(out_0[4]), .A(n_143), .B(n_137), .CI(n_41));
  ADDFX1 g330(.CO(n_41), .S(out_0[3]), .A(n_142), .B(n_136), .CI(n_39));
  ADDFX1 g331(.CO(n_39), .S(out_0[2]), .A(n_141), .B(n_37), .CI(n_135));
  ADDFX1 g332(.CO(n_37), .S(out_0[1]), .A(n_140), .B(n_32), .CI(n_134));
  OAI21X1 g333(.Y(n_36), .A0(n_30), .A1(n_34), .B0(n_35));
  NAND2X1 g334(.Y(n_35), .A(n_30), .B(n_34));
  INVX1 g335(.Y(n_34), .A(n_55));
  ADDFX1 g336(.CO(n_32), .S(out_0[0]), .A(n_132), .B(n_139), .CI(n_133));
  AO21XL g337(.Y(n_31), .A0(n_26), .A1(n_98), .B0(n_30));
  NOR2X1 g338(.Y(n_30), .A(n_26), .B(n_98));
  OAI2BB1X1 g339(.Y(n_29), .A0N(in_29[0]), .A1N(in_19[0]), .B0(n_27));
  OAI21X1 g340(.Y(n_28), .A0(in_15[2]), .A1(in_35[0]), .B0(n_26));
  NAND2X1 g341(.Y(n_27), .A(n_12), .B(n_1));
  NAND2X1 g342(.Y(n_26), .A(in_35[0]), .B(in_15[2]));
  INVX1 g343(.Y(n_25), .A(in_6[1]));
  INVX1 g344(.Y(n_24), .A(in_31[1]));
  INVX1 g345(.Y(n_23), .A(in_44[1]));
  INVX1 g346(.Y(n_22), .A(in_22[0]));
  INVX1 g347(.Y(n_21), .A(in_1[0]));
  INVX1 g348(.Y(n_20), .A(in_3[1]));
  INVX1 g349(.Y(n_19), .A(in_0[0]));
  INVX1 g350(.Y(n_18), .A(in_41[1]));
  INVX1 g351(.Y(n_17), .A(in_7[2]));
  INVX1 g352(.Y(n_16), .A(in_28[0]));
  INVX1 g353(.Y(n_15), .A(in_34[0]));
  INVX1 g354(.Y(n_14), .A(in_43[0]));
  INVX1 g355(.Y(n_13), .A(in_37[0]));
  INVX1 g356(.Y(n_12), .A(in_29[0]));
  INVX1 g357(.Y(n_11), .A(in_2[0]));
  INVX1 g358(.Y(n_10), .A(in_32[0]));
  INVX1 g359(.Y(n_9), .A(in_12[1]));
  INVX1 g360(.Y(n_8), .A(in_10[2]));
  INVX1 g361(.Y(n_7), .A(in_4[1]));
  INVX1 g362(.Y(n_6), .A(in_33[1]));
  INVX1 g363(.Y(n_5), .A(in_14[2]));
  INVX1 g364(.Y(n_4), .A(in_17[1]));
  INVX1 g365(.Y(n_3), .A(in_26[1]));
  INVX1 g366(.Y(n_2), .A(in_36[1]));
  INVX1 g367(.Y(n_1), .A(in_19[0]));
endmodule

module WALLACE_CSA_DUMMY_OP754_group_359252(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, out_0);
input  in_24, in_26;
input   [4:0] in_0;
input   [4:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [4:0] in_15;
input   [2:0] in_16;
input   [4:0] in_17;
input   [1:0] in_18;
input   [1:0] in_19;
input   [1:0] in_20;
input   [1:0] in_21;
input   [1:0] in_22;
input   [2:0] in_23;
input   [1:0] in_25;
input   [4:0] in_27;
input   [3:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [2:0] in_33;
input   [1:0] in_34;
input   [2:0] in_35;
input   [1:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [4:0] in_40;
input   [1:0] in_41;
input   [1:0] in_42;
input   [1:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [2:0] in_46;
output  [9:0] out_0;
wire  n_133, n_130, n_128, n_126, n_125, n_124, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_26, 
    in_24;
wire   [9:0] out_0;
wire   [3:0] in_28;
wire   [1:0] in_45;
wire   [1:0] in_43;
wire   [1:0] in_42;
wire   [1:0] in_41;
wire   [1:0] in_37;
wire   [1:0] in_36;
wire   [1:0] in_34;
wire   [1:0] in_25;
wire   [1:0] in_22;
wire   [1:0] in_21;
wire   [1:0] in_20;
wire   [1:0] in_19;
wire   [1:0] in_18;
wire   [2:0] in_46;
wire   [2:0] in_39;
wire   [2:0] in_35;
wire   [2:0] in_33;
wire   [2:0] in_32;
wire   [2:0] in_30;
wire   [2:0] in_23;
wire   [2:0] in_16;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [4:0] in_44;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_17;
wire   [4:0] in_15;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  AO21X1 g4222(.Y(out_0[6]), .A0(n_113), .A1(n_133), .B0(out_0[9]));
  NOR2X1 g4223(.Y(out_0[9]), .A(n_113), .B(n_133));
  ADDFX1 g4224(.CO(n_133), .S(out_0[5]), .A(n_112), .B(n_120), .CI(n_130));
  ADDFX1 g4225(.CO(n_130), .S(out_0[4]), .A(n_121), .B(n_124), .CI(n_128));
  ADDFX1 g4226(.CO(n_128), .S(out_0[3]), .A(n_118), .B(n_125), .CI(n_126));
  ADDFX1 g4227(.CO(n_126), .S(out_0[2]), .A(n_108), .B(n_122), .CI(n_119));
  ADDFX1 g4228(.CO(n_124), .S(n_125), .A(n_107), .B(n_106), .CI(n_117));
  ADDFX1 g4229(.CO(n_122), .S(out_0[1]), .A(n_95), .B(n_98), .CI(n_115));
  ADDFX1 g4230(.CO(n_120), .S(n_121), .A(n_105), .B(n_111), .CI(n_116));
  ADDFX1 g4231(.CO(n_118), .S(n_119), .A(n_102), .B(n_110), .CI(n_114));
  ADDFX1 g4232(.CO(n_116), .S(n_117), .A(n_101), .B(n_104), .CI(n_109));
  ADDFX1 g4233(.CO(n_114), .S(n_115), .A(n_84), .B(n_88), .CI(n_100));
  INVX1 g4234(.Y(n_112), .A(n_113));
  ADDFX1 g4235(.CO(n_113), .S(n_111), .A(n_19), .B(n_89), .CI(n_103));
  ADDFX1 g4236(.CO(n_109), .S(n_110), .A(n_86), .B(n_94), .CI(n_99));
  ADDFX1 g4237(.CO(n_107), .S(n_108), .A(n_87), .B(n_92), .CI(n_97));
  ADDFX1 g4238(.CO(n_105), .S(n_106), .A(n_90), .B(n_91), .CI(n_85));
  ADDFX1 g4239(.CO(n_103), .S(n_104), .A(n_73), .B(n_79), .CI(n_93));
  ADDFX1 g4240(.CO(n_101), .S(n_102), .A(n_72), .B(n_81), .CI(n_83));
  ADDFX1 g4241(.CO(n_99), .S(n_100), .A(n_58), .B(n_69), .CI(n_76));
  ADDFX1 g4242(.CO(n_97), .S(n_98), .A(n_82), .B(n_62), .CI(n_77));
  ADDFX1 g4243(.CO(n_95), .S(out_0[0]), .A(n_64), .B(n_70), .CI(n_78));
  ADDFX1 g4244(.CO(n_93), .S(n_94), .A(n_25), .B(n_65), .CI(n_75));
  ADDFX1 g4245(.CO(n_91), .S(n_92), .A(n_74), .B(n_67), .CI(n_61));
  ADDFX1 g4246(.CO(n_89), .S(n_90), .A(n_20), .B(n_59), .CI(n_71));
  ADDFX1 g4247(.CO(n_87), .S(n_88), .A(n_66), .B(n_63), .CI(n_68));
  ADDFX1 g4248(.CO(n_85), .S(n_86), .A(n_57), .B(n_60), .CI(n_80));
  ADDFX1 g4249(.CO(n_83), .S(n_84), .A(n_54), .B(n_31), .CI(n_29));
  ADDFX1 g4250(.CO(n_81), .S(n_82), .A(n_56), .B(n_46), .CI(n_40));
  ADDFX1 g4251(.CO(n_79), .S(n_80), .A(n_18), .B(n_39), .CI(n_5));
  ADDFX1 g4252(.CO(n_77), .S(n_78), .A(n_24), .B(n_32), .CI(n_30));
  ADDFX1 g4253(.CO(n_75), .S(n_76), .A(n_37), .B(n_33), .CI(in_2[1]));
  ADDFX1 g4254(.CO(n_73), .S(n_74), .A(n_47), .B(n_41), .CI(n_55));
  ADDFX1 g4255(.CO(n_71), .S(n_72), .A(n_27), .B(n_53), .CI(n_45));
  ADDFX1 g4256(.CO(n_69), .S(n_70), .A(n_38), .B(n_50), .CI(n_36));
  ADDFX1 g4257(.CO(n_67), .S(n_68), .A(n_49), .B(n_42), .CI(n_28));
  ADDFX1 g4258(.CO(n_65), .S(n_66), .A(n_35), .B(n_21), .CI(n_43));
  ADDFX1 g4259(.CO(n_63), .S(n_64), .A(n_22), .B(n_44), .CI(n_34));
  ADDFX1 g4260(.CO(n_61), .S(n_62), .A(n_52), .B(n_48), .CI(n_26));
  ADDFX1 g4261(.CO(n_59), .S(n_60), .A(in_23[2]), .B(n_1), .CI(n_51));
  ADDFX1 g4262(.CO(n_57), .S(n_58), .A(in_9[1]), .B(n_13), .CI(n_23));
  ADDFX1 g4263(.CO(n_55), .S(n_56), .A(in_6[1]), .B(in_8[1]), .CI(in_21[1]));
  ADDFX1 g4264(.CO(n_53), .S(n_54), .A(in_30[1]), .B(in_36[1]), .CI(n_16));
  ADDFX1 g4265(.CO(n_51), .S(n_52), .A(in_34[1]), .B(in_16[1]), .CI(in_37[1]));
  ADDFX1 g4266(.CO(n_49), .S(n_50), .A(in_8[0]), .B(n_2), .CI(in_33[0]));
  ADDFX1 g4267(.CO(n_47), .S(n_48), .A(in_25[0]), .B(in_10[1]), .CI(n_8));
  ADDFX1 g4268(.CO(n_45), .S(n_46), .A(in_5[1]), .B(in_32[1]), .CI(in_45[0]));
  ADDFX1 g4269(.CO(n_43), .S(n_44), .A(in_26), .B(in_6[0]), .CI(n_9));
  ADDFX1 g4270(.CO(n_41), .S(n_42), .A(in_20[1]), .B(n_3), .CI(in_43[1]));
  ADDFX1 g4271(.CO(n_39), .S(n_40), .A(in_19[1]), .B(in_4[1]), .CI(in_35[0]));
  ADDFX1 g4272(.CO(n_37), .S(n_38), .A(in_10[0]), .B(n_4), .CI(n_7));
  ADDFX1 g4273(.CO(n_35), .S(n_36), .A(in_18[0]), .B(n_12), .CI(in_35[0]));
  ADDFX1 g4274(.CO(n_33), .S(n_34), .A(in_7[0]), .B(n_11), .CI(n_15));
  ADDFX1 g4275(.CO(n_31), .S(n_32), .A(in_25[0]), .B(in_45[0]), .CI(in_9[0]));
  ADDFX1 g4276(.CO(n_29), .S(n_30), .A(in_14[0]), .B(in_11[0]), .CI(in_2[0]));
  ADDFX1 g4277(.CO(n_27), .S(n_28), .A(in_22[1]), .B(n_10), .CI(in_39[0]));
  ADDFX1 g4278(.CO(n_25), .S(n_26), .A(in_12[1]), .B(in_42[1]), .CI(n_6));
  ADDFX1 g4279(.CO(n_23), .S(n_24), .A(in_24), .B(in_3[0]), .CI(in_41[0]));
  ADDFX1 g4280(.CO(n_21), .S(n_22), .A(in_39[0]), .B(in_13[0]), .CI(n_14));
  XNOR2X1 g4281(.Y(n_20), .A(in_28[0]), .B(n_17));
  NOR2X1 g4282(.Y(n_19), .A(n_9), .B(n_17));
  AO21X1 g4283(.Y(n_18), .A0(in_46[2]), .A1(in_33[0]), .B0(n_17));
  NOR2X1 g4284(.Y(n_17), .A(in_46[2]), .B(in_33[0]));
  INVX1 g4285(.Y(n_16), .A(in_38[1]));
  INVX1 g4286(.Y(n_15), .A(in_27[0]));
  INVX1 g4287(.Y(n_14), .A(in_40[0]));
  INVX1 g4288(.Y(n_13), .A(in_14[1]));
  INVX1 g4289(.Y(n_12), .A(in_1[0]));
  INVX1 g4290(.Y(n_11), .A(in_17[0]));
  INVX1 g4291(.Y(n_10), .A(in_0[1]));
  INVX1 g4292(.Y(n_9), .A(in_28[0]));
  INVX1 g4293(.Y(n_8), .A(in_31[1]));
  INVX1 g4294(.Y(n_7), .A(in_44[0]));
  INVX1 g4295(.Y(n_6), .A(in_11[1]));
  INVX1 g4296(.Y(n_5), .A(in_2[2]));
  INVX1 g4297(.Y(n_4), .A(in_29[0]));
  INVX1 g4298(.Y(n_3), .A(in_13[1]));
  INVX1 g4299(.Y(n_2), .A(in_15[0]));
  INVX1 g4300(.Y(n_1), .A(in_9[2]));
endmodule

module WALLACE_CSA_DUMMY_OP758_group_359250(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, out_0);
input  in_29, in_34, in_35;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [6:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [4:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [1:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [1:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [2:0] in_27;
input   [4:0] in_28;
input   [2:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [4:0] in_33;
input   [4:0] in_36;
input   [4:0] in_37;
input   [1:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [1:0] in_42;
input   [4:0] in_43;
output  [9:0] out_0;
wire  n_136, n_134, n_132, n_130, n_129, n_128, n_127, n_126, n_124, n_123, 
    n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
    n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, 
    n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, 
    n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
    n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_0, in_35, in_34, in_29;
wire   [9:0] out_0;
wire   [1:0] in_42;
wire   [1:0] in_38;
wire   [1:0] in_23;
wire   [1:0] in_22;
wire   [1:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [6:0] in_5;
wire   [2:0] in_32;
wire   [2:0] in_30;
wire   [2:0] in_27;
wire   [2:0] in_3;
wire   [4:0] in_43;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_10;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1659(.Y(out_0[9]), .A(n_136));
  ADDFX1 g1660(.CO(n_136), .S(out_0[5]), .A(n_110), .B(n_126), .CI(n_134));
  ADDFX1 g1661(.CO(n_134), .S(out_0[4]), .A(n_128), .B(n_127), .CI(n_132));
  ADDFX1 g1662(.CO(n_132), .S(out_0[3]), .A(n_122), .B(n_129), .CI(n_130));
  ADDFX1 g1663(.CO(n_130), .S(out_0[2]), .A(n_119), .B(n_124), .CI(n_123));
  ADDFX1 g1664(.CO(n_128), .S(n_129), .A(n_113), .B(n_118), .CI(n_121));
  ADDFX1 g1665(.CO(n_126), .S(n_127), .A(n_111), .B(n_112), .CI(n_120));
  ADDFX1 g1666(.CO(n_124), .S(out_0[1]), .A(n_107), .B(n_108), .CI(n_117));
  ADDFX1 g1667(.CO(n_122), .S(n_123), .A(n_106), .B(n_116), .CI(n_115));
  ADDFX1 g1668(.CO(n_120), .S(n_121), .A(n_104), .B(n_97), .CI(n_114));
  ADDFX1 g1669(.CO(n_118), .S(n_119), .A(n_100), .B(n_105), .CI(n_95));
  ADDFX1 g1670(.CO(n_116), .S(n_117), .A(n_101), .B(n_90), .CI(n_103));
  ADDFX1 g1671(.CO(n_114), .S(n_115), .A(n_92), .B(n_99), .CI(n_102));
  ADDFX1 g1672(.CO(n_112), .S(n_113), .A(n_76), .B(n_98), .CI(n_94));
  ADDFX1 g1673(.CO(n_110), .S(n_111), .A(n_21), .B(n_67), .CI(n_96));
  ADDFX1 g1674(.CO(n_108), .S(out_0[0]), .A(n_79), .B(n_73), .CI(n_91));
  ADDFX1 g1675(.CO(n_106), .S(n_107), .A(n_75), .B(n_89), .CI(n_93));
  ADDFX1 g1676(.CO(n_104), .S(n_105), .A(n_74), .B(n_88), .CI(n_77));
  ADDFX1 g1677(.CO(n_102), .S(n_103), .A(n_78), .B(n_82), .CI(n_63));
  ADDFX1 g1678(.CO(n_100), .S(n_101), .A(n_71), .B(n_85), .CI(n_87));
  ADDFX1 g1679(.CO(n_98), .S(n_99), .A(n_65), .B(n_86), .CI(n_70));
  ADDFX1 g1680(.CO(n_96), .S(n_97), .A(n_80), .B(n_0), .CI(n_68));
  ADDFX1 g1681(.CO(n_94), .S(n_95), .A(n_81), .B(n_84), .CI(n_69));
  ADDFX1 g1682(.CO(n_92), .S(n_93), .A(n_37), .B(n_66), .CI(n_72));
  ADDFX1 g1683(.CO(n_90), .S(n_91), .A(n_38), .B(n_83), .CI(n_64));
  ADDFX1 g1684(.CO(n_88), .S(n_89), .A(n_28), .B(n_49), .CI(n_34));
  ADDFX1 g1685(.CO(n_86), .S(n_87), .A(n_23), .B(n_55), .CI(n_57));
  ADDFX1 g1686(.CO(n_84), .S(n_85), .A(n_42), .B(n_46), .CI(in_5[1]));
  ADDFX1 g1687(.CO(n_82), .S(n_83), .A(n_24), .B(n_36), .CI(n_54));
  ADDFX1 g1689(.CO(n_80), .S(n_81), .A(n_27), .B(n_25), .CI(n_59));
  ADDFX1 g1690(.CO(n_78), .S(n_79), .A(n_30), .B(n_56), .CI(n_58));
  ADDFX1 g1691(.CO(n_76), .S(n_77), .A(n_52), .B(n_45), .CI(n_33));
  ADDFX1 g1692(.CO(n_74), .S(n_75), .A(n_29), .B(n_26), .CI(n_60));
  ADDFX1 g1693(.CO(n_72), .S(n_73), .A(n_32), .B(n_47), .CI(n_41));
  ADDFX1 g1694(.CO(n_70), .S(n_71), .A(n_31), .B(n_53), .CI(n_40));
  ADDFX1 g1696(.CO(n_68), .S(n_69), .A(n_22), .B(n_48), .CI(n_9));
  OAI22X1 g1697(.Y(n_67), .A0(n_44), .A1(n_61), .B0(n_21), .B1(n_51));
  ADDFX1 g1698(.CO(n_65), .S(n_66), .A(in_16[1]), .B(n_5), .CI(n_35));
  ADDFX1 g1699(.CO(n_63), .S(n_64), .A(in_14[0]), .B(n_43), .CI(in_5[0]));
  XNOR2X1 g1700(.Y(n_62), .A(n_44), .B(n_51));
  AND2XL g1701(.Y(n_61), .A(n_21), .B(n_51));
  ADDFX1 g1702(.CO(n_59), .S(n_60), .A(in_22[0]), .B(in_6[0]), .CI(in_27[1]));
  ADDFX1 g1703(.CO(n_57), .S(n_58), .A(in_25[0]), .B(n_15), .CI(in_26[0]));
  ADDFX1 g1704(.CO(n_55), .S(n_56), .A(in_32[0]), .B(n_6), .CI(in_33[0]));
  ADDFX1 g1705(.CO(n_53), .S(n_54), .A(n_4), .B(n_20), .CI(in_15[0]));
  INVX1 g1706(.Y(n_52), .A(n_50));
  ADDFX1 g1707(.CO(n_51), .S(n_50), .A(in_25[0]), .B(in_33[0]), .CI(in_40[0]));
  ADDFX1 g1708(.CO(n_48), .S(n_49), .A(in_23[1]), .B(n_13), .CI(n_8));
  ADDFX1 g1709(.CO(n_46), .S(n_47), .A(in_17[0]), .B(n_3), .CI(in_35));
  INVX1 g1710(.Y(n_45), .A(n_39));
  ADDFX1 g1711(.CO(n_42), .S(n_43), .A(in_10[0]), .B(n_11), .CI(n_19));
  ADDFX1 g1712(.CO(n_40), .S(n_41), .A(in_3[0]), .B(n_17), .CI(in_43[0]));
  ADDFX1 g1713(.CO(n_44), .S(n_39), .A(in_10[0]), .B(in_26[0]), .CI(in_43[0]));
  ADDFX1 g1714(.CO(n_37), .S(n_38), .A(in_9[0]), .B(in_16[0]), .CI(in_12[0]));
  ADDFX1 g1715(.CO(n_35), .S(n_36), .A(in_34), .B(in_8[0]), .CI(in_40[0]));
  ADDFX1 g1716(.CO(n_33), .S(n_34), .A(in_11[1]), .B(n_2), .CI(n_18));
  ADDFX1 g1717(.CO(n_31), .S(n_32), .A(in_6[0]), .B(n_16), .CI(n_7));
  ADDFX1 g1718(.CO(n_29), .S(n_30), .A(in_29), .B(n_10), .CI(in_38[0]));
  ADDFX1 g1719(.CO(n_27), .S(n_28), .A(in_13[1]), .B(n_14), .CI(in_32[0]));
  ADDFX1 g1720(.CO(n_25), .S(n_26), .A(in_3[0]), .B(in_7[1]), .CI(in_15[0]));
  ADDFX1 g1721(.CO(n_23), .S(n_24), .A(in_22[0]), .B(in_42[0]), .CI(n_12));
  XNOR2X1 g1722(.Y(n_22), .A(in_30[2]), .B(in_15[0]));
  NOR2BX1 g1723(.Y(n_21), .AN(in_30[2]), .B(in_15[0]));
  INVX1 g1724(.Y(n_20), .A(in_41[0]));
  INVX1 g1725(.Y(n_19), .A(in_39[0]));
  INVX1 g1726(.Y(n_18), .A(in_14[1]));
  INVX1 g1727(.Y(n_17), .A(in_24[0]));
  INVX1 g1728(.Y(n_16), .A(in_2[0]));
  INVX1 g1729(.Y(n_15), .A(in_0[0]));
  INVX1 g1730(.Y(n_14), .A(in_31[1]));
  INVX1 g1731(.Y(n_13), .A(in_21[1]));
  INVX1 g1732(.Y(n_12), .A(in_37[0]));
  INVX1 g1733(.Y(n_11), .A(in_19[0]));
  INVX1 g1734(.Y(n_10), .A(in_1[0]));
  INVX1 g1735(.Y(n_9), .A(in_5[2]));
  INVX1 g1736(.Y(n_8), .A(in_28[1]));
  INVX1 g1737(.Y(n_7), .A(in_36[0]));
  INVX1 g1738(.Y(n_6), .A(in_18[0]));
  INVX1 g1739(.Y(n_5), .A(in_9[1]));
  INVX1 g1740(.Y(n_4), .A(in_20[0]));
  INVX1 g1741(.Y(n_3), .A(in_4[0]));
  INVX1 g1742(.Y(n_2), .A(in_12[1]));
  CLKXOR2X1 g2(.Y(n_0), .A(n_21), .B(n_62));
endmodule

module WALLACE_CSA_DUMMY_OP791_group_359281(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, out_0);
input  in_23, in_31;
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [4:0] in_4;
input   [4:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [1:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [1:0] in_32;
input   [1:0] in_33;
input   [1:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
output  [9:0] out_0;
wire  n_108, n_106, n_104, n_102, n_101, n_100, n_99, n_98, n_96, n_95, n_94, 
    n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, 
    n_81, n_80, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, 
    n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, 
    n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
    n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, 
    n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, 
    n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, 
    n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_31, in_23;
wire   [9:0] out_0;
wire   [2:0] in_39;
wire   [1:0] in_34;
wire   [1:0] in_33;
wire   [1:0] in_32;
wire   [1:0] in_29;
wire   [1:0] in_26;
wire   [1:0] in_24;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_25;
wire   [4:0] in_5;
wire   [4:0] in_4;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g3391(.Y(out_0[9]), .A(n_108));
  ADDFX1 g3392(.CO(n_108), .S(out_0[5]), .A(n_72), .B(n_98), .CI(n_106));
  ADDFX1 g3393(.CO(n_106), .S(out_0[4]), .A(n_99), .B(n_100), .CI(n_104));
  ADDFX1 g3394(.CO(n_104), .S(out_0[3]), .A(n_94), .B(n_101), .CI(n_102));
  ADDFX1 g3395(.CO(n_102), .S(out_0[2]), .A(n_93), .B(n_96), .CI(n_95));
  ADDFX1 g3396(.CO(n_100), .S(n_101), .A(n_87), .B(n_92), .CI(n_91));
  ADDFX1 g3397(.CO(n_98), .S(n_99), .A(n_73), .B(n_86), .CI(n_90));
  ADDFX1 g3398(.CO(n_96), .S(out_0[1]), .A(n_78), .B(n_83), .CI(n_89));
  ADDFX1 g3399(.CO(n_94), .S(n_95), .A(n_77), .B(n_81), .CI(n_88));
  ADDFX1 g3400(.CO(n_92), .S(n_93), .A(n_84), .B(n_82), .CI(n_75));
  ADDFX1 g3401(.CO(n_90), .S(n_91), .A(n_74), .B(n_76), .CI(n_80));
  ADDFX1 g3402(.CO(n_88), .S(n_89), .A(n_56), .B(n_70), .CI(n_85));
  ADDFX1 g3403(.CO(n_86), .S(n_87), .A(n_51), .B(n_59), .CI(n_71));
  ADDFX1 g3404(.CO(n_84), .S(n_85), .A(n_54), .B(n_67), .CI(n_65));
  ADDFX1 g3405(.CO(n_82), .S(n_83), .A(n_49), .B(n_58), .CI(n_62));
  ADDFX1 g3406(.CO(n_80), .S(n_81), .A(n_61), .B(n_60), .CI(n_69));
  ADDFX1 g3407(.CO(n_78), .S(out_0[0]), .A(n_50), .B(n_66), .CI(n_68));
  ADDFX1 g3408(.CO(n_76), .S(n_77), .A(n_53), .B(n_64), .CI(n_55));
  ADDFX1 g3409(.CO(n_74), .S(n_75), .A(n_47), .B(n_57), .CI(n_52));
  INVX1 g3410(.Y(n_73), .A(n_72));
  ADDFX1 g3411(.CO(n_72), .S(n_71), .A(n_7), .B(n_15), .CI(n_63));
  ADDFX1 g3412(.CO(n_69), .S(n_70), .A(n_30), .B(n_44), .CI(n_48));
  ADDFX1 g3413(.CO(n_67), .S(n_68), .A(n_34), .B(n_40), .CI(n_20));
  ADDFX1 g3414(.CO(n_65), .S(n_66), .A(n_36), .B(n_46), .CI(n_22));
  ADDFX1 g3415(.CO(n_63), .S(n_64), .A(n_41), .B(n_37), .CI(n_29));
  ADDFX1 g3416(.CO(n_61), .S(n_62), .A(n_45), .B(n_39), .CI(n_38));
  ADDFX1 g3417(.CO(n_59), .S(n_60), .A(n_43), .B(n_18), .CI(n_23));
  ADDFX1 g3418(.CO(n_57), .S(n_58), .A(n_21), .B(n_33), .CI(n_25));
  ADDFX1 g3419(.CO(n_55), .S(n_56), .A(n_42), .B(n_28), .CI(n_24));
  ADDFX1 g3420(.CO(n_53), .S(n_54), .A(in_20[1]), .B(n_35), .CI(n_19));
  ADDFX1 g3421(.CO(n_51), .S(n_52), .A(n_16), .B(n_5), .CI(n_27));
  ADDFX1 g3422(.CO(n_49), .S(n_50), .A(n_8), .B(in_12[0]), .CI(n_26));
  ADDFX1 g3423(.CO(n_47), .S(n_48), .A(in_26[0]), .B(n_17), .CI(in_11[1]));
  ADDFX1 g3424(.CO(n_45), .S(n_46), .A(in_29[0]), .B(n_9), .CI(in_35[0]));
  ADDFX1 g3425(.CO(n_43), .S(n_44), .A(in_6[1]), .B(n_1), .CI(in_33[1]));
  ADDFX1 g3426(.CO(n_41), .S(n_42), .A(n_6), .B(n_12), .CI(in_39[1]));
  ADDFX1 g3427(.CO(n_39), .S(n_40), .A(in_15[0]), .B(in_11[0]), .CI(in_23));
  ADDFX1 g3428(.CO(n_37), .S(n_38), .A(in_24[1]), .B(in_32[1]), .CI(n_11));
  ADDFX1 g3429(.CO(n_35), .S(n_36), .A(in_21[0]), .B(in_19[0]), .CI(n_14));
  INVX1 g3430(.Y(n_34), .A(n_32));
  INVX1 g3431(.Y(n_33), .A(n_31));
  ADDFX1 g3432(.CO(n_31), .S(n_32), .A(in_0[0]), .B(in_2[0]), .CI(in_27[0]));
  ADDFX1 g3433(.CO(n_29), .S(n_30), .A(in_22[1]), .B(in_7[1]), .CI(in_34[1]));
  ADDFX1 g3434(.CO(n_27), .S(n_28), .A(in_15[1]), .B(in_10[1]), .CI(in_16[1]));
  ADDFX1 g3435(.CO(n_25), .S(n_26), .A(in_9[0]), .B(in_8[0]), .CI(n_13));
  ADDFX1 g3436(.CO(n_23), .S(n_24), .A(n_10), .B(in_35[0]), .CI(in_12[1]));
  ADDFX1 g3437(.CO(n_21), .S(n_22), .A(n_2), .B(n_4), .CI(in_31));
  ADDFX1 g3438(.CO(n_19), .S(n_20), .A(in_13[0]), .B(n_3), .CI(in_20[0]));
  OAI21X1 g3439(.Y(n_18), .A0(in_12[2]), .A1(in_20[2]), .B0(n_15));
  XOR2XL g3440(.Y(n_17), .A(in_38[1]), .B(in_36[1]));
  NOR2X1 g3441(.Y(n_16), .A(in_38[1]), .B(in_36[1]));
  NAND2X1 g3442(.Y(n_15), .A(in_12[2]), .B(in_20[2]));
  INVX1 g3443(.Y(n_14), .A(in_28[0]));
  INVX1 g3444(.Y(n_13), .A(in_37[0]));
  INVX1 g3445(.Y(n_12), .A(in_1[1]));
  INVX1 g3446(.Y(n_11), .A(in_30[1]));
  INVX1 g3447(.Y(n_10), .A(in_5[1]));
  INVX1 g3448(.Y(n_9), .A(in_3[0]));
  INVX1 g3449(.Y(n_8), .A(in_26[0]));
  INVX1 g3450(.Y(n_7), .A(in_35[0]));
  INVX1 g3451(.Y(n_6), .A(in_17[1]));
  INVX1 g3452(.Y(n_5), .A(in_11[2]));
  INVX1 g3453(.Y(n_4), .A(in_14[0]));
  INVX1 g3454(.Y(n_3), .A(in_18[0]));
  INVX1 g3455(.Y(n_2), .A(in_4[0]));
  INVX1 g3456(.Y(n_1), .A(in_25[1]));
endmodule

module WALLACE_CSA_DUMMY_OP800_group_359276(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, out_0);
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [7:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [1:0] in_14;
input   [4:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [1:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [2:0] in_33;
input   [4:0] in_34;
output  [9:0] out_0;
wire  n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_46, n_44, n_42, n_40, n_38, n_37, n_36, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [9:0] out_0;
wire   [2:0] in_33;
wire   [1:0] in_31;
wire   [1:0] in_27;
wire   [1:0] in_21;
wire   [1:0] in_20;
wire   [1:0] in_14;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [7:0] in_4;
wire   [4:0] in_34;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_15;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_106), .S(n_86), .A(in_19[0]), .B(in_7[0]), .CI(n_6));
  ADDFX1 cdnfadd_000_2(.CO(n_85), .S(n_84), .A(n_31), .B(in_30[0]), .CI(n_17));
  ADDFX1 cdnfadd_000_3(.CO(n_105), .S(n_104), .A(in_27[0]), .B(in_5[0]), .CI(
    in_33[0]));
  ADDFX1 cdnfadd_000_4(.CO(n_103), .S(n_102), .A(n_5), .B(in_9[0]), .CI(n_3));
  ADDFX1 cdnfadd_000_5(.CO(n_101), .S(n_100), .A(n_2), .B(n_18), .CI(in_29[0]));
  ADDFX1 cdnfadd_000_6(.CO(n_99), .S(n_98), .A(n_15), .B(in_31[0]), .CI(in_22[0]));
  ADDFX1 cdnfadd_000_7(.CO(n_97), .S(n_96), .A(in_14[0]), .B(in_11[0]), .CI(n_1));
  ADDFX1 cdnfadd_000_8(.CO(n_95), .S(n_107), .A(n_13), .B(in_18[0]), .CI(in_4[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_76), .S(n_108), .A(n_102), .B(n_84), .CI(n_98));
  ADDFX1 cdnfadd_000_10(.CO(n_83), .S(n_114), .A(n_100), .B(n_96), .CI(n_104));
  ADDFX1 cdnfadd_001_0(.CO(n_94), .S(n_93), .A(n_10), .B(n_7), .CI(n_19));
  ADDFX1 cdnfadd_001_1(.CO(n_82), .S(n_81), .A(n_24), .B(n_106), .CI(n_93));
  ADDFX1 cdnfadd_001_2(.CO(n_73), .S(n_72), .A(n_30), .B(n_81), .CI(n_16));
  ADDFX1 cdnfadd_001_3(.CO(n_92), .S(n_91), .A(n_4), .B(n_8), .CI(in_29[0]));
  ADDFX1 cdnfadd_001_4(.CO(n_90), .S(n_89), .A(n_14), .B(in_33[0]), .CI(in_21[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_88), .S(n_87), .A(in_20[1]), .B(in_6[1]), .CI(
    in_18[1]));
  ADDFX1 cdnfadd_001_6(.CO(n_75), .S(n_74), .A(n_85), .B(n_101), .CI(n_103));
  ADDFX1 cdnfadd_001_7(.CO(n_65), .S(n_64), .A(n_99), .B(n_72), .CI(n_105));
  ADDFX1 cdnfadd_001_8(.CO(n_80), .S(n_79), .A(n_97), .B(n_89), .CI(n_87));
  ADDFX1 cdnfadd_001_9(.CO(n_78), .S(n_77), .A(n_91), .B(in_4[1]), .CI(n_95));
  ADDFX1 cdnfadd_001_10(.CO(n_53), .S(n_115), .A(n_83), .B(n_74), .CI(n_64));
  ADDFX1 cdnfadd_001_11(.CO(n_61), .S(n_109), .A(n_76), .B(n_79), .CI(n_77));
  ADDFX1 cdnfadd_002_1(.CO(n_71), .S(n_70), .A(n_94), .B(n_26), .CI(n_82));
  ADDFX1 cdnfadd_002_2(.CO(n_69), .S(n_68), .A(n_12), .B(n_11), .CI(n_70));
  ADDFX1 cdnfadd_002_3(.CO(n_63), .S(n_62), .A(n_92), .B(n_73), .CI(n_90));
  ADDFX1 cdnfadd_002_4(.CO(n_55), .S(n_54), .A(n_88), .B(n_68), .CI(n_65));
  ADDFX1 cdnfadd_002_5(.CO(n_60), .S(n_59), .A(in_4[2]), .B(n_75), .CI(n_80));
  ADDFX1 cdnfadd_002_6(.CO(n_49), .S(n_116), .A(n_62), .B(n_78), .CI(n_54));
  ADDFX1 cdnfadd_002_7(.CO(n_117), .S(n_110), .A(n_59), .B(n_53), .CI(n_61));
  ADDFX1 cdnfadd_003_0(.CO(n_67), .S(n_66), .A(n_29), .B(in_29[0]), .CI(n_71));
  ADDFX1 cdnfadd_003_1(.CO(n_58), .S(n_57), .A(n_69), .B(n_66), .CI(n_63));
  ADDFX1 cdnfadd_003_2(.CO(n_51), .S(n_50), .A(in_4[3]), .B(n_55), .CI(n_57));
  ADDFX1 cdnfadd_003_3(.CO(n_112), .S(n_111), .A(n_60), .B(n_49), .CI(n_50));
  ADDFX1 cdnfadd_004_1(.CO(n_52), .S(n_56), .A(n_67), .B(n_33), .CI(n_9));
  ADDFX1 cdnfadd_004_2(.CO(n_113), .S(n_118), .A(n_56), .B(n_58), .CI(n_51));
  NAND2BX1 g338(.Y(out_0[9]), .AN(n_36), .B(n_46));
  ADDFX1 g339(.CO(n_46), .S(out_0[5]), .A(n_37), .B(n_113), .CI(n_44));
  ADDFX1 g340(.CO(n_44), .S(out_0[4]), .A(n_118), .B(n_112), .CI(n_42));
  ADDFX1 g341(.CO(n_42), .S(out_0[3]), .A(n_117), .B(n_111), .CI(n_40));
  ADDFX1 g342(.CO(n_40), .S(out_0[2]), .A(n_38), .B(n_116), .CI(n_110));
  ADDFX1 g343(.CO(n_38), .S(out_0[1]), .A(n_34), .B(n_109), .CI(n_115));
  AO21X1 g344(.Y(n_37), .A0(n_32), .A1(n_52), .B0(n_36));
  NOR2X1 g345(.Y(n_36), .A(n_32), .B(n_52));
  ADDFX1 g346(.CO(n_34), .S(out_0[0]), .A(n_107), .B(n_114), .CI(n_108));
  OAI21X1 g347(.Y(n_33), .A0(in_29[0]), .A1(n_27), .B0(n_32));
  NAND2X1 g348(.Y(n_32), .A(in_29[0]), .B(n_27));
  OAI21X1 g349(.Y(n_31), .A0(n_22), .A1(n_28), .B0(n_30));
  NAND2X1 g350(.Y(n_30), .A(n_22), .B(n_28));
  OA21X1 g351(.Y(n_29), .A0(n_21), .A1(n_25), .B0(n_27));
  INVX1 g352(.Y(n_28), .A(n_86));
  NAND2X1 g353(.Y(n_27), .A(n_21), .B(n_25));
  OAI2BB1X1 g354(.Y(n_26), .A0N(n_20), .A1N(n_23), .B0(n_25));
  OR2X1 g355(.Y(n_25), .A(n_20), .B(n_23));
  AOI21X1 g356(.Y(n_24), .A0(in_16[1]), .A1(in_17[1]), .B0(n_20));
  XOR2XL g357(.Y(n_23), .A(in_7[0]), .B(in_19[0]));
  XNOR2X1 g358(.Y(n_22), .A(in_12[0]), .B(in_13[0]));
  NOR2XL g359(.Y(n_21), .A(in_7[0]), .B(in_19[0]));
  NOR2X1 g360(.Y(n_20), .A(in_17[1]), .B(in_16[1]));
  NOR2X1 g361(.Y(n_19), .A(in_13[0]), .B(in_12[0]));
  INVX1 g362(.Y(n_18), .A(in_15[0]));
  INVX1 g363(.Y(n_17), .A(in_26[0]));
  INVX1 g364(.Y(n_16), .A(in_24[1]));
  INVX1 g365(.Y(n_15), .A(in_25[0]));
  INVX1 g366(.Y(n_14), .A(in_0[1]));
  INVX1 g367(.Y(n_13), .A(in_32[0]));
  INVX1 g368(.Y(n_12), .A(in_22[0]));
  INVX1 g369(.Y(n_11), .A(in_30[0]));
  INVX1 g370(.Y(n_10), .A(in_5[1]));
  INVX1 g371(.Y(n_9), .A(in_4[4]));
  INVX1 g372(.Y(n_8), .A(in_23[1]));
  INVX1 g373(.Y(n_7), .A(in_8[1]));
  INVX1 g374(.Y(n_6), .A(in_10[0]));
  INVX1 g375(.Y(n_5), .A(in_2[0]));
  INVX1 g376(.Y(n_4), .A(in_28[1]));
  INVX1 g377(.Y(n_3), .A(in_1[0]));
  INVX1 g378(.Y(n_2), .A(in_34[0]));
  INVX1 g379(.Y(n_1), .A(in_3[0]));
endmodule

module WALLACE_CSA_DUMMY_OP818_group_359286(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, out_0);
input   [4:0] in_0;
input   [4:0] in_1;
input   [4:0] in_2;
input   [2:0] in_3;
input   [4:0] in_4;
input   [6:0] in_5;
input   [4:0] in_6;
input   [2:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [1:0] in_17;
input   [1:0] in_18;
input   [2:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [2:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [4:0] in_33;
input   [2:0] in_34;
input   [4:0] in_35;
input   [2:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [4:0] in_40;
input   [2:0] in_41;
input   [2:0] in_42;
input   [4:0] in_43;
input   [1:0] in_44;
output  [9:0] out_0;
wire  n_125, n_123, n_121, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_0;
wire   [9:0] out_0;
wire   [1:0] in_44;
wire   [1:0] in_29;
wire   [1:0] in_27;
wire   [1:0] in_18;
wire   [1:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [6:0] in_5;
wire   [2:0] in_42;
wire   [2:0] in_41;
wire   [2:0] in_39;
wire   [2:0] in_36;
wire   [2:0] in_34;
wire   [2:0] in_32;
wire   [2:0] in_22;
wire   [2:0] in_19;
wire   [2:0] in_7;
wire   [2:0] in_3;
wire   [4:0] in_43;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_6;
wire   [4:0] in_4;
wire   [4:0] in_2;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1556(.Y(out_0[9]), .A(n_125));
  ADDFX1 g1557(.CO(n_125), .S(out_0[5]), .A(n_89), .B(n_115), .CI(n_123));
  ADDFX1 g1558(.CO(n_123), .S(out_0[4]), .A(n_116), .B(n_117), .CI(n_121));
  ADDFX1 g1559(.CO(n_121), .S(out_0[3]), .A(n_113), .B(n_118), .CI(n_119));
  ADDFX1 g1560(.CO(n_119), .S(out_0[2]), .A(n_101), .B(n_114), .CI(n_111));
  ADDFX1 g1561(.CO(n_117), .S(n_118), .A(n_108), .B(n_105), .CI(n_110));
  ADDFX1 g1562(.CO(n_115), .S(n_116), .A(n_96), .B(n_107), .CI(n_109));
  ADDFX1 g1563(.CO(n_113), .S(n_114), .A(n_97), .B(n_104), .CI(n_106));
  ADDFX1 g1564(.CO(n_111), .S(out_0[1]), .A(n_99), .B(n_98), .CI(n_102));
  ADDFX1 g1565(.CO(n_109), .S(n_110), .A(n_87), .B(n_90), .CI(n_103));
  ADDFX1 g1566(.CO(n_107), .S(n_108), .A(n_75), .B(n_92), .CI(n_83));
  ADDFX1 g1567(.CO(n_105), .S(n_106), .A(n_93), .B(n_84), .CI(n_91));
  ADDFX1 g1568(.CO(n_103), .S(n_104), .A(n_65), .B(n_94), .CI(n_85));
  ADDFX1 g1569(.CO(n_101), .S(n_102), .A(n_81), .B(n_95), .CI(n_86));
  ADDFX1 g1570(.CO(n_99), .S(out_0[0]), .A(n_74), .B(n_78), .CI(n_82));
  ADDFX1 g1571(.CO(n_97), .S(n_98), .A(n_68), .B(n_70), .CI(n_66));
  OAI2BB1X1 g1572(.Y(n_96), .A0N(n_56), .A1N(n_88), .B0(n_89));
  ADDFX1 g1573(.CO(n_94), .S(n_95), .A(n_72), .B(n_60), .CI(n_73));
  ADDFX1 g1574(.CO(n_92), .S(n_93), .A(n_25), .B(n_58), .CI(n_71));
  ADDFX1 g1575(.CO(n_90), .S(n_91), .A(n_69), .B(n_80), .CI(n_67));
  OR2X1 g1576(.Y(n_89), .A(n_56), .B(n_88));
  ADDFX1 g1577(.CO(n_88), .S(n_87), .A(n_57), .B(n_0), .CI(n_79));
  ADDFX1 g1578(.CO(n_85), .S(n_86), .A(n_77), .B(n_62), .CI(n_63));
  ADDFX1 g1579(.CO(n_83), .S(n_84), .A(n_61), .B(n_59), .CI(n_76));
  ADDFX1 g1580(.CO(n_81), .S(n_82), .A(n_24), .B(n_50), .CI(n_64));
  ADDFX1 g1581(.CO(n_79), .S(n_80), .A(n_21), .B(n_15), .CI(n_43));
  ADDFX1 g1582(.CO(n_77), .S(n_78), .A(n_32), .B(n_38), .CI(n_40));
  ADDFX1 g1583(.CO(n_75), .S(n_76), .A(n_47), .B(n_51), .CI(n_55));
  ADDFX1 g1584(.CO(n_73), .S(n_74), .A(n_18), .B(n_46), .CI(n_36));
  ADDFX1 g1585(.CO(n_71), .S(n_72), .A(in_30[1]), .B(n_41), .CI(n_39));
  ADDFX1 g1586(.CO(n_69), .S(n_70), .A(n_22), .B(n_52), .CI(n_44));
  ADDFX1 g1587(.CO(n_67), .S(n_68), .A(n_35), .B(n_48), .CI(n_34));
  ADDFX1 g1588(.CO(n_65), .S(n_66), .A(n_16), .B(n_49), .CI(n_26));
  ADDFX1 g1589(.CO(n_63), .S(n_64), .A(in_5[0]), .B(n_20), .CI(n_42));
  ADDFX1 g1590(.CO(n_61), .S(n_62), .A(n_31), .B(n_45), .CI(n_37));
  ADDFX1 g1591(.CO(n_59), .S(n_60), .A(n_23), .B(n_17), .CI(n_19));
  ADDFX1 g1592(.CO(n_57), .S(n_58), .A(in_40[0]), .B(n_8), .CI(n_33));
  NOR2X1 g1594(.Y(n_56), .A(in_40[0]), .B(n_54));
  INVX1 g1595(.Y(n_55), .A(n_53));
  ADDFX1 g1596(.CO(n_54), .S(n_53), .A(in_20[0]), .B(in_21[0]), .CI(in_37[0]));
  ADDFX1 g1597(.CO(n_51), .S(n_52), .A(in_3[1]), .B(n_3), .CI(in_41[1]));
  ADDFX1 g1598(.CO(n_49), .S(n_50), .A(in_9[0]), .B(in_12[0]), .CI(in_13[0]));
  ADDFX1 g1599(.CO(n_47), .S(n_48), .A(in_18[1]), .B(n_12), .CI(in_36[0]));
  ADDFX1 g1600(.CO(n_45), .S(n_46), .A(in_15[0]), .B(n_10), .CI(in_21[0]));
  ADDFX1 g1601(.CO(n_43), .S(n_44), .A(in_7[1]), .B(in_8[0]), .CI(n_7));
  INVX1 g1602(.Y(n_42), .A(n_30));
  INVX1 g1603(.Y(n_41), .A(n_29));
  INVX1 g1604(.Y(n_40), .A(n_28));
  INVX1 g1605(.Y(n_39), .A(n_27));
  ADDFX1 g1606(.CO(n_37), .S(n_38), .A(in_14[0]), .B(in_20[0]), .CI(n_4));
  ADDFX1 g1607(.CO(n_35), .S(n_36), .A(in_17[0]), .B(in_22[0]), .CI(in_36[0]));
  ADDFX1 g1608(.CO(n_33), .S(n_34), .A(in_15[0]), .B(in_17[0]), .CI(in_34[1]));
  ADDFX1 g1609(.CO(n_31), .S(n_32), .A(n_9), .B(n_13), .CI(in_40[0]));
  ADDFX1 g1610(.CO(n_29), .S(n_30), .A(in_2[0]), .B(in_10[0]), .CI(in_11[0]));
  ADDFX1 g1611(.CO(n_27), .S(n_28), .A(in_0[0]), .B(in_23[0]), .CI(in_25[0]));
  ADDFX1 g1612(.CO(n_25), .S(n_26), .A(in_32[1]), .B(n_11), .CI(in_5[1]));
  ADDFX1 g1613(.CO(n_23), .S(n_24), .A(in_16[0]), .B(in_37[0]), .CI(in_39[0]));
  ADDFX1 g1614(.CO(n_21), .S(n_22), .A(in_22[0]), .B(in_19[1]), .CI(n_14));
  ADDFX1 g1615(.CO(n_19), .S(n_20), .A(in_8[0]), .B(in_27[0]), .CI(n_6));
  ADDFX1 g1616(.CO(n_17), .S(n_18), .A(in_29[0]), .B(n_2), .CI(in_44[0]));
  ADDFX1 g1617(.CO(n_15), .S(n_16), .A(in_39[0]), .B(in_42[1]), .CI(n_5));
  INVX1 g1618(.Y(n_14), .A(in_31[1]));
  INVX1 g1619(.Y(n_13), .A(in_38[0]));
  INVX1 g1620(.Y(n_12), .A(in_4[1]));
  INVX1 g1621(.Y(n_11), .A(in_13[1]));
  INVX1 g1622(.Y(n_10), .A(in_1[0]));
  INVX1 g1623(.Y(n_9), .A(in_26[0]));
  INVX1 g1624(.Y(n_8), .A(in_30[1]));
  INVX1 g1626(.Y(n_7), .A(in_35[1]));
  INVX1 g1627(.Y(n_6), .A(in_28[0]));
  INVX1 g1628(.Y(n_5), .A(in_43[1]));
  INVX1 g1629(.Y(n_4), .A(in_24[0]));
  INVX1 g1630(.Y(n_3), .A(in_6[1]));
  INVX1 g1631(.Y(n_2), .A(in_33[0]));
  CLKXOR2X1 g2(.Y(n_0), .A(in_40[0]), .B(n_54));
endmodule

module WALLACE_CSA_DUMMY_OP850_group_359289(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, out_0);
input  in_24, in_27, in_29, in_37, in_38, in_46, in_49;
input   [4:0] in_0;
input   [4:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [1:0] in_18;
input   [1:0] in_19;
input   [4:0] in_20;
input   [3:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [1:0] in_25;
input   [1:0] in_26;
input   [1:0] in_28;
input   [1:0] in_30;
input   [2:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [1:0] in_39;
input   [4:0] in_40;
input   [2:0] in_41;
input   [1:0] in_42;
input   [4:0] in_43;
input   [1:0] in_44;
input   [4:0] in_45;
input   [1:0] in_47;
input   [1:0] in_48;
output  [9:0] out_0;
wire  n_136, n_133, n_131, n_129, n_128, n_127, n_126, n_125, n_124, n_123, 
    n_122, n_121, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, 
    n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, in_49, in_46, in_38, in_37, in_29, in_27, in_24;
wire   [9:0] out_0;
wire   [2:0] in_41;
wire   [2:0] in_31;
wire   [3:0] in_21;
wire   [1:0] in_48;
wire   [1:0] in_47;
wire   [1:0] in_44;
wire   [1:0] in_42;
wire   [1:0] in_39;
wire   [1:0] in_36;
wire   [1:0] in_30;
wire   [1:0] in_28;
wire   [1:0] in_26;
wire   [1:0] in_25;
wire   [1:0] in_19;
wire   [1:0] in_18;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [4:0] in_45;
wire   [4:0] in_43;
wire   [4:0] in_40;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  AO21X1 g1693(.Y(out_0[6]), .A0(n_115), .A1(n_136), .B0(out_0[9]));
  NOR2X1 g1694(.Y(out_0[9]), .A(n_115), .B(n_136));
  ADDFX1 g1695(.CO(n_136), .S(out_0[5]), .A(n_118), .B(n_125), .CI(n_133));
  ADDFX1 g1696(.CO(n_133), .S(out_0[4]), .A(n_126), .B(n_127), .CI(n_131));
  ADDFX1 g1697(.CO(n_131), .S(out_0[3]), .A(n_121), .B(n_128), .CI(n_129));
  ADDFX1 g1698(.CO(n_129), .S(out_0[2]), .A(n_117), .B(n_122), .CI(n_119));
  ADDFX1 g1699(.CO(n_127), .S(n_128), .A(n_107), .B(n_116), .CI(n_124));
  ADDFX1 g1700(.CO(n_125), .S(n_126), .A(n_113), .B(n_111), .CI(n_123));
  ADDFX1 g1701(.CO(n_123), .S(n_124), .A(n_103), .B(n_98), .CI(n_112));
  ADDFX1 g1702(.CO(n_121), .S(n_122), .A(n_108), .B(n_105), .CI(n_109));
  ADDFX1 g1703(.CO(n_119), .S(out_0[1]), .A(n_95), .B(n_110), .CI(n_106));
  AOI2BB1X1 g1704(.Y(n_118), .A0N(n_54), .A1N(n_114), .B0(n_115));
  ADDFX1 g1705(.CO(n_116), .S(n_117), .A(n_91), .B(n_102), .CI(n_104));
  AND2X1 g1706(.Y(n_115), .A(n_114), .B(n_54));
  ADDFX1 g1707(.CO(n_114), .S(n_113), .A(n_53), .B(n_99), .CI(n_97));
  ADDFX1 g1708(.CO(n_111), .S(n_112), .A(n_85), .B(n_100), .CI(n_101));
  ADDFX1 g1709(.CO(n_109), .S(n_110), .A(n_81), .B(n_94), .CI(n_92));
  ADDFX1 g1710(.CO(n_107), .S(n_108), .A(n_73), .B(n_86), .CI(n_93));
  ADDFX1 g1711(.CO(n_105), .S(n_106), .A(n_76), .B(n_74), .CI(n_90));
  ADDFX1 g1712(.CO(n_103), .S(n_104), .A(n_75), .B(n_62), .CI(n_88));
  ADDFX1 g1713(.CO(n_101), .S(n_102), .A(n_68), .B(n_84), .CI(n_89));
  ADDFX1 g1714(.CO(n_99), .S(n_100), .A(n_53), .B(n_71), .CI(n_87));
  ADDFX1 g1715(.CO(n_97), .S(n_98), .A(n_67), .B(n_61), .CI(n_83));
  ADDFX1 g1716(.CO(n_95), .S(out_0[0]), .A(n_56), .B(n_80), .CI(n_82));
  ADDFX1 g1717(.CO(n_93), .S(n_94), .A(n_55), .B(n_59), .CI(n_66));
  ADDFX1 g1718(.CO(n_91), .S(n_92), .A(n_79), .B(n_78), .CI(n_58));
  ADDFX1 g1719(.CO(n_89), .S(n_90), .A(n_46), .B(n_28), .CI(n_64));
  ADDFX1 g1720(.CO(n_87), .S(n_88), .A(n_27), .B(n_29), .CI(n_63));
  ADDFX1 g1721(.CO(n_85), .S(n_86), .A(n_77), .B(n_57), .CI(n_65));
  ADDFX1 g1722(.CO(n_83), .S(n_84), .A(n_8), .B(in_31[2]), .CI(n_72));
  ADDFX1 g1723(.CO(n_81), .S(n_82), .A(n_34), .B(n_36), .CI(n_60));
  ADDFX1 g1724(.CO(n_79), .S(n_80), .A(n_44), .B(n_48), .CI(n_38));
  ADDFX1 g1725(.CO(n_77), .S(n_78), .A(n_47), .B(n_41), .CI(n_37));
  ADDFX1 g1726(.CO(n_75), .S(n_76), .A(n_30), .B(n_26), .CI(n_16));
  ADDFX1 g1727(.CO(n_73), .S(n_74), .A(n_32), .B(n_40), .CI(n_35));
  INVX1 g1728(.Y(n_72), .A(n_70));
  INVX1 g1729(.Y(n_71), .A(n_69));
  ADDFX1 g1730(.CO(n_69), .S(n_70), .A(in_2[2]), .B(in_45[0]), .CI(n_49));
  ADDFX1 g1731(.CO(n_67), .S(n_68), .A(n_15), .B(n_25), .CI(n_31));
  ADDFX1 g1732(.CO(n_65), .S(n_66), .A(n_33), .B(n_21), .CI(n_43));
  ADDFX1 g1733(.CO(n_63), .S(n_64), .A(in_28[0]), .B(in_30[1]), .CI(n_51));
  ADDFX1 g1734(.CO(n_61), .S(n_62), .A(n_45), .B(n_52), .CI(n_39));
  ADDFX1 g1735(.CO(n_59), .S(n_60), .A(n_18), .B(n_42), .CI(n_20));
  ADDFX1 g1736(.CO(n_57), .S(n_58), .A(n_19), .B(n_17), .CI(n_23));
  ADDFX1 g1737(.CO(n_55), .S(n_56), .A(in_9[0]), .B(n_22), .CI(n_24));
  INVX1 g1738(.Y(n_53), .A(n_54));
  ADDFX1 g1739(.CO(n_54), .S(n_52), .A(in_8[2]), .B(n_14), .CI(in_21[2]));
  INVX1 g1740(.Y(n_51), .A(n_50));
  ADDFX1 g1741(.CO(n_49), .S(n_50), .A(in_13[1]), .B(in_3[1]), .CI(in_15[1]));
  ADDFX1 g1742(.CO(n_47), .S(n_48), .A(in_5[0]), .B(in_19[0]), .CI(n_6));
  ADDFX1 g1743(.CO(n_45), .S(n_46), .A(n_13), .B(n_7), .CI(in_36[0]));
  ADDFX1 g1744(.CO(n_43), .S(n_44), .A(in_12[0]), .B(in_6[0]), .CI(in_42[0]));
  ADDFX1 g1745(.CO(n_41), .S(n_42), .A(in_26[0]), .B(n_12), .CI(in_44[0]));
  ADDFX1 g1746(.CO(n_39), .S(n_40), .A(in_10[1]), .B(in_9[1]), .CI(n_3));
  ADDFX1 g1747(.CO(n_37), .S(n_38), .A(in_13[0]), .B(n_11), .CI(in_36[0]));
  ADDFX1 g1748(.CO(n_35), .S(n_36), .A(in_4[0]), .B(in_49), .CI(in_7[0]));
  ADDFX1 g1749(.CO(n_33), .S(n_34), .A(in_18[0]), .B(in_47[0]), .CI(n_2));
  ADDFX1 g1750(.CO(n_31), .S(n_32), .A(in_5[1]), .B(in_11[1]), .CI(in_25[1]));
  ADDFX1 g1751(.CO(n_29), .S(n_30), .A(in_4[0]), .B(in_18[0]), .CI(in_41[1]));
  ADDFX1 g1752(.CO(n_27), .S(n_28), .A(n_4), .B(n_5), .CI(in_48[1]));
  ADDFX1 g1753(.CO(n_25), .S(n_26), .A(in_12[1]), .B(in_47[0]), .CI(in_26[0]));
  ADDFX1 g1754(.CO(n_23), .S(n_24), .A(in_45[0]), .B(in_38), .CI(in_46));
  ADDFX1 g1755(.CO(n_21), .S(n_22), .A(in_14[0]), .B(n_10), .CI(in_37));
  ADDFX1 g1756(.CO(n_19), .S(n_20), .A(in_17[0]), .B(in_24), .CI(in_28[0]));
  ADDFX1 g1757(.CO(n_17), .S(n_18), .A(in_27), .B(n_1), .CI(in_29));
  ADDFX1 g1758(.CO(n_15), .S(n_16), .A(in_39[1]), .B(in_19[0]), .CI(n_9));
  INVX1 g1759(.Y(n_14), .A(in_32[2]));
  INVX1 g1760(.Y(n_13), .A(in_23[1]));
  INVX1 g1761(.Y(n_12), .A(in_43[0]));
  INVX1 g1762(.Y(n_11), .A(in_0[0]));
  INVX1 g1763(.Y(n_10), .A(in_33[0]));
  INVX1 g1764(.Y(n_9), .A(in_34[1]));
  INVX1 g1765(.Y(n_8), .A(in_17[0]));
  INVX1 g1766(.Y(n_7), .A(in_40[1]));
  INVX1 g1767(.Y(n_6), .A(in_35[0]));
  INVX1 g1768(.Y(n_5), .A(in_16[1]));
  INVX1 g1769(.Y(n_4), .A(in_1[1]));
  INVX1 g1770(.Y(n_3), .A(in_7[1]));
  INVX1 g1771(.Y(n_2), .A(in_20[0]));
  INVX1 g1772(.Y(n_1), .A(in_22[0]));
endmodule

module WALLACE_CSA_DUMMY_OP875_group_359275(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, out_0);
input  in_26, in_27, in_33;
input   [4:0] in_0;
input   [4:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [4:0] in_4;
input   [4:0] in_5;
input   [4:0] in_6;
input   [4:0] in_7;
input   [4:0] in_8;
input   [4:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [1:0] in_28;
input   [4:0] in_29;
input   [2:0] in_30;
input   [4:0] in_31;
input   [2:0] in_32;
input   [4:0] in_34;
output  [9:0] out_0;
wire  n_104, n_102, n_100, n_98, n_97, n_96, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_82, n_81, n_80, n_79, n_78, n_77, n_76, 
    n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, 
    n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, 
    n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
    n_1, in_33, in_27, in_26;
wire   [9:0] out_0;
wire   [2:0] in_32;
wire   [2:0] in_30;
wire   [1:0] in_28;
wire   [1:0] in_25;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [4:0] in_34;
wire   [4:0] in_31;
wire   [4:0] in_29;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_9;
wire   [4:0] in_8;
wire   [4:0] in_7;
wire   [4:0] in_6;
wire   [4:0] in_5;
wire   [4:0] in_4;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1363(.Y(out_0[9]), .A(n_104));
  ADDFX1 g1364(.CO(n_104), .S(out_0[5]), .A(n_12), .B(n_92), .CI(n_102));
  ADDFX1 g1365(.CO(n_102), .S(out_0[4]), .A(n_93), .B(n_96), .CI(n_100));
  ADDFX1 g1366(.CO(n_100), .S(out_0[3]), .A(n_97), .B(n_90), .CI(n_98));
  ADDFX1 g1367(.CO(n_98), .S(out_0[2]), .A(n_84), .B(n_94), .CI(n_91));
  ADDFX1 g1368(.CO(n_96), .S(n_97), .A(n_80), .B(n_89), .CI(n_86));
  ADDFX1 g1369(.CO(n_94), .S(out_0[1]), .A(n_79), .B(n_82), .CI(n_85));
  ADDFX1 g1370(.CO(n_92), .S(n_93), .A(n_14), .B(n_70), .CI(n_88));
  ADDFX1 g1371(.CO(n_90), .S(n_91), .A(n_78), .B(n_81), .CI(n_87));
  ADDFX1 g1372(.CO(n_88), .S(n_89), .A(n_66), .B(n_71), .CI(n_76));
  ADDFX1 g1373(.CO(n_86), .S(n_87), .A(n_68), .B(n_74), .CI(n_77));
  ADDFX1 g1374(.CO(n_84), .S(n_85), .A(n_72), .B(n_69), .CI(n_75));
  ADDFX1 g1375(.CO(n_82), .S(out_0[0]), .A(n_53), .B(n_55), .CI(n_73));
  ADDFX1 g1376(.CO(n_80), .S(n_81), .A(n_58), .B(n_63), .CI(n_67));
  ADDFX1 g1377(.CO(n_78), .S(n_79), .A(n_52), .B(n_59), .CI(n_61));
  ADDFX1 g1378(.CO(n_76), .S(n_77), .A(n_48), .B(n_60), .CI(n_64));
  ADDFX1 g1379(.CO(n_74), .S(n_75), .A(n_49), .B(n_54), .CI(n_65));
  ADDFX1 g1380(.CO(n_72), .S(n_73), .A(n_20), .B(n_18), .CI(n_57));
  ADDFX1 g1381(.CO(n_70), .S(n_71), .A(n_14), .B(n_46), .CI(n_62));
  ADDFX1 g1382(.CO(n_68), .S(n_69), .A(n_17), .B(n_38), .CI(n_56));
  ADDFX1 g1383(.CO(n_66), .S(n_67), .A(n_21), .B(n_37), .CI(n_47));
  ADDFX1 g1384(.CO(n_64), .S(n_65), .A(n_30), .B(n_41), .CI(n_51));
  ADDFX1 g1385(.CO(n_62), .S(n_63), .A(in_32[2]), .B(n_23), .CI(n_50));
  ADDFX1 g1386(.CO(n_60), .S(n_61), .A(n_32), .B(n_15), .CI(n_34));
  ADDFX1 g1387(.CO(n_58), .S(n_59), .A(n_39), .B(n_24), .CI(n_22));
  ADDFX1 g1388(.CO(n_56), .S(n_57), .A(in_20[0]), .B(in_22[0]), .CI(n_43));
  ADDFX1 g1389(.CO(n_54), .S(n_55), .A(n_42), .B(n_31), .CI(n_16));
  ADDFX1 g1390(.CO(n_52), .S(n_53), .A(n_29), .B(n_40), .CI(n_33));
  ADDFX1 g1391(.CO(n_50), .S(n_51), .A(in_10[1]), .B(n_13), .CI(n_26));
  ADDFX1 g1392(.CO(n_48), .S(n_49), .A(n_9), .B(n_19), .CI(n_28));
  INVX1 g1393(.Y(n_47), .A(n_45));
  INVX1 g1394(.Y(n_46), .A(n_44));
  ADDFX1 g1395(.CO(n_44), .S(n_45), .A(in_24[2]), .B(in_34[0]), .CI(n_12));
  OAI21X1 g1396(.Y(n_43), .A0(in_8[0]), .A1(n_27), .B0(n_34));
  ADDFX1 g1397(.CO(n_41), .S(n_42), .A(in_10[0]), .B(in_17[0]), .CI(n_6));
  ADDFX1 g1398(.CO(n_39), .S(n_40), .A(in_12[0]), .B(in_27), .CI(in_18[0]));
  INVX1 g1399(.Y(n_38), .A(n_36));
  INVX1 g1400(.Y(n_37), .A(n_35));
  ADDFX1 g1401(.CO(n_35), .S(n_36), .A(in_19[1]), .B(in_22[1]), .CI(in_20[1]));
  NAND2X1 g1402(.Y(n_34), .A(in_8[0]), .B(n_27));
  ADDFX1 g1403(.CO(n_32), .S(n_33), .A(n_8), .B(n_7), .CI(in_15[0]));
  ADDFX1 g1404(.CO(n_30), .S(n_31), .A(n_10), .B(n_4), .CI(in_33));
  ADDFX1 g1405(.CO(n_28), .S(n_29), .A(in_28[0]), .B(n_3), .CI(in_34[0]));
  INVX1 g1406(.Y(n_26), .A(n_25));
  ADDFX1 g1407(.CO(n_25), .S(n_27), .A(in_2[0]), .B(in_3[0]), .CI(in_13[0]));
  ADDFX1 g1408(.CO(n_23), .S(n_24), .A(in_14[0]), .B(in_11[1]), .CI(in_30[1]));
  ADDFX1 g1409(.CO(n_21), .S(n_22), .A(in_12[1]), .B(n_11), .CI(in_16[1]));
  ADDFX1 g1410(.CO(n_19), .S(n_20), .A(in_16[0]), .B(in_26), .CI(n_2));
  ADDFX1 g1411(.CO(n_17), .S(n_18), .A(in_25[0]), .B(in_21[0]), .CI(in_19[0]));
  ADDFX1 g1412(.CO(n_15), .S(n_16), .A(in_14[0]), .B(n_1), .CI(n_5));
  INVX1 g1413(.Y(n_14), .A(n_12));
  XOR2XL g1414(.Y(n_13), .A(in_15[1]), .B(in_17[1]));
  NOR2X1 g1415(.Y(n_12), .A(in_17[1]), .B(in_15[1]));
  INVX1 g1416(.Y(n_11), .A(in_5[1]));
  INVX1 g1417(.Y(n_10), .A(in_1[0]));
  INVX1 g1418(.Y(n_9), .A(in_21[1]));
  INVX1 g1419(.Y(n_8), .A(in_0[0]));
  INVX1 g1420(.Y(n_7), .A(in_6[0]));
  INVX1 g1421(.Y(n_6), .A(in_31[0]));
  INVX1 g1422(.Y(n_5), .A(in_29[0]));
  INVX1 g1423(.Y(n_4), .A(in_4[0]));
  INVX1 g1424(.Y(n_3), .A(in_9[0]));
  INVX1 g1425(.Y(n_2), .A(in_7[0]));
  INVX1 g1426(.Y(n_1), .A(in_23[0]));
endmodule

module WALLACE_CSA_DUMMY_OP1315_group_109833(in_0, in_1, in_2, in_3, in_4, in_5
    , in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, out_0);
input  in_24, in_36, in_38, in_41;
input   [1:0] in_0;
input   [1:0] in_1;
input   [4:0] in_2;
input   [4:0] in_3;
input   [2:0] in_4;
input   [4:0] in_5;
input   [4:0] in_6;
input   [9:0] in_7;
input   [5:0] in_8;
input   [4:0] in_9;
input   [1:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [1:0] in_25;
input   [4:0] in_26;
input   [2:0] in_27;
input   [4:0] in_28;
input   [2:0] in_29;
input   [1:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [2:0] in_35;
input   [1:0] in_37;
input   [1:0] in_39;
input   [1:0] in_40;
input   [1:0] in_42;
output  [9:0] out_0;
wire  n_132, n_130, n_128, n_126, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_41, in_38, 
    in_36, in_24;
wire   [9:0] out_0;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_8;
wire   [9:0] in_7;
wire   [2:0] in_35;
wire   [2:0] in_29;
wire   [2:0] in_27;
wire   [2:0] in_4;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_28;
wire   [4:0] in_26;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_9;
wire   [4:0] in_6;
wire   [4:0] in_5;
wire   [4:0] in_3;
wire   [4:0] in_2;
wire   [1:0] in_42;
wire   [1:0] in_40;
wire   [1:0] in_39;
wire   [1:0] in_37;
wire   [1:0] in_31;
wire   [1:0] in_30;
wire   [1:0] in_25;
wire   [1:0] in_10;
wire   [1:0] in_1;
wire   [1:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  INVX1 g4054(.Y(out_0[9]), .A(n_132));
  ADDFX1 g4055(.CO(n_132), .S(out_0[6]), .A(n_18), .B(n_110), .CI(n_130));
  ADDFX1 g4056(.CO(n_130), .S(out_0[5]), .A(n_111), .B(n_120), .CI(n_128));
  ADDFX1 g4057(.CO(n_128), .S(out_0[4]), .A(n_122), .B(n_121), .CI(n_126));
  ADDFX1 g4058(.CO(n_126), .S(out_0[3]), .A(n_118), .B(n_123), .CI(n_124));
  ADDFX1 g4059(.CO(n_124), .S(out_0[2]), .A(n_119), .B(n_116), .CI(n_113));
  ADDFX1 g4060(.CO(n_122), .S(n_123), .A(n_115), .B(n_105), .CI(n_112));
  ADDFX1 g4061(.CO(n_120), .S(n_121), .A(n_114), .B(n_104), .CI(n_108));
  ADDFX1 g4062(.CO(n_118), .S(n_119), .A(n_103), .B(n_106), .CI(n_94));
  ADDFX1 g4063(.CO(n_116), .S(out_0[1]), .A(n_107), .B(n_98), .CI(n_95));
  ADDFX1 g4064(.CO(n_114), .S(n_115), .A(n_97), .B(n_100), .CI(n_102));
  ADDFX1 g4065(.CO(n_112), .S(n_113), .A(n_92), .B(n_101), .CI(in_7[2]));
  OAI2BB1X1 g4066(.Y(n_111), .A0N(in_7[5]), .A1N(n_109), .B0(n_110));
  OR2X1 g4067(.Y(n_110), .A(in_7[5]), .B(n_109));
  ADDFX1 g4068(.CO(n_109), .S(n_108), .A(n_78), .B(n_96), .CI(in_7[4]));
  ADDFX1 g4069(.CO(n_106), .S(n_107), .A(n_89), .B(n_85), .CI(n_93));
  ADDFX1 g4070(.CO(n_104), .S(n_105), .A(n_86), .B(n_90), .CI(in_7[3]));
  ADDFX1 g4071(.CO(n_102), .S(n_103), .A(n_87), .B(n_84), .CI(n_91));
  ADDFX1 g4072(.CO(n_100), .S(n_101), .A(n_81), .B(n_56), .CI(n_88));
  ADDFX1 g4073(.CO(n_98), .S(out_0[0]), .A(n_71), .B(n_83), .CI(in_7[0]));
  ADDFX1 g4074(.CO(n_96), .S(n_97), .A(n_64), .B(n_79), .CI(n_80));
  ADDFX1 g4075(.CO(n_94), .S(n_95), .A(n_57), .B(n_82), .CI(in_7[1]));
  ADDFX1 g4076(.CO(n_92), .S(n_93), .A(n_62), .B(n_67), .CI(n_77));
  ADDFX1 g4077(.CO(n_90), .S(n_91), .A(n_65), .B(n_66), .CI(n_76));
  ADDFX1 g4078(.CO(n_88), .S(n_89), .A(n_37), .B(n_61), .CI(n_70));
  ADDFX1 g4079(.CO(n_86), .S(n_87), .A(n_74), .B(n_60), .CI(n_59));
  ADDFX1 g4080(.CO(n_84), .S(n_85), .A(n_69), .B(n_75), .CI(n_72));
  ADDFX1 g4081(.CO(n_82), .S(n_83), .A(n_46), .B(n_63), .CI(n_73));
  ADDFX1 g4082(.CO(n_80), .S(n_81), .A(n_55), .B(n_27), .CI(n_68));
  ADDHX1 g4083(.CO(n_78), .S(n_79), .A(n_54), .B(n_58));
  ADDFX1 g4084(.CO(n_76), .S(n_77), .A(n_53), .B(n_44), .CI(n_24));
  ADDFX1 g4085(.CO(n_74), .S(n_75), .A(n_7), .B(n_47), .CI(n_49));
  ADDFX1 g4086(.CO(n_72), .S(n_73), .A(n_50), .B(n_36), .CI(n_48));
  ADDFX1 g4087(.CO(n_70), .S(n_71), .A(n_40), .B(n_34), .CI(n_52));
  ADDFX1 g4088(.CO(n_68), .S(n_69), .A(n_19), .B(n_41), .CI(n_51));
  ADDFX1 g4089(.CO(n_66), .S(n_67), .A(n_21), .B(n_32), .CI(n_26));
  ADDFX1 g4090(.CO(n_64), .S(n_65), .A(n_20), .B(n_29), .CI(n_31));
  ADDFX1 g4091(.CO(n_62), .S(n_63), .A(n_22), .B(n_42), .CI(n_38));
  ADDFX1 g4092(.CO(n_60), .S(n_61), .A(n_39), .B(n_33), .CI(n_35));
  ADDFX1 g4093(.CO(n_58), .S(n_59), .A(n_43), .B(n_23), .CI(n_25));
  ADDFX1 g4094(.CO(n_56), .S(n_57), .A(n_30), .B(n_45), .CI(n_28));
  INVX1 g4095(.Y(n_55), .A(n_54));
  ADDFX1 g4096(.CO(n_54), .S(n_53), .A(in_25[1]), .B(in_37[1]), .CI(in_21[0]));
  ADDFX1 g4097(.CO(n_51), .S(n_52), .A(n_5), .B(in_42[0]), .CI(n_3));
  ADDFX1 g4098(.CO(n_49), .S(n_50), .A(in_1[0]), .B(n_13), .CI(in_39[0]));
  ADDFX1 g4099(.CO(n_47), .S(n_48), .A(in_17[0]), .B(n_6), .CI(n_17));
  ADDFX1 g4100(.CO(n_45), .S(n_46), .A(in_12[0]), .B(in_16[0]), .CI(in_8[0]));
  ADDFX1 g4101(.CO(n_43), .S(n_44), .A(n_4), .B(n_12), .CI(in_29[0]));
  ADDFX1 g4102(.CO(n_41), .S(n_42), .A(in_13[0]), .B(n_11), .CI(in_41));
  ADDFX1 g4103(.CO(n_39), .S(n_40), .A(in_10[0]), .B(n_16), .CI(in_36));
  ADDFX1 g4104(.CO(n_37), .S(n_38), .A(in_15[0]), .B(in_24), .CI(in_19[0]));
  ADDFX1 g4105(.CO(n_35), .S(n_36), .A(in_18[0]), .B(n_2), .CI(in_21[0]));
  ADDFX1 g4106(.CO(n_33), .S(n_34), .A(in_11[0]), .B(in_35[0]), .CI(in_38));
  ADDFX1 g4107(.CO(n_31), .S(n_32), .A(n_14), .B(n_10), .CI(in_40[1]));
  ADDFX1 g4108(.CO(n_29), .S(n_30), .A(in_1[0]), .B(in_17[1]), .CI(n_8));
  ADDFX1 g4109(.CO(n_27), .S(n_28), .A(in_19[1]), .B(n_9), .CI(n_15));
  ADDFX1 g4110(.CO(n_25), .S(n_26), .A(in_27[1]), .B(in_4[1]), .CI(in_30[1]));
  ADDFX1 g4111(.CO(n_23), .S(n_24), .A(in_31[1]), .B(in_15[0]), .CI(in_35[0]));
  OAI21X1 g4112(.Y(n_22), .A0(in_23[0]), .A1(n_1), .B0(n_19));
  OAI2BB1X1 g4113(.Y(n_21), .A0N(in_0[1]), .A1N(in_39[0]), .B0(n_20));
  OR2X1 g4114(.Y(n_20), .A(in_0[1]), .B(in_39[0]));
  NAND2X1 g4115(.Y(n_19), .A(in_23[0]), .B(n_1));
  INVX1 g4116(.Y(n_18), .A(in_7[6]));
  INVX1 g4117(.Y(n_17), .A(in_34[0]));
  INVX1 g4118(.Y(n_16), .A(in_5[0]));
  INVX1 g4119(.Y(n_15), .A(in_12[1]));
  INVX1 g4120(.Y(n_14), .A(in_32[1]));
  INVX1 g4121(.Y(n_13), .A(in_14[0]));
  INVX1 g4122(.Y(n_12), .A(in_22[1]));
  INVX1 g4123(.Y(n_11), .A(in_20[0]));
  INVX1 g4124(.Y(n_10), .A(in_33[1]));
  INVX1 g4125(.Y(n_9), .A(in_16[1]));
  INVX1 g4126(.Y(n_8), .A(in_26[1]));
  INVX1 g4127(.Y(n_7), .A(in_8[1]));
  INVX1 g4128(.Y(n_6), .A(in_2[0]));
  INVX1 g4129(.Y(n_5), .A(in_9[0]));
  INVX1 g4130(.Y(n_4), .A(in_6[1]));
  INVX1 g4131(.Y(n_3), .A(in_28[0]));
  INVX1 g4132(.Y(n_2), .A(in_3[0]));
  INVX1 g4133(.Y(n_1), .A(in_29[0]));
endmodule

module WALLACE_CSA_DUMMY_OP1318_group_109815(in_0, in_1, in_2, in_3, in_4, in_5
    , in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, out_0);
input  in_2, in_37;
input   [3:0] in_0;
input   [2:0] in_1;
input   [4:0] in_3;
input   [4:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [4:0] in_8;
input   [4:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [4:0] in_18;
input   [4:0] in_19;
input   [1:0] in_20;
input   [1:0] in_21;
input   [1:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [2:0] in_25;
input   [3:0] in_26;
input   [4:0] in_27;
input   [2:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [2:0] in_38;
input   [1:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [1:0] in_42;
input   [2:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [2:0] in_46;
output  [9:0] out_0;
wire  n_134, n_132, n_130, n_128, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, 
    n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, 
    n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, 
    n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, 
    n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, 
    n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, 
    n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, 
    n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, 
    in_37, in_2;
wire   [9:0] out_0;
wire   [1:0] in_45;
wire   [1:0] in_42;
wire   [1:0] in_39;
wire   [1:0] in_31;
wire   [1:0] in_22;
wire   [1:0] in_21;
wire   [1:0] in_20;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [4:0] in_44;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_27;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_19;
wire   [4:0] in_18;
wire   [4:0] in_9;
wire   [4:0] in_8;
wire   [4:0] in_4;
wire   [4:0] in_3;
wire   [2:0] in_46;
wire   [2:0] in_43;
wire   [2:0] in_38;
wire   [2:0] in_28;
wire   [2:0] in_25;
wire   [2:0] in_1;
wire   [3:0] in_26;
wire   [3:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g4120(.Y(out_0[9]), .A(n_134));
  ADDFX1 g4121(.CO(n_134), .S(out_0[5]), .A(n_108), .B(n_120), .CI(n_132));
  ADDFX1 g4122(.CO(n_132), .S(out_0[4]), .A(n_121), .B(n_124), .CI(n_130));
  ADDFX1 g4123(.CO(n_130), .S(out_0[3]), .A(n_122), .B(n_125), .CI(n_128));
  ADDFX1 g4124(.CO(n_128), .S(out_0[2]), .A(n_115), .B(n_126), .CI(n_123));
  ADDFX1 g4125(.CO(n_126), .S(out_0[1]), .A(n_105), .B(n_106), .CI(n_117));
  ADDFX1 g4126(.CO(n_124), .S(n_125), .A(n_111), .B(n_114), .CI(n_119));
  ADDFX1 g4127(.CO(n_122), .S(n_123), .A(n_104), .B(n_113), .CI(n_116));
  ADDFX1 g4128(.CO(n_120), .S(n_121), .A(n_109), .B(n_110), .CI(n_118));
  ADDFX1 g4129(.CO(n_118), .S(n_119), .A(n_102), .B(n_100), .CI(n_112));
  ADDFX1 g4130(.CO(n_116), .S(n_117), .A(n_90), .B(n_99), .CI(n_97));
  ADDFX1 g4131(.CO(n_114), .S(n_115), .A(n_98), .B(n_103), .CI(n_101));
  ADDFX1 g4132(.CO(n_112), .S(n_113), .A(n_82), .B(n_95), .CI(n_96));
  ADDFX1 g4133(.CO(n_110), .S(n_111), .A(n_87), .B(n_94), .CI(n_93));
  ADDFX1 g4134(.CO(n_108), .S(n_109), .A(n_44), .B(n_86), .CI(n_92));
  ADDFX1 g4135(.CO(n_106), .S(out_0[0]), .A(n_79), .B(n_81), .CI(n_91));
  ADDFX1 g4136(.CO(n_104), .S(n_105), .A(n_85), .B(n_89), .CI(n_83));
  ADDFX1 g4137(.CO(n_102), .S(n_103), .A(n_64), .B(n_67), .CI(n_88));
  ADDFX1 g4138(.CO(n_100), .S(n_101), .A(n_71), .B(n_84), .CI(n_75));
  ADDFX1 g4139(.CO(n_98), .S(n_99), .A(n_80), .B(n_77), .CI(n_78));
  ADDFX1 g4140(.CO(n_96), .S(n_97), .A(n_69), .B(n_65), .CI(n_72));
  ADDFX1 g4141(.CO(n_94), .S(n_95), .A(n_62), .B(n_76), .CI(n_68));
  ADDFX1 g4142(.CO(n_92), .S(n_93), .A(n_70), .B(n_66), .CI(n_74));
  ADDFX1 g4143(.CO(n_90), .S(n_91), .A(n_46), .B(n_48), .CI(n_73));
  ADDFX1 g4144(.CO(n_88), .S(n_89), .A(n_57), .B(n_30), .CI(n_32));
  ADDFX1 g4145(.CO(n_86), .S(n_87), .A(n_55), .B(n_61), .CI(n_63));
  ADDFX1 g4146(.CO(n_84), .S(n_85), .A(n_52), .B(n_42), .CI(n_33));
  ADDFX1 g4147(.CO(n_82), .S(n_83), .A(n_28), .B(n_38), .CI(n_47));
  ADDFX1 g4148(.CO(n_80), .S(n_81), .A(n_36), .B(n_54), .CI(n_34));
  ADDFX1 g4149(.CO(n_78), .S(n_79), .A(n_21), .B(n_40), .CI(n_50));
  ADDFX1 g4150(.CO(n_76), .S(n_77), .A(n_20), .B(n_49), .CI(n_45));
  ADDFX1 g4151(.CO(n_74), .S(n_75), .A(n_56), .B(n_24), .CI(n_37));
  ADDFX1 g4152(.CO(n_72), .S(n_73), .A(n_58), .B(n_23), .CI(n_26));
  ADDFX1 g4153(.CO(n_70), .S(n_71), .A(in_1[1]), .B(n_51), .CI(n_31));
  ADDFX1 g4154(.CO(n_68), .S(n_69), .A(n_1), .B(n_53), .CI(n_39));
  ADDFX1 g4155(.CO(n_66), .S(n_67), .A(n_41), .B(n_27), .CI(n_29));
  ADDFX1 g4156(.CO(n_64), .S(n_65), .A(n_22), .B(n_25), .CI(n_35));
  OAI2BB1X1 g4157(.Y(n_63), .A0N(n_9), .A1N(n_43), .B0(n_44));
  INVX1 g4158(.Y(n_62), .A(n_60));
  INVX1 g4159(.Y(n_61), .A(n_59));
  ADDFX1 g4160(.CO(n_59), .S(n_60), .A(in_9[0]), .B(in_33[0]), .CI(in_40[0]));
  ADDFX1 g4161(.CO(n_57), .S(n_58), .A(in_19[0]), .B(in_42[0]), .CI(in_43[0]));
  ADDFX1 g4162(.CO(n_55), .S(n_56), .A(n_10), .B(n_2), .CI(in_46[0]));
  ADDFX1 g4163(.CO(n_53), .S(n_54), .A(in_33[0]), .B(n_14), .CI(in_40[0]));
  ADDFX1 g4164(.CO(n_51), .S(n_52), .A(in_16[1]), .B(in_25[1]), .CI(n_17));
  ADDFX1 g4165(.CO(n_49), .S(n_50), .A(in_32[0]), .B(n_12), .CI(in_46[0]));
  ADDFX1 g4166(.CO(n_47), .S(n_48), .A(in_1[0]), .B(in_5[0]), .CI(in_14[0]));
  ADDFX1 g4167(.CO(n_45), .S(n_46), .A(in_18[0]), .B(in_22[0]), .CI(n_5));
  OR2X1 g4168(.Y(n_44), .A(n_9), .B(n_43));
  ADDFX1 g4169(.CO(n_41), .S(n_42), .A(n_3), .B(n_7), .CI(in_45[0]));
  ADDFX1 g4170(.CO(n_39), .S(n_40), .A(in_9[0]), .B(in_6[0]), .CI(in_37));
  ADDFX1 g4171(.CO(n_37), .S(n_38), .A(in_28[1]), .B(in_5[1]), .CI(n_15));
  ADDFX1 g4172(.CO(n_35), .S(n_36), .A(in_11[0]), .B(n_4), .CI(n_19));
  ADDFX1 g4173(.CO(n_33), .S(n_34), .A(in_12[0]), .B(in_39[0]), .CI(in_2));
  ADDFX1 g4174(.CO(n_31), .S(n_32), .A(in_20[1]), .B(n_16), .CI(in_43[0]));
  ADDFX1 g4175(.CO(n_29), .S(n_30), .A(in_7[1]), .B(in_10[1]), .CI(n_18));
  ADDFX1 g4176(.CO(n_27), .S(n_28), .A(in_21[1]), .B(n_13), .CI(in_32[0]));
  ADDFX1 g4177(.CO(n_25), .S(n_26), .A(in_15[0]), .B(in_8[0]), .CI(in_45[0]));
  ADDFX1 g4178(.CO(n_43), .S(n_24), .A(in_26[2]), .B(in_38[2]), .CI(n_11));
  ADDFX1 g4179(.CO(n_22), .S(n_23), .A(in_31[0]), .B(n_6), .CI(n_8));
  OAI2BB1X1 g4180(.Y(n_21), .A0N(in_17[0]), .A1N(in_16[0]), .B0(n_20));
  OR2X1 g4181(.Y(n_20), .A(in_17[0]), .B(in_16[0]));
  INVX1 g4182(.Y(n_19), .A(in_13[0]));
  INVX1 g4183(.Y(n_18), .A(in_41[1]));
  INVX1 g4184(.Y(n_17), .A(in_36[1]));
  INVX1 g4185(.Y(n_16), .A(in_29[1]));
  INVX1 g4186(.Y(n_15), .A(in_14[1]));
  INVX1 g4187(.Y(n_14), .A(in_30[0]));
  INVX1 g4188(.Y(n_13), .A(in_23[1]));
  INVX1 g4189(.Y(n_12), .A(in_34[0]));
  INVX1 g4190(.Y(n_11), .A(in_8[0]));
  INVX1 g4191(.Y(n_10), .A(in_18[0]));
  INVX1 g4192(.Y(n_9), .A(in_32[0]));
  INVX1 g4193(.Y(n_8), .A(in_44[0]));
  INVX1 g4194(.Y(n_7), .A(in_24[1]));
  INVX1 g4195(.Y(n_6), .A(in_35[0]));
  INVX1 g4196(.Y(n_5), .A(in_4[0]));
  INVX1 g4197(.Y(n_4), .A(in_3[0]));
  INVX1 g4198(.Y(n_3), .A(in_27[1]));
  INVX1 g4199(.Y(n_2), .A(in_19[0]));
  INVX1 g4200(.Y(n_1), .A(in_1[1]));
endmodule

module WALLACE_CSA_DUMMY_OP_group_109839_6286_6339(in_0, in_1, in_2, in_3, in_4
    , in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, 
    in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26
    , in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, 
    in_37, in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47
    , in_48, in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, 
    in_58, in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, out_0);
input  in_60;
input   [4:0] in_0;
input   [4:0] in_1;
input   [2:0] in_2;
input   [4:0] in_3;
input   [9:0] in_4;
input   [8:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [4:0] in_19;
input   [2:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [4:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [4:0] in_49;
input   [2:0] in_50;
input   [4:0] in_51;
input   [1:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [2:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [1:0] in_59;
input   [4:0] in_61;
input   [2:0] in_62;
input   [1:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
output  [9:0] out_0;
wire  n_244, n_241, n_239, n_237, n_236, n_235, n_234, n_233, n_231, n_230, 
    n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, 
    n_219, n_218, n_217, n_216, n_214, n_213, n_212, n_211, n_210, n_209, 
    n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_199, n_198, 
    n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, 
    n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, 
    n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, 
    n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, in_60;
wire   [9:0] out_0;
wire   [1:0] in_63;
wire   [1:0] in_59;
wire   [1:0] in_52;
wire   [1:0] in_37;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [8:0] in_5;
wire   [9:0] in_4;
wire   [2:0] in_62;
wire   [2:0] in_56;
wire   [2:0] in_50;
wire   [2:0] in_20;
wire   [2:0] in_2;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_61;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_51;
wire   [4:0] in_49;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_23;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_19;
wire   [4:0] in_3;
wire   [4:0] in_1;
wire   [4:0] in_0;
  assign out_0[8] = 1'b0;
  OA21X1 g7127(.Y(out_0[7]), .A0(n_213), .A1(n_244), .B0(out_0[9]));
  NAND2X1 g7128(.Y(out_0[9]), .A(n_213), .B(n_244));
  ADDFX1 g7129(.CO(n_244), .S(out_0[6]), .A(n_218), .B(n_229), .CI(n_241));
  ADDFX1 g7130(.CO(n_241), .S(out_0[5]), .A(n_235), .B(n_230), .CI(n_239));
  ADDFX1 g7131(.CO(n_239), .S(out_0[4]), .A(n_233), .B(n_236), .CI(n_237));
  ADDFX1 g7132(.CO(n_237), .S(out_0[3]), .A(n_223), .B(n_234), .CI(n_231));
  ADDFX1 g7133(.CO(n_235), .S(n_236), .A(n_217), .B(n_225), .CI(n_228));
  ADDFX1 g7134(.CO(n_233), .S(n_234), .A(n_219), .B(n_209), .CI(n_226));
  ADDFX1 g7135(.CO(n_231), .S(out_0[2]), .A(n_220), .B(n_214), .CI(n_224));
  ADDFX1 g7136(.CO(n_229), .S(n_230), .A(n_216), .B(n_211), .CI(n_227));
  ADDFX1 g7137(.CO(n_227), .S(n_228), .A(n_221), .B(n_196), .CI(n_207));
  ADDFX1 g7138(.CO(n_225), .S(n_226), .A(n_198), .B(n_222), .CI(n_208));
  ADDFX1 g7139(.CO(n_223), .S(n_224), .A(n_190), .B(n_203), .CI(n_210));
  ADDFX1 g7140(.CO(n_221), .S(n_222), .A(n_189), .B(n_205), .CI(n_187));
  ADDFX1 g7141(.CO(n_219), .S(n_220), .A(n_206), .B(n_185), .CI(n_201));
  OAI2BB1X1 g7142(.Y(n_218), .A0N(n_182), .A1N(n_212), .B0(n_213));
  ADDFX1 g7143(.CO(n_216), .S(n_217), .A(n_197), .B(n_194), .CI(n_191));
  ADDFX1 g7144(.CO(n_214), .S(out_0[1]), .A(n_199), .B(n_202), .CI(n_204));
  OR2X1 g7145(.Y(n_213), .A(n_182), .B(n_212));
  ADDFX1 g7146(.CO(n_212), .S(n_211), .A(n_193), .B(n_195), .CI(n_163));
  ADDFX1 g7147(.CO(n_209), .S(n_210), .A(n_188), .B(n_180), .CI(n_175));
  ADDFX1 g7148(.CO(n_207), .S(n_208), .A(n_184), .B(n_174), .CI(n_192));
  ADDFX1 g7149(.CO(n_205), .S(n_206), .A(n_160), .B(n_172), .CI(n_157));
  ADDFX1 g7150(.CO(n_203), .S(n_204), .A(n_173), .B(n_181), .CI(n_186));
  ADDFX1 g7151(.CO(n_201), .S(n_202), .A(n_171), .B(n_178), .CI(n_152));
  ADDFX1 g7152(.CO(n_199), .S(out_0[0]), .A(n_131), .B(n_179), .CI(n_153));
  ADDFX1 g7153(.CO(n_197), .S(n_198), .A(n_166), .B(n_176), .CI(n_162));
  ADDFX1 g7154(.CO(n_195), .S(n_196), .A(n_161), .B(n_183), .CI(in_4[4]));
  ADDFX1 g7155(.CO(n_193), .S(n_194), .A(n_124), .B(n_164), .CI(n_154));
  ADDFX1 g7156(.CO(n_191), .S(n_192), .A(n_165), .B(n_168), .CI(in_4[3]));
  ADDFX1 g7157(.CO(n_189), .S(n_190), .A(n_167), .B(n_177), .CI(n_170));
  ADDFX1 g7158(.CO(n_187), .S(n_188), .A(n_137), .B(n_169), .CI(n_150));
  ADDFX1 g7159(.CO(n_185), .S(n_186), .A(n_115), .B(n_158), .CI(n_151));
  ADDFX1 g7160(.CO(n_183), .S(n_184), .A(n_136), .B(n_159), .CI(in_5[3]));
  AOI21X1 g7161(.Y(n_182), .A0(n_36), .A1(in_4[5]), .B0(n_156));
  ADDFX1 g7162(.CO(n_180), .S(n_181), .A(n_145), .B(n_139), .CI(in_4[1]));
  ADDFX1 g7163(.CO(n_178), .S(n_179), .A(n_149), .B(n_141), .CI(n_129));
  ADDFX1 g7164(.CO(n_176), .S(n_177), .A(n_116), .B(n_135), .CI(n_146));
  ADDFX1 g7165(.CO(n_174), .S(n_175), .A(n_144), .B(n_114), .CI(in_4[2]));
  ADDFX1 g7166(.CO(n_172), .S(n_173), .A(n_130), .B(n_143), .CI(n_148));
  ADDFX1 g7167(.CO(n_170), .S(n_171), .A(n_120), .B(n_140), .CI(n_147));
  ADDFX1 g7168(.CO(n_168), .S(n_169), .A(n_142), .B(n_126), .CI(in_5[2]));
  ADDFX1 g7169(.CO(n_166), .S(n_167), .A(n_133), .B(n_113), .CI(n_138));
  ADDFX1 g7170(.CO(n_164), .S(n_165), .A(n_110), .B(n_132), .CI(n_134));
  AO21XL g7171(.Y(n_163), .A0(n_155), .A1(n_47), .B0(n_156));
  ADDFX1 g7172(.CO(n_161), .S(n_162), .A(n_109), .B(n_112), .CI(n_125));
  ADDFX1 g7173(.CO(n_159), .S(n_160), .A(n_118), .B(n_89), .CI(n_111));
  ADDFX1 g7174(.CO(n_157), .S(n_158), .A(n_117), .B(n_127), .CI(n_128));
  NOR2X1 g7175(.Y(n_156), .A(n_155), .B(n_47));
  ADDFX1 g7176(.CO(n_155), .S(n_154), .A(n_36), .B(n_108), .CI(n_20));
  ADDFX1 g7177(.CO(n_152), .S(n_153), .A(n_57), .B(n_121), .CI(in_4[0]));
  ADDFX1 g7178(.CO(n_150), .S(n_151), .A(n_119), .B(n_90), .CI(in_5[1]));
  ADDFX1 g7179(.CO(n_148), .S(n_149), .A(n_98), .B(n_73), .CI(n_61));
  ADDFX1 g7180(.CO(n_146), .S(n_147), .A(n_81), .B(n_107), .CI(n_83));
  ADDFX1 g7181(.CO(n_144), .S(n_145), .A(n_92), .B(n_87), .CI(n_96));
  ADDFX1 g7182(.CO(n_142), .S(n_143), .A(n_58), .B(n_62), .CI(n_99));
  ADDFX1 g7183(.CO(n_140), .S(n_141), .A(n_46), .B(n_71), .CI(n_100));
  ADDFX1 g7184(.CO(n_138), .S(n_139), .A(n_52), .B(n_69), .CI(n_75));
  ADDFX1 g7185(.CO(n_136), .S(n_137), .A(n_88), .B(n_76), .CI(n_103));
  ADDFX1 g7186(.CO(n_134), .S(n_135), .A(n_86), .B(n_95), .CI(n_91));
  ADDFX1 g7187(.CO(n_132), .S(n_133), .A(n_37), .B(n_68), .CI(n_106));
  ADDFX1 g7188(.CO(n_130), .S(n_131), .A(n_63), .B(n_65), .CI(n_79));
  ADDFX1 g7189(.CO(n_128), .S(n_129), .A(n_53), .B(n_85), .CI(in_5[0]));
  ADDFX1 g7190(.CO(n_126), .S(n_127), .A(n_72), .B(n_78), .CI(n_44));
  INVX1 g7191(.Y(n_125), .A(n_123));
  INVX1 g7192(.Y(n_124), .A(n_122));
  ADDFX1 g7193(.CO(n_122), .S(n_123), .A(n_54), .B(n_43), .CI(n_101));
  ADDFX1 g7194(.CO(n_120), .S(n_121), .A(in_18[0]), .B(n_67), .CI(n_59));
  ADDFX1 g7195(.CO(n_118), .S(n_119), .A(n_97), .B(n_84), .CI(n_66));
  ADDFX1 g7196(.CO(n_116), .S(n_117), .A(n_60), .B(n_64), .CI(n_70));
  ADDFX1 g7197(.CO(n_114), .S(n_115), .A(n_42), .B(n_56), .CI(n_77));
  ADDFX1 g7198(.CO(n_112), .S(n_113), .A(n_82), .B(n_74), .CI(n_45));
  ADDFX1 g7199(.CO(n_110), .S(n_111), .A(in_10[2]), .B(n_0), .CI(n_80));
  ADDFX1 g7200(.CO(n_108), .S(n_109), .A(n_35), .B(n_3), .CI(n_39));
  INVX1 g7201(.Y(n_107), .A(n_105));
  INVX1 g7202(.Y(n_106), .A(n_104));
  ADDFX1 g7203(.CO(n_104), .S(n_105), .A(in_44[1]), .B(in_29[1]), .CI(in_48[1]));
  INVX1 g7204(.Y(n_103), .A(n_102));
  ADDFX1 g7205(.CO(n_101), .S(n_102), .A(in_8[2]), .B(in_11[2]), .CI(in_15[2]));
  ADDFX1 g7206(.CO(n_99), .S(n_100), .A(in_40[0]), .B(in_14[0]), .CI(n_32));
  ADDFX1 g7207(.CO(n_97), .S(n_98), .A(n_19), .B(n_28), .CI(in_60));
  INVX1 g7208(.Y(n_96), .A(n_94));
  INVX1 g7209(.Y(n_95), .A(n_93));
  ADDFX1 g7210(.CO(n_93), .S(n_94), .A(in_54[1]), .B(in_14[1]), .CI(in_57[1]));
  ADDFX1 g7211(.CO(n_91), .S(n_92), .A(in_28[0]), .B(n_31), .CI(in_56[0]));
  ADDFX1 g7212(.CO(n_89), .S(n_90), .A(in_15[1]), .B(n_5), .CI(in_11[1]));
  INVX1 g7213(.Y(n_88), .A(n_55));
  INVX1 g7214(.Y(n_87), .A(n_51));
  INVX1 g7215(.Y(n_86), .A(n_50));
  INVX1 g7216(.Y(n_85), .A(n_49));
  INVX1 g7217(.Y(n_84), .A(n_48));
  ADDFX1 g7218(.CO(n_82), .S(n_83), .A(in_2[1]), .B(in_10[0]), .CI(n_12));
  ADDFX1 g7219(.CO(n_80), .S(n_81), .A(in_22[0]), .B(n_25), .CI(in_62[1]));
  ADDFX1 g7220(.CO(n_78), .S(n_79), .A(in_22[0]), .B(n_21), .CI(n_13));
  ADDFX1 g7221(.CO(n_76), .S(n_77), .A(n_9), .B(in_8[1]), .CI(n_30));
  ADDFX1 g7222(.CO(n_74), .S(n_75), .A(in_20[1]), .B(n_24), .CI(in_59[1]));
  ADDFX1 g7223(.CO(n_72), .S(n_73), .A(in_36[0]), .B(n_6), .CI(in_63[0]));
  ADDFX1 g7224(.CO(n_70), .S(n_71), .A(in_28[0]), .B(n_10), .CI(in_65[0]));
  ADDFX1 g7225(.CO(n_68), .S(n_69), .A(n_7), .B(n_2), .CI(in_50[0]));
  ADDFX1 g7226(.CO(n_66), .S(n_67), .A(in_9[0]), .B(n_23), .CI(in_42[0]));
  ADDFX1 g7227(.CO(n_64), .S(n_65), .A(n_26), .B(n_17), .CI(in_52[0]));
  ADDFX1 g7228(.CO(n_62), .S(n_63), .A(in_15[0]), .B(n_27), .CI(n_29));
  ADDFX1 g7229(.CO(n_60), .S(n_61), .A(n_4), .B(n_8), .CI(in_56[0]));
  ADDFX1 g7230(.CO(n_58), .S(n_59), .A(n_11), .B(n_18), .CI(in_37[0]));
  ADDFX1 g7231(.CO(n_56), .S(n_57), .A(in_8[0]), .B(in_12[0]), .CI(in_16[0]));
  ADDFX1 g7232(.CO(n_54), .S(n_55), .A(in_35[0]), .B(in_42[0]), .CI(in_65[0]));
  ADDFX1 g7233(.CO(n_52), .S(n_53), .A(in_10[0]), .B(n_22), .CI(in_50[0]));
  ADDFX1 g7234(.CO(n_50), .S(n_51), .A(in_46[1]), .B(in_23[1]), .CI(in_47[1]));
  ADDFX1 g7235(.CO(n_48), .S(n_49), .A(in_38[0]), .B(in_41[0]), .CI(in_51[0]));
  XNOR2X1 g7236(.Y(n_47), .A(n_36), .B(in_4[5]));
  XNOR2X1 g7237(.Y(n_46), .A(in_19[0]), .B(n_40));
  XNOR2X1 g7238(.Y(n_45), .A(in_31[0]), .B(n_41));
  OAI21X1 g7239(.Y(n_44), .A0(n_16), .A1(n_38), .B0(n_34));
  AOI21X1 g7240(.Y(n_43), .A0(n_15), .A1(n_34), .B0(n_38));
  OAI2BB1X1 g7241(.Y(n_42), .A0N(in_7[1]), .A1N(n_33), .B0(n_37));
  MX2XL g7242(.Y(n_41), .A(in_36[0]), .B(n_15), .S0(in_19[0]));
  MX2XL g7244(.Y(n_40), .A(n_16), .B(in_35[0]), .S0(in_31[0]));
  OAI22XL g7245(.Y(n_39), .A0(in_28[0]), .A1(n_14), .B0(in_22[0]), .B1(n_1));
  NOR2X1 g7246(.Y(n_38), .A(in_19[0]), .B(in_31[0]));
  OR2X1 g7247(.Y(n_37), .A(in_7[1]), .B(n_33));
  NAND2X1 g7248(.Y(n_36), .A(n_1), .B(n_14));
  NOR2X1 g7249(.Y(n_35), .A(in_61[2]), .B(in_40[0]));
  NAND2X1 g7250(.Y(n_34), .A(in_31[0]), .B(in_19[0]));
  INVX1 g7251(.Y(n_33), .A(in_66[1]));
  INVX1 g7252(.Y(n_32), .A(in_55[0]));
  INVX1 g7253(.Y(n_31), .A(in_64[1]));
  INVX1 g7254(.Y(n_30), .A(in_18[1]));
  INVX1 g7255(.Y(n_29), .A(in_34[0]));
  INVX1 g7256(.Y(n_28), .A(in_53[0]));
  INVX1 g7257(.Y(n_27), .A(in_25[0]));
  INVX1 g7258(.Y(n_26), .A(in_1[0]));
  INVX1 g7259(.Y(n_25), .A(in_43[1]));
  INVX1 g7260(.Y(n_24), .A(in_27[1]));
  INVX1 g7261(.Y(n_23), .A(in_26[0]));
  INVX1 g7262(.Y(n_22), .A(in_21[0]));
  INVX1 g7263(.Y(n_21), .A(in_0[0]));
  INVX1 g7264(.Y(n_20), .A(in_5[4]));
  INVX1 g7265(.Y(n_19), .A(in_13[0]));
  INVX1 g7266(.Y(n_18), .A(in_32[0]));
  INVX1 g7267(.Y(n_17), .A(in_17[0]));
  INVX1 g7268(.Y(n_16), .A(in_35[0]));
  INVX1 g7269(.Y(n_15), .A(in_36[0]));
  INVX1 g7270(.Y(n_14), .A(in_22[0]));
  INVX1 g7271(.Y(n_13), .A(in_24[0]));
  INVX1 g7272(.Y(n_12), .A(in_58[1]));
  INVX1 g7273(.Y(n_11), .A(in_6[0]));
  INVX1 g7274(.Y(n_10), .A(in_30[0]));
  INVX1 g7275(.Y(n_9), .A(in_16[1]));
  INVX1 g7276(.Y(n_8), .A(in_33[0]));
  INVX1 g7277(.Y(n_7), .A(in_3[1]));
  INVX1 g7278(.Y(n_6), .A(in_49[0]));
  INVX1 g7279(.Y(n_5), .A(in_12[1]));
  INVX1 g7280(.Y(n_4), .A(in_39[0]));
  INVX1 g7281(.Y(n_3), .A(in_10[3]));
  INVX1 g7282(.Y(n_2), .A(in_45[1]));
  INVX1 g7284(.Y(n_1), .A(in_28[0]));
  CLKXOR2X1 g2(.Y(n_0), .A(in_40[0]), .B(in_61[2]));
endmodule

module WALLACE_CSA_DUMMY_OP_group_109839(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, out_0);
input  in_34, in_35, in_37, in_38;
input   [1:0] in_0;
input   [1:0] in_1;
input   [6:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [4:0] in_9;
input   [1:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [1:0] in_14;
input   [1:0] in_15;
input   [4:0] in_16;
input   [4:0] in_17;
input   [2:0] in_18;
input   [4:0] in_19;
input   [2:0] in_20;
input   [4:0] in_21;
input   [1:0] in_22;
input   [1:0] in_23;
input   [4:0] in_24;
input   [4:0] in_25;
input   [2:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [4:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [3:0] in_32;
input   [4:0] in_33;
input   [4:0] in_36;
output  [9:0] out_0;
wire  n_111, n_109, n_107, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_38, in_37, 
    in_35, in_34;
wire   [9:0] out_0;
wire   [3:0] in_32;
wire   [2:0] in_26;
wire   [2:0] in_20;
wire   [2:0] in_18;
wire   [4:0] in_36;
wire   [4:0] in_33;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_29;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_25;
wire   [4:0] in_24;
wire   [4:0] in_21;
wire   [4:0] in_19;
wire   [4:0] in_17;
wire   [4:0] in_16;
wire   [4:0] in_9;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [6:0] in_2;
wire   [1:0] in_23;
wire   [1:0] in_22;
wire   [1:0] in_15;
wire   [1:0] in_14;
wire   [1:0] in_10;
wire   [1:0] in_1;
wire   [1:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1355(.Y(out_0[9]), .A(n_111));
  ADDFX1 g1356(.CO(n_111), .S(out_0[5]), .A(n_54), .B(n_101), .CI(n_109));
  ADDFX1 g1357(.CO(n_109), .S(out_0[4]), .A(n_102), .B(n_103), .CI(n_107));
  ADDFX1 g1358(.CO(n_107), .S(out_0[3]), .A(n_99), .B(n_105), .CI(n_104));
  ADDFX1 g1359(.CO(n_105), .S(out_0[2]), .A(n_94), .B(n_97), .CI(n_100));
  ADDFX1 g1360(.CO(n_103), .S(n_104), .A(n_85), .B(n_93), .CI(n_96));
  ADDFX1 g1361(.CO(n_101), .S(n_102), .A(n_72), .B(n_89), .CI(n_95));
  ADDFX1 g1362(.CO(n_99), .S(n_100), .A(n_84), .B(n_86), .CI(n_91));
  ADDFX1 g1363(.CO(n_97), .S(out_0[1]), .A(n_81), .B(n_88), .CI(n_92));
  ADDFX1 g1364(.CO(n_95), .S(n_96), .A(n_77), .B(n_83), .CI(n_90));
  ADDFX1 g1365(.CO(n_93), .S(n_94), .A(n_78), .B(n_79), .CI(n_87));
  ADDFX1 g1366(.CO(n_91), .S(n_92), .A(n_64), .B(n_71), .CI(n_80));
  ADDFX1 g1367(.CO(n_89), .S(n_90), .A(n_75), .B(n_66), .CI(n_61));
  ADDFX1 g1368(.CO(n_87), .S(n_88), .A(n_69), .B(n_57), .CI(n_74));
  ADDFX1 g1369(.CO(n_85), .S(n_86), .A(n_68), .B(n_73), .CI(n_70));
  ADDFX1 g1370(.CO(n_83), .S(n_84), .A(n_67), .B(n_59), .CI(n_76));
  ADDFX1 g1371(.CO(n_81), .S(out_0[0]), .A(n_58), .B(n_63), .CI(n_65));
  ADDFX1 g1372(.CO(n_79), .S(n_80), .A(n_56), .B(n_60), .CI(n_62));
  ADDFX1 g1373(.CO(n_77), .S(n_78), .A(n_49), .B(n_55), .CI(n_53));
  ADDFX1 g1374(.CO(n_75), .S(n_76), .A(n_37), .B(n_47), .CI(n_7));
  ADDFX1 g1375(.CO(n_73), .S(n_74), .A(n_38), .B(n_36), .CI(n_48));
  INVX1 g1376(.Y(n_72), .A(n_54));
  ADDFX1 g1377(.CO(n_70), .S(n_71), .A(n_46), .B(n_33), .CI(n_50));
  ADDFX1 g1378(.CO(n_68), .S(n_69), .A(n_31), .B(n_39), .CI(n_42));
  ADDFX1 g1379(.CO(n_66), .S(n_67), .A(n_41), .B(n_45), .CI(n_35));
  ADDFX1 g1380(.CO(n_64), .S(n_65), .A(n_28), .B(n_22), .CI(n_34));
  ADDFX1 g1381(.CO(n_62), .S(n_63), .A(n_40), .B(n_24), .CI(n_32));
  OAI21X1 g1382(.Y(n_61), .A0(n_19), .A1(n_52), .B0(n_54));
  ADDFX1 g1383(.CO(n_59), .S(n_60), .A(n_21), .B(n_23), .CI(in_2[1]));
  ADDFX1 g1384(.CO(n_57), .S(n_58), .A(n_30), .B(n_44), .CI(n_26));
  ADDFX1 g1385(.CO(n_55), .S(n_56), .A(n_25), .B(n_29), .CI(n_27));
  NAND2X1 g1386(.Y(n_54), .A(n_19), .B(n_52));
  INVX1 g1387(.Y(n_53), .A(n_51));
  ADDFX1 g1388(.CO(n_52), .S(n_51), .A(in_31[0]), .B(in_6[2]), .CI(n_20));
  ADDFX1 g1389(.CO(n_49), .S(n_50), .A(in_6[1]), .B(n_12), .CI(n_43));
  ADDFX1 g1390(.CO(n_47), .S(n_48), .A(n_9), .B(in_26[0]), .CI(n_18));
  ADDFX1 g1391(.CO(n_45), .S(n_46), .A(in_0[1]), .B(in_3[1]), .CI(n_4));
  ADDFX1 g1392(.CO(n_43), .S(n_44), .A(n_2), .B(in_11[0]), .CI(in_37));
  ADDFX1 g1393(.CO(n_41), .S(n_42), .A(in_18[1]), .B(n_10), .CI(in_20[0]));
  ADDFX1 g1394(.CO(n_39), .S(n_40), .A(in_7[0]), .B(in_12[0]), .CI(n_5));
  ADDFX1 g1395(.CO(n_37), .S(n_38), .A(in_14[1]), .B(in_15[1]), .CI(n_15));
  ADDFX1 g1396(.CO(n_35), .S(n_36), .A(in_1[1]), .B(n_3), .CI(n_13));
  ADDFX1 g1397(.CO(n_33), .S(n_34), .A(in_5[0]), .B(in_6[0]), .CI(in_4[0]));
  ADDFX1 g1398(.CO(n_31), .S(n_32), .A(n_1), .B(n_8), .CI(in_31[0]));
  ADDFX1 g1399(.CO(n_29), .S(n_30), .A(in_2[0]), .B(in_22[0]), .CI(n_14));
  ADDFX1 g1400(.CO(n_27), .S(n_28), .A(in_8[0]), .B(in_26[0]), .CI(in_38));
  ADDFX1 g1401(.CO(n_25), .S(n_26), .A(in_13[0]), .B(n_11), .CI(in_34));
  ADDFX1 g1402(.CO(n_23), .S(n_24), .A(n_6), .B(in_35), .CI(in_20[0]));
  ADDFX1 g1403(.CO(n_21), .S(n_22), .A(in_10[0]), .B(in_23[0]), .CI(n_16));
  XNOR2X1 g1404(.Y(n_20), .A(in_32[2]), .B(n_17));
  NAND2X1 g1405(.Y(n_19), .A(in_32[2]), .B(n_17));
  XNOR2X1 g1406(.Y(n_18), .A(in_13[1]), .B(in_11[0]));
  NAND2X1 g1407(.Y(n_17), .A(in_13[1]), .B(in_11[0]));
  INVX1 g1408(.Y(n_16), .A(in_33[0]));
  INVX1 g1409(.Y(n_15), .A(in_28[1]));
  INVX1 g1410(.Y(n_14), .A(in_30[0]));
  INVX1 g1411(.Y(n_13), .A(in_4[1]));
  INVX1 g1412(.Y(n_12), .A(in_5[1]));
  INVX1 g1413(.Y(n_11), .A(in_24[0]));
  INVX1 g1414(.Y(n_10), .A(in_17[1]));
  INVX1 g1415(.Y(n_9), .A(in_9[1]));
  INVX1 g1416(.Y(n_8), .A(in_19[0]));
  INVX1 g1417(.Y(n_7), .A(in_2[2]));
  INVX1 g1418(.Y(n_6), .A(in_21[0]));
  INVX1 g1419(.Y(n_5), .A(in_16[0]));
  INVX1 g1420(.Y(n_4), .A(in_36[1]));
  INVX1 g1421(.Y(n_3), .A(in_29[1]));
  INVX1 g1422(.Y(n_2), .A(in_27[0]));
  INVX1 g1423(.Y(n_1), .A(in_25[0]));
endmodule

module WALLACE_CSA_DUMMY_OP_group_109839_6286(in_0, in_1, in_2, in_3, in_4, in_5
    , in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27
    , in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, 
    in_38, in_39, in_40, in_41, in_42, in_43, in_44, in_45, in_46, in_47, in_48
    , in_49, in_50, in_51, in_52, in_53, in_54, in_55, in_56, in_57, in_58, 
    in_59, in_60, in_61, in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69
    , in_70, in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, 
    in_80, in_81, in_82, in_83, in_84, out_0);
input  in_42, in_43, in_50, in_68, in_71, in_78, in_79, in_81;
input   [5:0] in_0;
input   [4:0] in_1;
input   [9:0] in_2;
input   [9:0] in_3;
input   [6:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [5:0] in_32;
input   [5:0] in_33;
input   [5:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [4:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [3:0] in_40;
input   [4:0] in_41;
input   [4:0] in_44;
input   [4:0] in_45;
input   [4:0] in_46;
input   [4:0] in_47;
input   [4:0] in_48;
input   [2:0] in_49;
input   [4:0] in_51;
input   [4:0] in_52;
input   [4:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [4:0] in_56;
input   [1:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [1:0] in_60;
input   [1:0] in_61;
input   [4:0] in_62;
input   [1:0] in_63;
input   [4:0] in_64;
input   [4:0] in_65;
input   [2:0] in_66;
input   [1:0] in_67;
input   [4:0] in_69;
input   [4:0] in_70;
input   [2:0] in_72;
input   [1:0] in_73;
input   [1:0] in_74;
input   [2:0] in_75;
input   [4:0] in_76;
input   [2:0] in_77;
input   [1:0] in_80;
input   [1:0] in_82;
input   [2:0] in_83;
input   [4:0] in_84;
output  [9:0] out_0;
wire  n_278, n_276, n_274, n_272, n_270, n_269, n_268, n_267, n_266, n_264, 
    n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
    n_253, n_252, n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, 
    n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
    n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
    n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, 
    n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_204, n_203, n_202, 
    n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, 
    n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
    n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, 
    n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, 
    n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
    n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, 
    n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, 
    n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, 
    n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
    n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, 
    n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, 
    n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
    n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_1, n_0, in_81, in_79, in_78, in_71, in_68, in_50, in_43, 
    in_42;
wire   [9:0] out_0;
wire   [1:0] in_82;
wire   [1:0] in_80;
wire   [1:0] in_74;
wire   [1:0] in_73;
wire   [1:0] in_67;
wire   [1:0] in_63;
wire   [1:0] in_61;
wire   [1:0] in_60;
wire   [1:0] in_57;
wire   [3:0] in_40;
wire   [2:0] in_83;
wire   [2:0] in_77;
wire   [2:0] in_75;
wire   [2:0] in_72;
wire   [2:0] in_66;
wire   [2:0] in_49;
wire   [2:0] in_39;
wire   [6:0] in_4;
wire   [9:0] in_3;
wire   [9:0] in_2;
wire   [4:0] in_84;
wire   [4:0] in_76;
wire   [4:0] in_70;
wire   [4:0] in_69;
wire   [4:0] in_65;
wire   [4:0] in_64;
wire   [4:0] in_62;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_56;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_53;
wire   [4:0] in_52;
wire   [4:0] in_51;
wire   [4:0] in_48;
wire   [4:0] in_47;
wire   [4:0] in_46;
wire   [4:0] in_45;
wire   [4:0] in_44;
wire   [4:0] in_41;
wire   [4:0] in_38;
wire   [4:0] in_37;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_1;
wire   [5:0] in_34;
wire   [5:0] in_33;
wire   [5:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g9353(.Y(out_0[9]), .A(n_278));
  ADDFX1 g9354(.CO(n_278), .S(out_0[7]), .A(n_203), .B(n_260), .CI(n_276));
  ADDFX1 g9355(.CO(n_276), .S(out_0[6]), .A(n_261), .B(n_266), .CI(n_274));
  ADDFX1 g9356(.CO(n_274), .S(out_0[5]), .A(n_268), .B(n_267), .CI(n_272));
  ADDFX1 g9357(.CO(n_272), .S(out_0[4]), .A(n_262), .B(n_270), .CI(n_269));
  ADDFX1 g9358(.CO(n_270), .S(out_0[3]), .A(n_255), .B(n_263), .CI(n_264));
  ADDFX1 g9359(.CO(n_268), .S(n_269), .A(n_254), .B(n_247), .CI(n_259));
  ADDFX1 g9360(.CO(n_266), .S(n_267), .A(n_246), .B(n_257), .CI(n_258));
  ADDFX1 g9361(.CO(n_264), .S(out_0[2]), .A(n_253), .B(n_250), .CI(n_237));
  ADDFX1 g9362(.CO(n_262), .S(n_263), .A(n_252), .B(n_249), .CI(n_236));
  ADDFX1 g9363(.CO(n_260), .S(n_261), .A(n_244), .B(n_198), .CI(n_256));
  ADDFX1 g9364(.CO(n_258), .S(n_259), .A(n_248), .B(n_242), .CI(n_241));
  ADDFX1 g9365(.CO(n_256), .S(n_257), .A(n_167), .B(n_240), .CI(n_245));
  ADDFX1 g9366(.CO(n_254), .S(n_255), .A(n_230), .B(n_233), .CI(n_243));
  ADDFX1 g9367(.CO(n_252), .S(n_253), .A(n_231), .B(n_235), .CI(n_238));
  ADDFX1 g9368(.CO(n_250), .S(out_0[1]), .A(n_204), .B(n_207), .CI(n_239));
  ADDFX1 g9369(.CO(n_248), .S(n_249), .A(n_223), .B(n_234), .CI(n_218));
  ADDFX1 g9370(.CO(n_246), .S(n_247), .A(n_222), .B(n_232), .CI(n_229));
  ADDFX1 g9371(.CO(n_244), .S(n_245), .A(n_224), .B(in_2[5]), .CI(n_228));
  ADDFX1 g9372(.CO(n_242), .S(n_243), .A(n_220), .B(n_226), .CI(n_211));
  ADDFX1 g9373(.CO(n_240), .S(n_241), .A(n_208), .B(n_225), .CI(n_210));
  ADDFX1 g9374(.CO(n_238), .S(n_239), .A(n_217), .B(n_215), .CI(n_177));
  ADDFX1 g9375(.CO(n_236), .S(n_237), .A(n_227), .B(n_219), .CI(n_206));
  ADDFX1 g9376(.CO(n_234), .S(n_235), .A(n_216), .B(n_221), .CI(n_214));
  ADDFX1 g9377(.CO(n_232), .S(n_233), .A(n_201), .B(n_212), .CI(n_209));
  ADDFX1 g9378(.CO(n_230), .S(n_231), .A(n_189), .B(n_202), .CI(n_213));
  ADDFX1 g9379(.CO(n_228), .S(n_229), .A(n_199), .B(in_2[4]), .CI(in_3[4]));
  ADDFX1 g9380(.CO(n_226), .S(n_227), .A(n_193), .B(n_165), .CI(in_2[2]));
  ADDFX1 g9381(.CO(n_224), .S(n_225), .A(n_174), .B(n_196), .CI(n_160));
  ADDFX1 g9382(.CO(n_222), .S(n_223), .A(n_197), .B(n_188), .CI(n_200));
  ADDFX1 g9383(.CO(n_220), .S(n_221), .A(n_185), .B(n_180), .CI(n_179));
  ADDFX1 g9384(.CO(n_218), .S(n_219), .A(in_3[2]), .B(n_176), .CI(n_194));
  ADDFX1 g9385(.CO(n_216), .S(n_217), .A(n_169), .B(n_181), .CI(n_186));
  ADDFX1 g9386(.CO(n_214), .S(n_215), .A(n_191), .B(n_171), .CI(n_172));
  ADDFX1 g9387(.CO(n_212), .S(n_213), .A(n_170), .B(n_168), .CI(n_190));
  ADDFX1 g9388(.CO(n_210), .S(n_211), .A(n_192), .B(in_3[3]), .CI(in_2[3]));
  ADDFX1 g9389(.CO(n_208), .S(n_209), .A(n_184), .B(n_175), .CI(n_178));
  ADDFX1 g9390(.CO(n_206), .S(n_207), .A(n_166), .B(n_163), .CI(n_195));
  ADDFX1 g9391(.CO(n_204), .S(out_0[0]), .A(n_187), .B(n_173), .CI(n_164));
  OAI21X1 g9392(.Y(n_203), .A0(n_162), .A1(n_31), .B0(n_27));
  ADDFX1 g9393(.CO(n_201), .S(n_202), .A(n_135), .B(n_138), .CI(n_183));
  ADDFX1 g9394(.CO(n_199), .S(n_200), .A(n_137), .B(n_134), .CI(n_182));
  XOR2XL g9395(.Y(n_198), .A(n_162), .B(n_31));
  ADDFX1 g9396(.CO(n_196), .S(n_197), .A(n_79), .B(n_154), .CI(n_140));
  ADDFX1 g9397(.CO(n_194), .S(n_195), .A(n_139), .B(n_146), .CI(in_2[1]));
  ADDFX1 g9398(.CO(n_192), .S(n_193), .A(n_152), .B(n_112), .CI(n_114));
  ADDFX1 g9399(.CO(n_190), .S(n_191), .A(n_120), .B(n_153), .CI(n_128));
  ADDFX1 g9400(.CO(n_188), .S(n_189), .A(n_155), .B(n_141), .CI(n_156));
  ADDFX1 g9401(.CO(n_186), .S(n_187), .A(n_145), .B(n_129), .CI(n_149));
  ADDFX1 g9402(.CO(n_184), .S(n_185), .A(n_132), .B(n_130), .CI(n_109));
  ADDFX1 g9403(.CO(n_182), .S(n_183), .A(n_122), .B(n_150), .CI(n_118));
  ADDFX1 g9404(.CO(n_180), .S(n_181), .A(n_151), .B(n_131), .CI(n_148));
  ADDFX1 g9405(.CO(n_178), .S(n_179), .A(n_127), .B(n_159), .CI(n_124));
  ADDFX1 g9406(.CO(n_176), .S(n_177), .A(n_115), .B(n_157), .CI(in_3[1]));
  ADDFX1 g9407(.CO(n_174), .S(n_175), .A(n_108), .B(n_158), .CI(n_126));
  ADDFX1 g9408(.CO(n_172), .S(n_173), .A(n_143), .B(n_117), .CI(in_3[0]));
  ADDFX1 g9409(.CO(n_170), .S(n_171), .A(n_133), .B(n_142), .CI(n_116));
  ADDFX1 g9410(.CO(n_168), .S(n_169), .A(n_111), .B(n_123), .CI(n_144));
  AO21X1 g9411(.Y(n_167), .A0(n_161), .A1(in_3[5]), .B0(n_162));
  ADDFX1 g9412(.CO(n_165), .S(n_166), .A(n_119), .B(n_125), .CI(n_113));
  ADDFX1 g9413(.CO(n_163), .S(n_164), .A(n_121), .B(n_147), .CI(in_2[0]));
  NOR2X1 g9414(.Y(n_162), .A(n_161), .B(in_3[5]));
  ADDFX1 g9415(.CO(n_161), .S(n_160), .A(n_13), .B(n_78), .CI(n_136));
  ADDFX1 g9416(.CO(n_158), .S(n_159), .A(n_36), .B(n_76), .CI(n_44));
  ADDFX1 g9417(.CO(n_156), .S(n_157), .A(n_49), .B(n_80), .CI(n_54));
  ADDFX1 g9418(.CO(n_154), .S(n_155), .A(n_106), .B(n_68), .CI(n_52));
  ADDFX1 g9419(.CO(n_152), .S(n_153), .A(n_104), .B(n_38), .CI(n_70));
  ADDFX1 g9420(.CO(n_150), .S(n_151), .A(in_11[1]), .B(n_98), .CI(n_92));
  ADDFX1 g9421(.CO(n_148), .S(n_149), .A(n_47), .B(n_39), .CI(n_101));
  ADDFX1 g9422(.CO(n_146), .S(n_147), .A(n_83), .B(n_55), .CI(n_81));
  ADDFX1 g9423(.CO(n_144), .S(n_145), .A(n_103), .B(n_105), .CI(n_61));
  ADDFX1 g9424(.CO(n_142), .S(n_143), .A(n_85), .B(n_93), .CI(n_99));
  ADDFX1 g9425(.CO(n_140), .S(n_141), .A(n_75), .B(n_89), .CI(n_34));
  ADDFX1 g9426(.CO(n_138), .S(n_139), .A(n_45), .B(n_53), .CI(n_82));
  ADDFX1 g9427(.CO(n_136), .S(n_137), .A(n_74), .B(n_88), .CI(n_72));
  ADDFX1 g9428(.CO(n_134), .S(n_135), .A(n_73), .B(n_48), .CI(n_110));
  ADDFX1 g9429(.CO(n_132), .S(n_133), .A(n_26), .B(n_56), .CI(n_102));
  ADDFX1 g9430(.CO(n_130), .S(n_131), .A(n_32), .B(n_62), .CI(n_84));
  ADDFX1 g9431(.CO(n_128), .S(n_129), .A(n_33), .B(n_59), .CI(n_65));
  ADDFX1 g9432(.CO(n_126), .S(n_127), .A(n_96), .B(n_40), .CI(n_86));
  ADDFX1 g9433(.CO(n_124), .S(n_125), .A(n_87), .B(n_77), .CI(n_97));
  ADDFX1 g9434(.CO(n_122), .S(n_123), .A(n_58), .B(n_100), .CI(n_46));
  ADDFX1 g9435(.CO(n_120), .S(n_121), .A(n_30), .B(n_67), .CI(n_57));
  ADDFX1 g9436(.CO(n_118), .S(n_119), .A(n_64), .B(n_60), .CI(n_66));
  ADDFX1 g9437(.CO(n_116), .S(n_117), .A(n_71), .B(n_43), .CI(n_63));
  ADDFX1 g9438(.CO(n_114), .S(n_115), .A(n_37), .B(n_35), .CI(n_69));
  ADDFX1 g9439(.CO(n_112), .S(n_113), .A(n_42), .B(n_107), .CI(n_41));
  ADDFX1 g9440(.CO(n_110), .S(n_111), .A(n_29), .B(n_4), .CI(in_13[1]));
  ADDFX1 g9441(.CO(n_108), .S(n_109), .A(n_25), .B(n_19), .CI(n_28));
  INVX1 g9442(.Y(n_107), .A(n_95));
  INVX1 g9443(.Y(n_106), .A(n_94));
  INVX1 g9444(.Y(n_105), .A(n_91));
  INVX1 g9445(.Y(n_104), .A(n_90));
  ADDFX1 g9446(.CO(n_102), .S(n_103), .A(in_56[0]), .B(n_8), .CI(in_79));
  ADDFX1 g9447(.CO(n_100), .S(n_101), .A(in_32[0]), .B(in_61[0]), .CI(in_60[0]));
  ADDFX1 g9448(.CO(n_98), .S(n_99), .A(in_7[0]), .B(in_80[0]), .CI(in_21[0]));
  ADDFX1 g9449(.CO(n_96), .S(n_97), .A(in_73[1]), .B(n_11), .CI(n_7));
  ADDFX1 g9450(.CO(n_94), .S(n_95), .A(in_35[1]), .B(in_65[1]), .CI(in_52[1]));
  ADDFX1 g9451(.CO(n_92), .S(n_93), .A(in_24[0]), .B(in_55[0]), .CI(n_21));
  ADDFX1 g9452(.CO(n_90), .S(n_91), .A(in_41[0]), .B(in_46[0]), .CI(in_76[0]));
  ADDFX1 g9453(.CO(n_88), .S(n_89), .A(in_5[2]), .B(in_72[0]), .CI(n_15));
  ADDFX1 g9454(.CO(n_86), .S(n_87), .A(in_39[1]), .B(in_23[1]), .CI(in_83[1]));
  ADDFX1 g9455(.CO(n_84), .S(n_85), .A(in_0[0]), .B(in_30[0]), .CI(in_82[0]));
  ADDFX1 g9456(.CO(n_82), .S(n_83), .A(in_10[0]), .B(in_19[0]), .CI(in_22[0]));
  ADDFX1 g9457(.CO(n_80), .S(n_81), .A(in_4[0]), .B(in_17[0]), .CI(in_26[0]));
  ADDFX1 g9458(.CO(n_78), .S(n_79), .A(n_14), .B(in_55[0]), .CI(n_0));
  ADDFX1 g9459(.CO(n_76), .S(n_77), .A(in_21[0]), .B(n_10), .CI(in_37[0]));
  INVX1 g9460(.Y(n_75), .A(n_51));
  INVX1 g9461(.Y(n_74), .A(n_50));
  ADDFX1 g9462(.CO(n_72), .S(n_73), .A(in_49[0]), .B(n_16), .CI(n_6));
  ADDFX1 g9463(.CO(n_70), .S(n_71), .A(in_9[0]), .B(in_11[0]), .CI(in_40[0]));
  ADDFX1 g9464(.CO(n_68), .S(n_69), .A(in_27[1]), .B(in_74[1]), .CI(in_67[0]));
  ADDFX1 g9465(.CO(n_66), .S(n_67), .A(in_8[0]), .B(in_13[0]), .CI(n_22));
  ADDFX1 g9466(.CO(n_64), .S(n_65), .A(in_23[0]), .B(in_49[0]), .CI(in_63[0]));
  ADDFX1 g9467(.CO(n_62), .S(n_63), .A(in_57[0]), .B(in_68), .CI(n_23));
  ADDFX1 g9468(.CO(n_60), .S(n_61), .A(in_20[0]), .B(in_43), .CI(n_12));
  ADDFX1 g9469(.CO(n_58), .S(n_59), .A(in_12[0]), .B(in_29[0]), .CI(in_81));
  ADDFX1 g9470(.CO(n_56), .S(n_57), .A(in_34[0]), .B(n_5), .CI(in_48[0]));
  ADDFX1 g9471(.CO(n_54), .S(n_55), .A(in_6[0]), .B(in_25[0]), .CI(in_28[0]));
  ADDFX1 g9472(.CO(n_52), .S(n_53), .A(in_28[1]), .B(n_9), .CI(n_3));
  ADDFX1 g9473(.CO(n_50), .S(n_51), .A(in_47[2]), .B(in_48[0]), .CI(in_54[0]));
  ADDFX1 g9474(.CO(n_48), .S(n_49), .A(in_17[1]), .B(in_26[1]), .CI(n_1));
  ADDFX1 g9475(.CO(n_46), .S(n_47), .A(in_37[0]), .B(in_54[0]), .CI(in_67[0]));
  ADDFX1 g9476(.CO(n_44), .S(n_45), .A(n_18), .B(in_66[1]), .CI(in_55[0]));
  ADDFX1 g9477(.CO(n_42), .S(n_43), .A(in_42), .B(in_72[0]), .CI(in_78));
  ADDFX1 g9478(.CO(n_40), .S(n_41), .A(n_2), .B(in_77[1]), .CI(in_82[0]));
  ADDFX1 g9479(.CO(n_38), .S(n_39), .A(in_16[0]), .B(n_20), .CI(in_50));
  ADDFX1 g9480(.CO(n_36), .S(n_37), .A(in_31[1]), .B(in_15[1]), .CI(in_34[0]));
  ADDFX1 g9481(.CO(n_34), .S(n_35), .A(n_17), .B(in_75[1]), .CI(in_19[1]));
  ADDFX1 g9482(.CO(n_32), .S(n_33), .A(in_33[0]), .B(in_58[0]), .CI(n_24));
  OAI2BB1X1 g9483(.Y(n_31), .A0N(in_3[6]), .A1N(in_2[6]), .B0(n_27));
  OAI2BB1X1 g9484(.Y(n_30), .A0N(in_18[0]), .A1N(in_71), .B0(n_26));
  XNOR2X1 g9485(.Y(n_29), .A(in_30[1]), .B(in_53[1]));
  XNOR2X1 g9486(.Y(n_28), .A(in_29[0]), .B(in_40[0]));
  OR2X1 g9487(.Y(n_27), .A(in_3[6]), .B(in_2[6]));
  OR2X1 g9488(.Y(n_26), .A(in_18[0]), .B(in_71));
  NOR2BX1 g9489(.Y(n_25), .AN(in_30[1]), .B(in_53[1]));
  INVX1 g9491(.Y(n_24), .A(in_62[0]));
  INVX1 g9492(.Y(n_23), .A(in_69[0]));
  INVX1 g9493(.Y(n_22), .A(in_51[0]));
  INVX1 g9494(.Y(n_21), .A(in_64[0]));
  INVX1 g9495(.Y(n_20), .A(in_45[0]));
  INVX1 g9496(.Y(n_19), .A(in_11[2]));
  INVX1 g9497(.Y(n_18), .A(in_59[1]));
  INVX1 g9498(.Y(n_17), .A(in_44[1]));
  INVX1 g9499(.Y(n_16), .A(in_58[0]));
  INVX1 g9500(.Y(n_15), .A(in_56[0]));
  INVX1 g9501(.Y(n_14), .A(in_37[0]));
  INVX1 g9502(.Y(n_13), .A(in_55[0]));
  INVX1 g9503(.Y(n_12), .A(in_70[0]));
  INVX1 g9504(.Y(n_11), .A(in_84[1]));
  INVX1 g9505(.Y(n_10), .A(in_38[1]));
  INVX1 g9506(.Y(n_9), .A(in_4[1]));
  INVX1 g9507(.Y(n_8), .A(in_1[0]));
  INVX1 g9508(.Y(n_7), .A(in_14[1]));
  INVX1 g9509(.Y(n_6), .A(in_13[2]));
  INVX1 g9510(.Y(n_5), .A(in_36[0]));
  INVX1 g9511(.Y(n_4), .A(in_22[1]));
  INVX1 g9512(.Y(n_3), .A(in_25[1]));
  INVX1 g9513(.Y(n_2), .A(in_12[1]));
  INVX1 g9514(.Y(n_1), .A(in_6[1]));
  NOR2BX1 g2(.Y(n_0), .AN(in_40[0]), .B(in_29[0]));
endmodule

module csa_tree_dot_product_and_ReLU_0__product_terms_gen_255__final_adder_adder_inst_add_47_23_group_359257
    (in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, 
    in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22
    , in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, 
    in_33, in_34, in_35, in_36, in_37, in_38, in_39, in_40, in_41, in_42, in_43
    , in_44, in_45, in_46, in_47, in_48, in_49, in_50, in_51, in_52, in_53, 
    in_54, in_55, in_56, in_57, in_58, in_59, in_60, in_61, in_62, in_63, in_64
    , in_65, in_66, in_67, in_68, in_69, in_70, in_71, in_72, in_73, in_74, 
    in_75, in_76, in_77, in_78, in_79, in_80, in_81, in_82, out_0);
input  in_46, in_47, in_52, in_80;
input   [9:0] in_0;
input   [9:0] in_1;
input   [6:0] in_2;
input   [6:0] in_3;
input   [6:0] in_4;
input   [6:0] in_5;
input   [6:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [5:0] in_20;
input   [5:0] in_21;
input   [5:0] in_22;
input   [5:0] in_23;
input   [5:0] in_24;
input   [5:0] in_25;
input   [5:0] in_26;
input   [5:0] in_27;
input   [5:0] in_28;
input   [5:0] in_29;
input   [5:0] in_30;
input   [5:0] in_31;
input   [4:0] in_32;
input   [4:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [2:0] in_37;
input   [4:0] in_38;
input   [1:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [4:0] in_42;
input   [4:0] in_43;
input   [4:0] in_44;
input   [2:0] in_45;
input   [2:0] in_48;
input   [4:0] in_49;
input   [4:0] in_50;
input   [4:0] in_51;
input   [1:0] in_53;
input   [4:0] in_54;
input   [4:0] in_55;
input   [1:0] in_56;
input   [4:0] in_57;
input   [4:0] in_58;
input   [4:0] in_59;
input   [4:0] in_60;
input   [2:0] in_61;
input   [1:0] in_62;
input   [4:0] in_63;
input   [1:0] in_64;
input   [4:0] in_65;
input   [4:0] in_66;
input   [4:0] in_67;
input   [1:0] in_68;
input   [4:0] in_69;
input   [4:0] in_70;
input   [2:0] in_71;
input   [4:0] in_72;
input   [4:0] in_73;
input   [1:0] in_74;
input   [4:0] in_75;
input   [4:0] in_76;
input   [1:0] in_77;
input   [4:0] in_78;
input   [1:0] in_79;
input   [1:0] in_81;
input   [4:0] in_82;
output  [9:0] out_0;
wire  n_265, n_263, n_261, n_259, n_257, n_256, n_255, n_254, n_253, n_251, 
    n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, 
    n_240, n_239, n_238, n_237, n_235, n_234, n_233, n_232, n_231, n_230, 
    n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, 
    n_219, n_218, n_217, n_216, n_215, n_213, n_212, n_211, n_210, n_209, 
    n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, 
    n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, 
    n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, 
    n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, 
    n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, 
    n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, 
    n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, 
    in_80, in_52, in_47, in_46;
wire   [9:0] out_0;
wire   [1:0] in_81;
wire   [1:0] in_79;
wire   [1:0] in_77;
wire   [1:0] in_74;
wire   [1:0] in_68;
wire   [1:0] in_64;
wire   [1:0] in_62;
wire   [1:0] in_56;
wire   [1:0] in_53;
wire   [1:0] in_39;
wire   [2:0] in_71;
wire   [2:0] in_61;
wire   [2:0] in_48;
wire   [2:0] in_45;
wire   [2:0] in_37;
wire   [4:0] in_82;
wire   [4:0] in_78;
wire   [4:0] in_76;
wire   [4:0] in_75;
wire   [4:0] in_73;
wire   [4:0] in_72;
wire   [4:0] in_70;
wire   [4:0] in_69;
wire   [4:0] in_67;
wire   [4:0] in_66;
wire   [4:0] in_65;
wire   [4:0] in_63;
wire   [4:0] in_60;
wire   [4:0] in_59;
wire   [4:0] in_58;
wire   [4:0] in_57;
wire   [4:0] in_55;
wire   [4:0] in_54;
wire   [4:0] in_51;
wire   [4:0] in_50;
wire   [4:0] in_49;
wire   [4:0] in_44;
wire   [4:0] in_43;
wire   [4:0] in_42;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_33;
wire   [4:0] in_32;
wire   [5:0] in_31;
wire   [5:0] in_30;
wire   [5:0] in_29;
wire   [5:0] in_28;
wire   [5:0] in_27;
wire   [5:0] in_26;
wire   [5:0] in_25;
wire   [5:0] in_24;
wire   [5:0] in_23;
wire   [5:0] in_22;
wire   [5:0] in_21;
wire   [5:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [6:0] in_6;
wire   [6:0] in_5;
wire   [6:0] in_4;
wire   [6:0] in_3;
wire   [6:0] in_2;
wire   [9:0] in_1;
wire   [9:0] in_0;
  assign out_0[8] = 1'b0;
  INVX1 g8467(.Y(out_0[9]), .A(n_265));
  ADDFX1 g8468(.CO(n_265), .S(out_0[7]), .A(n_27), .B(n_247), .CI(n_263));
  ADDFX1 g8469(.CO(n_263), .S(out_0[6]), .A(n_248), .B(n_253), .CI(n_261));
  ADDFX1 g8470(.CO(n_261), .S(out_0[5]), .A(n_255), .B(n_254), .CI(n_259));
  ADDFX1 g8471(.CO(n_259), .S(out_0[4]), .A(n_249), .B(n_256), .CI(n_257));
  ADDFX1 g8472(.CO(n_257), .S(out_0[3]), .A(n_241), .B(n_251), .CI(n_250));
  ADDFX1 g8473(.CO(n_255), .S(n_256), .A(n_240), .B(n_243), .CI(n_246));
  ADDFX1 g8474(.CO(n_253), .S(n_254), .A(n_239), .B(n_245), .CI(n_238));
  ADDFX1 g8475(.CO(n_251), .S(out_0[2]), .A(n_235), .B(n_242), .CI(n_232));
  ADDFX1 g8476(.CO(n_249), .S(n_250), .A(n_231), .B(n_234), .CI(n_244));
  ADDFX1 g8477(.CO(n_247), .S(n_248), .A(n_34), .B(n_225), .CI(n_237));
  ADDFX1 g8478(.CO(n_245), .S(n_246), .A(n_229), .B(n_220), .CI(n_233));
  ADDFX1 g8479(.CO(n_243), .S(n_244), .A(n_227), .B(n_215), .CI(n_230));
  ADDFX1 g8480(.CO(n_241), .S(n_242), .A(n_228), .B(n_221), .CI(n_216));
  ADDFX1 g8481(.CO(n_239), .S(n_240), .A(n_223), .B(n_201), .CI(n_218));
  ADDFX1 g8482(.CO(n_237), .S(n_238), .A(in_0[5]), .B(n_219), .CI(n_226));
  ADDFX1 g8483(.CO(n_235), .S(out_0[1]), .A(n_213), .B(n_204), .CI(n_222));
  ADDFX1 g8484(.CO(n_233), .S(n_234), .A(n_224), .B(n_207), .CI(n_202));
  ADDFX1 g8485(.CO(n_231), .S(n_232), .A(n_203), .B(n_196), .CI(n_208));
  ADDFX1 g8486(.CO(n_229), .S(n_230), .A(n_209), .B(n_195), .CI(n_206));
  ADDFX1 g8487(.CO(n_227), .S(n_228), .A(n_197), .B(n_210), .CI(n_212));
  ADDFX1 g8488(.CO(n_225), .S(n_226), .A(n_191), .B(in_1[5]), .CI(n_217));
  ADDFX1 g8489(.CO(n_223), .S(n_224), .A(n_176), .B(n_200), .CI(n_211));
  ADDFX1 g8490(.CO(n_221), .S(n_222), .A(n_190), .B(n_198), .CI(n_194));
  ADDFX1 g8491(.CO(n_219), .S(n_220), .A(n_192), .B(in_1[4]), .CI(n_205));
  ADDFX1 g8492(.CO(n_217), .S(n_218), .A(n_175), .B(n_199), .CI(in_0[4]));
  ADDFX1 g8493(.CO(n_215), .S(n_216), .A(n_189), .B(n_193), .CI(n_173));
  ADDFX1 g8494(.CO(n_213), .S(out_0[0]), .A(n_170), .B(n_188), .CI(n_122));
  ADDFX1 g8495(.CO(n_211), .S(n_212), .A(n_158), .B(n_172), .CI(n_183));
  ADDFX1 g8496(.CO(n_209), .S(n_210), .A(n_179), .B(n_161), .CI(n_181));
  ADDFX1 g8497(.CO(n_207), .S(n_208), .A(n_168), .B(n_186), .CI(in_1[2]));
  ADDFX1 g8498(.CO(n_205), .S(n_206), .A(n_178), .B(n_167), .CI(in_1[3]));
  ADDFX1 g8499(.CO(n_203), .S(n_204), .A(n_180), .B(n_187), .CI(n_174));
  ADDFX1 g8500(.CO(n_201), .S(n_202), .A(n_185), .B(n_165), .CI(in_0[3]));
  ADDFX1 g8501(.CO(n_199), .S(n_200), .A(n_159), .B(n_171), .CI(n_152));
  ADDFX1 g8502(.CO(n_197), .S(n_198), .A(n_162), .B(n_169), .CI(n_182));
  ADDFX1 g8503(.CO(n_195), .S(n_196), .A(n_160), .B(n_166), .CI(in_0[2]));
  ADDFX1 g8504(.CO(n_193), .S(n_194), .A(n_184), .B(n_121), .CI(in_0[1]));
  ADDFX1 g8505(.CO(n_191), .S(n_192), .A(n_76), .B(n_151), .CI(n_177));
  ADDFX1 g8506(.CO(n_189), .S(n_190), .A(n_141), .B(n_136), .CI(n_164));
  ADDFX1 g8507(.CO(n_187), .S(n_188), .A(n_126), .B(n_154), .CI(n_142));
  ADDFX1 g8508(.CO(n_185), .S(n_186), .A(n_120), .B(n_132), .CI(n_163));
  ADDFX1 g8509(.CO(n_183), .S(n_184), .A(n_147), .B(n_60), .CI(n_138));
  ADDFX1 g8510(.CO(n_181), .S(n_182), .A(n_156), .B(n_125), .CI(n_144));
  ADDFX1 g8511(.CO(n_179), .S(n_180), .A(n_123), .B(n_146), .CI(n_153));
  ADDFX1 g8512(.CO(n_177), .S(n_178), .A(n_129), .B(n_133), .CI(n_131));
  ADDFX1 g8513(.CO(n_175), .S(n_176), .A(n_105), .B(n_119), .CI(n_157));
  ADDFX1 g8514(.CO(n_173), .S(n_174), .A(n_114), .B(n_140), .CI(in_1[1]));
  ADDFX1 g8515(.CO(n_171), .S(n_172), .A(n_155), .B(n_115), .CI(n_143));
  ADDFX1 g8516(.CO(n_169), .S(n_170), .A(n_124), .B(n_118), .CI(n_148));
  ADDFX1 g8517(.CO(n_167), .S(n_168), .A(n_130), .B(n_139), .CI(n_134));
  ADDFX1 g8518(.CO(n_165), .S(n_166), .A(n_113), .B(n_135), .CI(n_137));
  ADDFX1 g8519(.CO(n_163), .S(n_164), .A(n_101), .B(n_107), .CI(n_109));
  ADDFX1 g8520(.CO(n_161), .S(n_162), .A(n_128), .B(n_116), .CI(n_117));
  ADDFX1 g8521(.CO(n_159), .S(n_160), .A(n_108), .B(n_127), .CI(n_112));
  ADDFX1 g8522(.CO(n_157), .S(n_158), .A(n_104), .B(n_106), .CI(n_145));
  ADDFX1 g8523(.CO(n_155), .S(n_156), .A(n_99), .B(n_97), .CI(n_64));
  ADDFX1 g8524(.CO(n_153), .S(n_154), .A(n_75), .B(n_94), .CI(n_98));
  INVX1 g8525(.Y(n_152), .A(n_150));
  INVX1 g8526(.Y(n_151), .A(n_149));
  ADDFX1 g8527(.CO(n_149), .S(n_150), .A(n_85), .B(n_110), .CI(in_2[3]));
  ADDFX1 g8528(.CO(n_147), .S(n_148), .A(n_78), .B(n_92), .CI(n_65));
  ADDFX1 g8529(.CO(n_145), .S(n_146), .A(n_68), .B(n_41), .CI(n_87));
  ADDFX1 g8530(.CO(n_143), .S(n_144), .A(n_49), .B(n_43), .CI(in_4[1]));
  ADDFX1 g8531(.CO(n_141), .S(n_142), .A(n_100), .B(n_102), .CI(n_56));
  ADDFX1 g8532(.CO(n_139), .S(n_140), .A(n_84), .B(n_103), .CI(n_67));
  ADDFX1 g8533(.CO(n_137), .S(n_138), .A(n_39), .B(n_77), .CI(in_2[1]));
  ADDFX1 g8534(.CO(n_135), .S(n_136), .A(n_96), .B(n_55), .CI(n_71));
  ADDFX1 g8535(.CO(n_133), .S(n_134), .A(n_26), .B(n_83), .CI(n_2));
  ADDFX1 g8536(.CO(n_131), .S(n_132), .A(n_89), .B(n_66), .CI(in_2[2]));
  ADDFX1 g8537(.CO(n_129), .S(n_130), .A(n_37), .B(n_95), .CI(n_51));
  ADDFX1 g8538(.CO(n_127), .S(n_128), .A(n_32), .B(n_79), .CI(n_47));
  ADDFX1 g8539(.CO(n_125), .S(n_126), .A(n_88), .B(n_48), .CI(n_69));
  ADDFX1 g8540(.CO(n_123), .S(n_124), .A(n_80), .B(n_63), .CI(n_42));
  ADDFX1 g8541(.CO(n_121), .S(n_122), .A(n_61), .B(in_0[0]), .CI(in_1[0]));
  ADDFX1 g8542(.CO(n_119), .S(n_120), .A(n_33), .B(n_73), .CI(n_70));
  ADDFX1 g8543(.CO(n_117), .S(n_118), .A(n_50), .B(n_44), .CI(n_40));
  ADDFX1 g8544(.CO(n_115), .S(n_116), .A(n_74), .B(n_62), .CI(n_91));
  ADDFX1 g8545(.CO(n_113), .S(n_114), .A(n_38), .B(n_90), .CI(n_52));
  INVX1 g8546(.Y(n_112), .A(n_111));
  ADDFX1 g8547(.CO(n_110), .S(n_111), .A(in_17[2]), .B(in_24[2]), .CI(n_81));
  ADDFX1 g8548(.CO(n_108), .S(n_109), .A(n_13), .B(in_24[1]), .CI(n_93));
  ADDFX1 g8549(.CO(n_106), .S(n_107), .A(n_28), .B(n_6), .CI(in_17[1]));
  OAI21X1 g8550(.Y(n_105), .A0(n_30), .A1(n_72), .B0(n_76));
  INVX1 g8551(.Y(n_104), .A(n_86));
  INVX1 g8552(.Y(n_103), .A(n_82));
  ADDFX1 g8553(.CO(n_101), .S(n_102), .A(in_6[0]), .B(n_31), .CI(in_9[0]));
  ADDFX1 g8554(.CO(n_99), .S(n_100), .A(in_52), .B(in_59[0]), .CI(in_80));
  ADDFX1 g8555(.CO(n_97), .S(n_98), .A(in_26[0]), .B(in_74[0]), .CI(in_72[0]));
  ADDFX1 g8556(.CO(n_95), .S(n_96), .A(n_1), .B(in_27[0]), .CI(in_48[1]));
  ADDFX1 g8557(.CO(n_93), .S(n_94), .A(in_31[0]), .B(n_12), .CI(n_4));
  ADDFX1 g8558(.CO(n_91), .S(n_92), .A(in_47), .B(in_81[0]), .CI(n_14));
  ADDFX1 g8559(.CO(n_89), .S(n_90), .A(in_61[1]), .B(n_10), .CI(n_21));
  ADDFX1 g8560(.CO(n_87), .S(n_88), .A(in_3[0]), .B(in_18[0]), .CI(in_54[0]));
  ADDFX1 g8561(.CO(n_85), .S(n_86), .A(in_35[0]), .B(in_82[2]), .CI(in_72[0]));
  ADDFX1 g8562(.CO(n_83), .S(n_84), .A(in_53[1]), .B(n_0), .CI(n_24));
  ADDFX1 g8563(.CO(n_81), .S(n_82), .A(in_11[1]), .B(in_44[1]), .CI(in_75[1]));
  ADDFX1 g8564(.CO(n_79), .S(n_80), .A(n_17), .B(n_5), .CI(in_39[0]));
  ADDFX1 g8565(.CO(n_77), .S(n_78), .A(n_9), .B(in_27[0]), .CI(in_46));
  NAND2X1 g8566(.Y(n_76), .A(n_30), .B(n_72));
  INVX1 g8567(.Y(n_75), .A(n_59));
  INVX1 g8568(.Y(n_74), .A(n_58));
  INVX1 g8569(.Y(n_73), .A(n_57));
  INVX1 g8570(.Y(n_71), .A(n_54));
  INVX1 g8571(.Y(n_70), .A(n_53));
  INVX1 g8572(.Y(n_69), .A(n_46));
  INVX1 g8573(.Y(n_68), .A(n_45));
  INVX1 g8574(.Y(n_67), .A(n_36));
  INVX1 g8575(.Y(n_66), .A(n_35));
  ADDFX1 g8576(.CO(n_64), .S(n_65), .A(in_30[0]), .B(n_8), .CI(in_77[0]));
  ADDFX1 g8577(.CO(n_62), .S(n_63), .A(in_35[0]), .B(in_62[0]), .CI(n_22));
  ADDFX1 g8578(.CO(n_60), .S(n_61), .A(in_21[0]), .B(in_4[0]), .CI(in_2[0]));
  ADDFX1 g8579(.CO(n_58), .S(n_59), .A(in_14[0]), .B(in_51[0]), .CI(in_70[0]));
  ADDFX1 g8580(.CO(n_72), .S(n_57), .A(in_12[0]), .B(in_40[0]), .CI(in_54[0]));
  ADDFX1 g8581(.CO(n_55), .S(n_56), .A(in_19[0]), .B(in_25[0]), .CI(in_23[0]));
  ADDFX1 g8582(.CO(n_53), .S(n_54), .A(in_6[1]), .B(in_9[1]), .CI(in_23[1]));
  ADDFX1 g8583(.CO(n_51), .S(n_52), .A(n_16), .B(in_37[1]), .CI(in_79[1]));
  ADDFX1 g8584(.CO(n_49), .S(n_50), .A(in_12[0]), .B(n_11), .CI(n_3));
  ADDFX1 g8585(.CO(n_47), .S(n_48), .A(in_29[0]), .B(in_16[0]), .CI(in_56[0]));
  ADDFX1 g8586(.CO(n_45), .S(n_46), .A(in_43[0]), .B(in_42[0]), .CI(in_73[0]));
  ADDFX1 g8587(.CO(n_43), .S(n_44), .A(in_24[0]), .B(n_7), .CI(in_68[0]));
  ADDFX1 g8588(.CO(n_41), .S(n_42), .A(in_40[0]), .B(n_19), .CI(in_69[0]));
  ADDFX1 g8589(.CO(n_39), .S(n_40), .A(n_18), .B(n_20), .CI(in_64[0]));
  ADDFX1 g8590(.CO(n_37), .S(n_38), .A(in_45[1]), .B(n_23), .CI(n_15));
  ADDFX1 g8591(.CO(n_35), .S(n_36), .A(in_34[1]), .B(in_78[1]), .CI(in_25[1]));
  AOI21X1 g8592(.Y(n_34), .A0(in_0[6]), .A1(in_1[6]), .B0(n_27));
  OAI21X1 g8593(.Y(n_33), .A0(in_59[0]), .A1(in_69[0]), .B0(n_29));
  OAI2BB1X1 g8594(.Y(n_32), .A0N(in_71[1]), .A1N(n_25), .B0(n_26));
  XOR2XL g8595(.Y(n_31), .A(in_33[0]), .B(in_22[0]));
  INVX1 g8596(.Y(n_30), .A(n_29));
  NAND2X1 g8597(.Y(n_29), .A(in_69[0]), .B(in_59[0]));
  NOR2X1 g8598(.Y(n_28), .A(in_33[0]), .B(in_22[0]));
  NOR2X1 g8599(.Y(n_27), .A(in_0[6]), .B(in_1[6]));
  OR2X1 g8600(.Y(n_26), .A(in_71[1]), .B(n_25));
  INVX1 g8601(.Y(n_25), .A(in_5[1]));
  INVX1 g8602(.Y(n_24), .A(in_66[1]));
  INVX1 g8603(.Y(n_23), .A(in_63[1]));
  INVX1 g8604(.Y(n_22), .A(in_65[0]));
  INVX1 g8605(.Y(n_21), .A(in_76[1]));
  INVX1 g8606(.Y(n_20), .A(in_8[0]));
  INVX1 g8607(.Y(n_19), .A(in_58[0]));
  INVX1 g8608(.Y(n_18), .A(in_7[0]));
  INVX1 g8609(.Y(n_17), .A(in_32[0]));
  INVX1 g8610(.Y(n_16), .A(in_38[1]));
  INVX1 g8611(.Y(n_15), .A(in_50[1]));
  INVX1 g8612(.Y(n_14), .A(in_15[0]));
  INVX1 g8613(.Y(n_13), .A(in_21[1]));
  INVX1 g8614(.Y(n_12), .A(in_60[0]));
  INVX1 g8615(.Y(n_11), .A(in_67[0]));
  INVX1 g8616(.Y(n_10), .A(in_57[1]));
  INVX1 g8617(.Y(n_9), .A(in_13[0]));
  INVX1 g8618(.Y(n_8), .A(in_55[0]));
  INVX1 g8619(.Y(n_7), .A(in_41[0]));
  INVX1 g8620(.Y(n_6), .A(in_19[1]));
  INVX1 g8621(.Y(n_5), .A(in_10[0]));
  INVX1 g8622(.Y(n_4), .A(in_20[0]));
  INVX1 g8623(.Y(n_3), .A(in_28[0]));
  INVX1 g8624(.Y(n_2), .A(in_4[2]));
  INVX1 g8625(.Y(n_1), .A(in_36[1]));
  INVX1 g8626(.Y(n_0), .A(in_49[1]));
endmodule

module csa_tree_dot_product_and_ReLU_1__product_terms_gen_127__adder_32s_adder_inst_add_38_20_group_100063
    (in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, 
    in_12, in_13, in_14, in_15, in_16, in_17, in_18, out_0);
input  in_2, in_3;
input   [1:0] in_0;
input   [4:0] in_1;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [4:0] in_9;
input   [4:0] in_10;
input   [4:0] in_11;
input   [4:0] in_12;
input   [1:0] in_13;
input   [4:0] in_14;
input   [2:0] in_15;
input   [4:0] in_16;
input   [1:0] in_17;
input   [1:0] in_18;
output  [9:0] out_0;
wire  n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_25, n_22, n_20, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
    n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, in_3, in_2;
wire   [9:0] out_0;
wire   [2:0] in_15;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [4:0] in_16;
wire   [4:0] in_14;
wire   [4:0] in_12;
wire   [4:0] in_11;
wire   [4:0] in_10;
wire   [4:0] in_9;
wire   [4:0] in_1;
wire   [1:0] in_18;
wire   [1:0] in_17;
wire   [1:0] in_13;
wire   [1:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  assign out_0[5] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_43), .S(n_42), .A(in_3), .B(in_2), .CI(in_15[0]));
  ADDFX1 cdnfadd_000_1(.CO(n_41), .S(n_44), .A(n_3), .B(in_7[0]), .CI(n_7));
  ADDFX1 cdnfadd_000_2(.CO(n_40), .S(n_49), .A(in_13[0]), .B(in_0[0]), .CI(n_11));
  ADDFX1 cdnfadd_000_3(.CO(n_33), .S(n_45), .A(in_5[0]), .B(in_4[0]), .CI(n_42));
  ADDFX1 cdnfadd_001_0(.CO(n_34), .S(n_39), .A(n_2), .B(in_17[1]), .CI(in_18[1]));
  ADDFX1 cdnfadd_001_1(.CO(n_38), .S(n_37), .A(in_6[1]), .B(n_8), .CI(n_1));
  ADDFX1 cdnfadd_001_2(.CO(n_36), .S(n_35), .A(n_6), .B(n_5), .CI(n_12));
  ADDFX1 cdnfadd_001_3(.CO(n_32), .S(n_31), .A(n_10), .B(n_43), .CI(n_41));
  ADDFX1 cdnfadd_001_4(.CO(n_30), .S(n_50), .A(n_37), .B(n_39), .CI(n_35));
  ADDFX1 cdnfadd_001_5(.CO(n_51), .S(n_46), .A(n_40), .B(n_33), .CI(n_31));
  ADDFX1 cdnfadd_002_0(.CO(n_28), .S(n_29), .A(n_38), .B(n_36), .CI(n_14));
  ADDFX1 cdnfadd_002_1(.CO(n_48), .S(n_47), .A(n_32), .B(n_30), .CI(n_29));
  AO21XL g230(.Y(out_0[4]), .A0(n_16), .A1(n_25), .B0(out_0[9]));
  NOR2X1 g231(.Y(out_0[9]), .A(n_16), .B(n_25));
  ADDFX1 g232(.CO(n_25), .S(out_0[3]), .A(n_17), .B(n_48), .CI(n_22));
  ADDFX1 g233(.CO(n_22), .S(out_0[2]), .A(n_51), .B(n_47), .CI(n_20));
  ADDFX1 g234(.CO(n_20), .S(out_0[1]), .A(n_18), .B(n_50), .CI(n_46));
  ADDFX1 g235(.CO(n_18), .S(out_0[0]), .A(n_44), .B(n_49), .CI(n_45));
  AOI21X1 g236(.Y(n_17), .A0(n_13), .A1(n_15), .B0(n_16));
  NOR2X1 g237(.Y(n_16), .A(n_13), .B(n_15));
  INVX1 g238(.Y(n_15), .A(n_28));
  XNOR2X1 g239(.Y(n_14), .A(n_9), .B(n_34));
  NAND2BX1 g240(.Y(n_13), .AN(n_9), .B(n_34));
  OA21X1 g241(.Y(n_12), .A0(in_15[0]), .A1(n_4), .B0(n_9));
  AOI21X1 g242(.Y(n_11), .A0(in_12[0]), .A1(in_8[0]), .B0(n_10));
  NOR2X1 g243(.Y(n_10), .A(in_12[0]), .B(in_8[0]));
  NAND2X1 g244(.Y(n_9), .A(n_4), .B(in_15[0]));
  INVX1 g245(.Y(n_8), .A(in_16[1]));
  INVX1 g246(.Y(n_7), .A(in_10[0]));
  INVX1 g247(.Y(n_6), .A(in_4[1]));
  INVX1 g248(.Y(n_5), .A(in_5[1]));
  INVX1 g249(.Y(n_4), .A(in_1[1]));
  INVX1 g250(.Y(n_3), .A(in_11[0]));
  INVX1 g251(.Y(n_2), .A(in_14[1]));
  INVX1 g252(.Y(n_1), .A(in_9[1]));
endmodule

module csa_tree_dot_product_and_ReLU_1__product_terms_gen_255__adder_64s_adder_inst_add_47_23_group_109831
    (in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, 
    in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22
    , in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, 
    in_33, in_34, in_35, in_36, in_37, in_38, in_39, in_40, in_41, in_42, out_0);
input   [5:0] in_0;
input   [5:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [4:0] in_17;
input   [4:0] in_18;
input   [5:0] in_19;
input   [4:0] in_20;
input   [4:0] in_21;
input   [4:0] in_22;
input   [1:0] in_23;
input   [4:0] in_24;
input   [2:0] in_25;
input   [4:0] in_26;
input   [1:0] in_27;
input   [1:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [4:0] in_31;
input   [4:0] in_32;
input   [1:0] in_33;
input   [4:0] in_34;
input   [4:0] in_35;
input   [4:0] in_36;
input   [1:0] in_37;
input   [4:0] in_38;
input   [2:0] in_39;
input   [4:0] in_40;
input   [2:0] in_41;
input   [4:0] in_42;
output  [9:0] out_0;
wire  n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_41, n_39, n_37, n_35, n_33, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [9:0] out_0;
wire   [2:0] in_41;
wire   [2:0] in_39;
wire   [2:0] in_25;
wire   [1:0] in_37;
wire   [1:0] in_33;
wire   [1:0] in_29;
wire   [1:0] in_28;
wire   [1:0] in_27;
wire   [1:0] in_23;
wire   [4:0] in_42;
wire   [4:0] in_40;
wire   [4:0] in_38;
wire   [4:0] in_36;
wire   [4:0] in_35;
wire   [4:0] in_34;
wire   [4:0] in_32;
wire   [4:0] in_31;
wire   [4:0] in_30;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_21;
wire   [4:0] in_20;
wire   [4:0] in_18;
wire   [4:0] in_17;
wire   [5:0] in_19;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [5:0] in_1;
wire   [5:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  ADDFX1 cdnfadd_000_0(.CO(n_129), .S(n_128), .A(in_18[0]), .B(in_37[0]), .CI(
    in_41[0]));
  ADDFX1 cdnfadd_000_1(.CO(n_127), .S(n_126), .A(n_23), .B(in_25[0]), .CI(
    in_31[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_125), .S(n_124), .A(n_5), .B(n_2), .CI(in_39[0]));
  ADDFX1 cdnfadd_000_3(.CO(n_123), .S(n_122), .A(in_17[0]), .B(n_9), .CI(n_10));
  ADDFX1 cdnfadd_000_4(.CO(n_121), .S(n_120), .A(in_9[0]), .B(in_23[0]), .CI(
    n_25));
  ADDFX1 cdnfadd_000_5(.CO(n_119), .S(n_118), .A(in_29[0]), .B(n_22), .CI(n_6));
  ADDFX1 cdnfadd_000_6(.CO(n_117), .S(n_116), .A(n_19), .B(n_15), .CI(n_14));
  ADDFX1 cdnfadd_000_7(.CO(n_115), .S(n_114), .A(in_40[0]), .B(n_20), .CI(
    in_13[0]));
  ADDFX1 cdnfadd_000_8(.CO(n_113), .S(n_112), .A(in_6[0]), .B(in_33[0]), .CI(
    in_3[0]));
  ADDFX1 cdnfadd_000_9(.CO(n_111), .S(n_110), .A(in_11[0]), .B(in_5[0]), .CI(
    in_10[0]));
  ADDFX1 cdnfadd_000_10(.CO(n_109), .S(n_108), .A(in_2[0]), .B(in_14[0]), .CI(
    in_0[0]));
  ADDFX1 cdnfadd_000_11(.CO(n_91), .S(n_90), .A(in_4[0]), .B(in_19[0]), .CI(
    n_116));
  ADDFX1 cdnfadd_000_12(.CO(n_89), .S(n_88), .A(n_120), .B(n_114), .CI(n_112));
  ADDFX1 cdnfadd_000_13(.CO(n_87), .S(n_131), .A(n_126), .B(n_128), .CI(n_124));
  ADDFX1 cdnfadd_000_14(.CO(n_86), .S(n_138), .A(n_122), .B(n_118), .CI(n_110));
  ADDFX1 cdnfadd_000_15(.CO(n_67), .S(n_132), .A(n_108), .B(n_90), .CI(n_88));
  ADDFX1 cdnfadd_001_0(.CO(n_107), .S(n_106), .A(n_4), .B(in_3[1]), .CI(in_27[1]));
  ADDFX1 cdnfadd_001_1(.CO(n_105), .S(n_104), .A(n_21), .B(in_28[1]), .CI(n_1));
  ADDFX1 cdnfadd_001_2(.CO(n_103), .S(n_102), .A(n_17), .B(in_39[0]), .CI(n_24));
  ADDFX1 cdnfadd_001_3(.CO(n_101), .S(n_100), .A(n_13), .B(in_4[1]), .CI(n_8));
  ADDFX1 cdnfadd_001_4(.CO(n_99), .S(n_98), .A(n_16), .B(n_7), .CI(in_19[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_97), .S(n_96), .A(n_29), .B(n_3), .CI(in_11[1]));
  ADDFX1 cdnfadd_001_6(.CO(n_85), .S(n_84), .A(n_127), .B(n_119), .CI(n_121));
  ADDFX1 cdnfadd_001_7(.CO(n_83), .S(n_82), .A(n_129), .B(n_125), .CI(n_113));
  ADDFX1 cdnfadd_001_8(.CO(n_81), .S(n_80), .A(n_117), .B(n_123), .CI(n_115));
  ADDFX1 cdnfadd_001_9(.CO(n_79), .S(n_78), .A(n_104), .B(n_106), .CI(n_102));
  ADDFX1 cdnfadd_001_10(.CO(n_77), .S(n_76), .A(n_111), .B(n_98), .CI(n_109));
  ADDFX1 cdnfadd_001_11(.CO(n_66), .S(n_65), .A(n_100), .B(n_96), .CI(n_87));
  ADDFX1 cdnfadd_001_12(.CO(n_64), .S(n_63), .A(n_82), .B(n_80), .CI(n_91));
  ADDFX1 cdnfadd_001_13(.CO(n_62), .S(n_61), .A(n_84), .B(n_89), .CI(n_78));
  ADDFX1 cdnfadd_001_14(.CO(n_52), .S(n_139), .A(n_76), .B(n_86), .CI(n_65));
  ADDFX1 cdnfadd_001_15(.CO(n_51), .S(n_133), .A(n_63), .B(n_67), .CI(n_61));
  ADDFX1 cdnfadd_002_0(.CO(n_95), .S(n_94), .A(in_7[2]), .B(n_12), .CI(n_11));
  ADDFX1 cdnfadd_002_1(.CO(n_93), .S(n_92), .A(n_26), .B(n_18), .CI(in_3[2]));
  ADDFX1 cdnfadd_002_2(.CO(n_75), .S(n_74), .A(in_31[0]), .B(n_28), .CI(n_107));
  ADDFX1 cdnfadd_002_3(.CO(n_73), .S(n_72), .A(n_105), .B(n_103), .CI(n_101));
  ADDFX1 cdnfadd_002_4(.CO(n_71), .S(n_70), .A(n_94), .B(n_99), .CI(n_92));
  ADDFX1 cdnfadd_002_5(.CO(n_60), .S(n_59), .A(n_97), .B(n_83), .CI(n_81));
  ADDFX1 cdnfadd_002_6(.CO(n_58), .S(n_57), .A(n_74), .B(n_85), .CI(n_72));
  ADDFX1 cdnfadd_002_7(.CO(n_56), .S(n_55), .A(n_79), .B(n_77), .CI(n_70));
  ADDFX1 cdnfadd_002_8(.CO(n_44), .S(n_50), .A(n_66), .B(n_57), .CI(n_59));
  ADDFX1 cdnfadd_002_9(.CO(n_49), .S(n_140), .A(n_64), .B(n_62), .CI(n_55));
  ADDFX1 cdnfadd_002_10(.CO(n_141), .S(n_134), .A(n_52), .B(n_51), .CI(n_50));
  ADDFX1 cdnfadd_003_0(.CO(n_69), .S(n_68), .A(n_95), .B(n_30), .CI(n_93));
  ADDFX1 cdnfadd_003_1(.CO(n_54), .S(n_53), .A(n_75), .B(n_73), .CI(n_68));
  ADDFX1 cdnfadd_003_2(.CO(n_48), .S(n_47), .A(n_71), .B(n_60), .CI(n_58));
  ADDFX1 cdnfadd_003_3(.CO(n_46), .S(n_45), .A(n_53), .B(n_56), .CI(n_44));
  ADDFX1 cdnfadd_003_4(.CO(n_142), .S(n_135), .A(n_47), .B(n_49), .CI(n_45));
  ADDFX1 cdnfadd_004_0(.CO(n_143), .S(n_130), .A(n_27), .B(n_69), .CI(n_54));
  ADDFX1 cdnfadd_004_1(.CO(n_137), .S(n_136), .A(n_48), .B(n_130), .CI(n_46));
  INVX1 g247(.Y(out_0[9]), .A(n_41));
  ADDFX1 g248(.CO(n_41), .S(out_0[5]), .A(n_143), .B(n_137), .CI(n_39));
  ADDFX1 g249(.CO(n_39), .S(out_0[4]), .A(n_142), .B(n_136), .CI(n_37));
  ADDFX1 g250(.CO(n_37), .S(out_0[3]), .A(n_141), .B(n_35), .CI(n_135));
  ADDFX1 g251(.CO(n_35), .S(out_0[2]), .A(n_140), .B(n_33), .CI(n_134));
  ADDFX1 g252(.CO(n_33), .S(out_0[1]), .A(n_31), .B(n_139), .CI(n_133));
  ADDFX1 g253(.CO(n_31), .S(out_0[0]), .A(n_131), .B(n_138), .CI(n_132));
  AOI21X1 g254(.Y(n_30), .A0(in_31[0]), .A1(in_3[3]), .B0(n_27));
  AOI2BB1X1 g255(.Y(n_29), .A0N(in_41[0]), .A1N(in_25[0]), .B0(n_28));
  AND2XL g256(.Y(n_28), .A(in_41[0]), .B(in_25[0]));
  NOR2X1 g257(.Y(n_27), .A(in_31[0]), .B(in_3[3]));
  INVX1 g258(.Y(n_26), .A(in_11[2]));
  INVX1 g259(.Y(n_25), .A(in_34[0]));
  INVX1 g260(.Y(n_24), .A(in_12[1]));
  INVX1 g261(.Y(n_23), .A(in_1[0]));
  INVX1 g262(.Y(n_22), .A(in_38[0]));
  INVX1 g263(.Y(n_21), .A(in_32[1]));
  INVX1 g264(.Y(n_20), .A(in_20[0]));
  INVX1 g265(.Y(n_19), .A(in_42[0]));
  INVX1 g266(.Y(n_18), .A(in_4[2]));
  INVX1 g267(.Y(n_17), .A(in_26[1]));
  INVX1 g268(.Y(n_16), .A(in_0[1]));
  INVX1 g269(.Y(n_15), .A(in_8[0]));
  INVX1 g270(.Y(n_14), .A(in_16[0]));
  INVX1 g271(.Y(n_13), .A(in_14[1]));
  INVX1 g272(.Y(n_12), .A(in_40[0]));
  INVX1 g273(.Y(n_11), .A(in_19[2]));
  INVX1 g274(.Y(n_10), .A(in_36[0]));
  INVX1 g275(.Y(n_9), .A(in_24[0]));
  INVX1 g276(.Y(n_8), .A(in_2[1]));
  INVX1 g277(.Y(n_7), .A(in_5[1]));
  INVX1 g278(.Y(n_6), .A(in_15[0]));
  INVX1 g279(.Y(n_5), .A(in_22[0]));
  INVX1 g280(.Y(n_4), .A(in_21[1]));
  INVX1 g281(.Y(n_3), .A(in_10[1]));
  INVX1 g282(.Y(n_2), .A(in_35[0]));
  INVX1 g283(.Y(n_1), .A(in_30[1]));
endmodule

module csa_tree_dot_product_and_ReLU_2__product_terms_gen_127__adder_64s_adder_inst_add_47_23_group_100071
    (in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, 
    in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22
    , in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, 
    in_33, in_34, in_35, in_36, in_37, in_38, out_0);
input  in_15, in_16, in_20, in_21, in_33, in_34, in_38;
input   [7:0] in_0;
input   [5:0] in_1;
input   [5:0] in_2;
input   [5:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [4:0] in_9;
input   [4:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [4:0] in_14;
input   [2:0] in_17;
input   [4:0] in_18;
input   [2:0] in_19;
input   [2:0] in_22;
input   [4:0] in_23;
input   [2:0] in_24;
input   [4:0] in_25;
input   [1:0] in_26;
input   [2:0] in_27;
input   [4:0] in_28;
input   [2:0] in_29;
input   [4:0] in_30;
input   [1:0] in_31;
input   [4:0] in_32;
input   [4:0] in_35;
input   [2:0] in_36;
input   [1:0] in_37;
output  [9:0] out_0;
wire  n_113, n_111, n_109, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_99, 
    n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_0, in_38, 
    in_34, in_33, in_21, in_20, in_16, in_15;
wire   [9:0] out_0;
wire   [1:0] in_37;
wire   [1:0] in_31;
wire   [1:0] in_26;
wire   [2:0] in_36;
wire   [2:0] in_29;
wire   [2:0] in_27;
wire   [2:0] in_24;
wire   [2:0] in_22;
wire   [2:0] in_19;
wire   [2:0] in_17;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_25;
wire   [4:0] in_23;
wire   [4:0] in_18;
wire   [4:0] in_14;
wire   [4:0] in_10;
wire   [4:0] in_9;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [5:0] in_3;
wire   [5:0] in_2;
wire   [5:0] in_1;
wire   [7:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  assign out_0[6] = 1'b0;
  INVX1 g1390(.Y(out_0[9]), .A(n_113));
  ADDFX1 g1391(.CO(n_113), .S(out_0[5]), .A(n_81), .B(n_105), .CI(n_111));
  ADDFX1 g1392(.CO(n_111), .S(out_0[4]), .A(n_106), .B(n_103), .CI(n_109));
  ADDFX1 g1393(.CO(n_109), .S(out_0[3]), .A(n_101), .B(n_104), .CI(n_107));
  ADDFX1 g1394(.CO(n_107), .S(out_0[2]), .A(n_91), .B(n_102), .CI(n_99));
  ADDFX1 g1395(.CO(n_105), .S(n_106), .A(n_93), .B(n_82), .CI(n_97));
  ADDFX1 g1396(.CO(n_103), .S(n_104), .A(n_95), .B(n_94), .CI(n_98));
  ADDFX1 g1397(.CO(n_101), .S(n_102), .A(n_71), .B(n_90), .CI(n_96));
  ADDFX1 g1398(.CO(n_99), .S(out_0[1]), .A(n_83), .B(n_72), .CI(n_92));
  ADDFX1 g1399(.CO(n_97), .S(n_98), .A(n_73), .B(n_79), .CI(n_89));
  ADDFX1 g1400(.CO(n_95), .S(n_96), .A(n_87), .B(n_74), .CI(n_86));
  ADDFX1 g1401(.CO(n_93), .S(n_94), .A(n_55), .B(n_77), .CI(n_85));
  ADDFX1 g1402(.CO(n_91), .S(n_92), .A(n_69), .B(n_76), .CI(n_88));
  ADDFX1 g1403(.CO(n_89), .S(n_90), .A(n_75), .B(n_78), .CI(n_49));
  ADDFX1 g1404(.CO(n_87), .S(n_88), .A(n_61), .B(n_59), .CI(n_68));
  ADDFX1 g1405(.CO(n_85), .S(n_86), .A(n_53), .B(n_67), .CI(in_0[2]));
  ADDFX1 g1406(.CO(n_83), .S(out_0[0]), .A(n_62), .B(n_60), .CI(n_70));
  OAI2BB1X1 g1407(.Y(n_82), .A0N(n_40), .A1N(n_80), .B0(n_81));
  OR2X1 g1408(.Y(n_81), .A(n_40), .B(n_80));
  ADDFX1 g1409(.CO(n_80), .S(n_79), .A(n_63), .B(n_46), .CI(n_3));
  ADDFX1 g1410(.CO(n_77), .S(n_78), .A(n_47), .B(n_39), .CI(n_65));
  ADDFX1 g1411(.CO(n_75), .S(n_76), .A(n_48), .B(n_32), .CI(n_66));
  ADDFX1 g1412(.CO(n_73), .S(n_74), .A(n_57), .B(n_56), .CI(n_64));
  ADDFX1 g1413(.CO(n_71), .S(n_72), .A(n_54), .B(n_58), .CI(n_50));
  ADDFX1 g1414(.CO(n_69), .S(n_70), .A(n_24), .B(n_33), .CI(n_52));
  ADDFX1 g1415(.CO(n_67), .S(n_68), .A(n_34), .B(n_25), .CI(n_51));
  ADDFX1 g1416(.CO(n_65), .S(n_66), .A(n_4), .B(in_8[1]), .CI(n_45));
  ADDFX1 g1417(.CO(n_63), .S(n_64), .A(n_21), .B(n_15), .CI(n_0));
  ADDFX1 g1418(.CO(n_61), .S(n_62), .A(n_20), .B(n_31), .CI(n_29));
  ADDFX1 g1419(.CO(n_59), .S(n_60), .A(n_18), .B(n_26), .CI(n_35));
  ADDFX1 g1420(.CO(n_57), .S(n_58), .A(n_30), .B(n_44), .CI(n_42));
  ADDFX1 g1421(.CO(n_55), .S(n_56), .A(n_13), .B(n_41), .CI(n_43));
  ADDFX1 g1422(.CO(n_53), .S(n_54), .A(n_19), .B(n_28), .CI(n_17));
  ADDFX1 g1423(.CO(n_51), .S(n_52), .A(in_15), .B(in_21), .CI(n_37));
  ADDFX1 g1424(.CO(n_49), .S(n_50), .A(n_22), .B(n_16), .CI(in_0[1]));
  ADDFX1 g1425(.CO(n_47), .S(n_48), .A(in_5[1]), .B(in_6[1]), .CI(n_23));
  XNOR2X1 g1426(.Y(n_46), .A(n_12), .B(n_38));
  XNOR2X1 g1427(.Y(n_45), .A(in_2[0]), .B(n_36));
  ADDFX1 g1428(.CO(n_43), .S(n_44), .A(in_24[0]), .B(n_7), .CI(in_29[1]));
  ADDFX1 g1429(.CO(n_41), .S(n_42), .A(in_7[0]), .B(in_36[1]), .CI(n_9));
  NOR2BX1 g1430(.Y(n_40), .AN(n_12), .B(n_38));
  INVX1 g1432(.Y(n_39), .A(n_27));
  INVX1 g1433(.Y(n_37), .A(n_14));
  ADDFX1 g1434(.CO(n_34), .S(n_35), .A(in_20), .B(in_27[0]), .CI(in_34));
  ADDFX1 g1435(.CO(n_32), .S(n_33), .A(in_33), .B(in_3[0]), .CI(in_0[0]));
  ADDFX1 g1436(.CO(n_30), .S(n_31), .A(in_24[0]), .B(in_31[0]), .CI(n_6));
  ADDFX1 g1437(.CO(n_28), .S(n_29), .A(in_5[0]), .B(in_10[0]), .CI(n_10));
  ADDFX1 g1438(.CO(n_38), .S(n_27), .A(in_5[2]), .B(in_6[2]), .CI(in_8[2]));
  ADDFX1 g1439(.CO(n_25), .S(n_26), .A(in_26[0]), .B(n_2), .CI(in_38));
  ADDFX1 g1440(.CO(n_23), .S(n_24), .A(n_8), .B(in_7[0]), .CI(n_11));
  ADDFX1 g1441(.CO(n_21), .S(n_22), .A(in_17[1]), .B(in_19[1]), .CI(in_37[1]));
  ADDFX1 g1442(.CO(n_19), .S(n_20), .A(in_1[0]), .B(in_4[0]), .CI(in_16));
  ADDFX1 g1443(.CO(n_17), .S(n_18), .A(in_2[0]), .B(in_6[0]), .CI(in_8[0]));
  ADDFX1 g1444(.CO(n_15), .S(n_16), .A(in_27[0]), .B(in_22[1]), .CI(n_5));
  ADDFX1 g1445(.CO(n_36), .S(n_14), .A(in_11[0]), .B(in_12[0]), .CI(in_13[0]));
  OAI21X1 g1446(.Y(n_13), .A0(in_10[0]), .A1(in_32[2]), .B0(n_12));
  NAND2X1 g1447(.Y(n_12), .A(in_32[2]), .B(in_10[0]));
  INVX1 g1448(.Y(n_11), .A(in_14[0]));
  INVX1 g1449(.Y(n_10), .A(in_23[0]));
  INVX1 g1450(.Y(n_9), .A(in_25[1]));
  INVX1 g1451(.Y(n_8), .A(in_9[0]));
  INVX1 g1452(.Y(n_7), .A(in_18[1]));
  INVX1 g1453(.Y(n_6), .A(in_35[0]));
  INVX1 g1454(.Y(n_5), .A(in_28[1]));
  INVX1 g1455(.Y(n_4), .A(in_3[1]));
  INVX1 g1456(.Y(n_3), .A(in_0[3]));
  INVX1 g1457(.Y(n_2), .A(in_30[0]));
  NOR2BX1 g2(.Y(n_0), .AN(in_2[0]), .B(n_36));
endmodule

module csa_tree_dot_product_and_ReLU_14__product_terms_gen_127__adder_128s_adder_inst_add_47_23_group_106211
    (in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, 
    in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22
    , in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, 
    in_33, in_34, in_35, in_36, in_37, in_38, in_39, in_40, in_41, in_42, in_43
    , in_44, in_45, in_46, in_47, in_48, in_49, in_50, in_51, in_52, in_53, 
    out_0);
input  in_33, in_49;
input   [9:0] in_0;
input   [8:0] in_1;
input   [6:0] in_2;
input   [6:0] in_3;
input   [5:0] in_4;
input   [5:0] in_5;
input   [5:0] in_6;
input   [5:0] in_7;
input   [5:0] in_8;
input   [5:0] in_9;
input   [5:0] in_10;
input   [5:0] in_11;
input   [5:0] in_12;
input   [5:0] in_13;
input   [5:0] in_14;
input   [5:0] in_15;
input   [5:0] in_16;
input   [5:0] in_17;
input   [5:0] in_18;
input   [5:0] in_19;
input   [4:0] in_20;
input   [1:0] in_21;
input   [4:0] in_22;
input   [1:0] in_23;
input   [4:0] in_24;
input   [1:0] in_25;
input   [4:0] in_26;
input   [4:0] in_27;
input   [4:0] in_28;
input   [1:0] in_29;
input   [4:0] in_30;
input   [2:0] in_31;
input   [4:0] in_32;
input   [1:0] in_34;
input   [4:0] in_35;
input   [1:0] in_36;
input   [4:0] in_37;
input   [2:0] in_38;
input   [4:0] in_39;
input   [4:0] in_40;
input   [4:0] in_41;
input   [3:0] in_42;
input   [1:0] in_43;
input   [4:0] in_44;
input   [1:0] in_45;
input   [4:0] in_46;
input   [2:0] in_47;
input   [4:0] in_48;
input   [1:0] in_50;
input   [4:0] in_51;
input   [1:0] in_52;
input   [4:0] in_53;
output  [9:0] out_0;
wire  n_179, n_177, n_175, n_173, n_171, n_170, n_169, n_168, n_167, n_166, 
    n_165, n_164, n_163, n_162, n_161, n_159, n_158, n_157, n_156, n_155, 
    n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, 
    n_144, n_143, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, 
    n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, 
    n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
    n_6, n_5, n_4, n_3, n_2, n_1, in_49, in_33;
wire   [9:0] out_0;
wire   [3:0] in_42;
wire   [2:0] in_47;
wire   [2:0] in_38;
wire   [2:0] in_31;
wire   [1:0] in_52;
wire   [1:0] in_50;
wire   [1:0] in_45;
wire   [1:0] in_43;
wire   [1:0] in_36;
wire   [1:0] in_34;
wire   [1:0] in_29;
wire   [1:0] in_25;
wire   [1:0] in_23;
wire   [1:0] in_21;
wire   [4:0] in_53;
wire   [4:0] in_51;
wire   [4:0] in_48;
wire   [4:0] in_46;
wire   [4:0] in_44;
wire   [4:0] in_41;
wire   [4:0] in_40;
wire   [4:0] in_39;
wire   [4:0] in_37;
wire   [4:0] in_35;
wire   [4:0] in_32;
wire   [4:0] in_30;
wire   [4:0] in_28;
wire   [4:0] in_27;
wire   [4:0] in_26;
wire   [4:0] in_24;
wire   [4:0] in_22;
wire   [4:0] in_20;
wire   [5:0] in_19;
wire   [5:0] in_18;
wire   [5:0] in_17;
wire   [5:0] in_16;
wire   [5:0] in_15;
wire   [5:0] in_14;
wire   [5:0] in_13;
wire   [5:0] in_12;
wire   [5:0] in_11;
wire   [5:0] in_10;
wire   [5:0] in_9;
wire   [5:0] in_8;
wire   [5:0] in_7;
wire   [5:0] in_6;
wire   [5:0] in_5;
wire   [5:0] in_4;
wire   [6:0] in_3;
wire   [6:0] in_2;
wire   [8:0] in_1;
wire   [9:0] in_0;
  assign out_0[8] = 1'b0;
  assign out_0[7] = 1'b0;
  INVX1 g5670(.Y(out_0[9]), .A(n_179));
  ADDFX1 g5671(.CO(n_179), .S(out_0[6]), .A(n_133), .B(n_165), .CI(n_177));
  ADDFX1 g5672(.CO(n_177), .S(out_0[5]), .A(n_166), .B(n_169), .CI(n_175));
  ADDFX1 g5673(.CO(n_175), .S(out_0[4]), .A(n_167), .B(n_170), .CI(n_173));
  ADDFX1 g5674(.CO(n_173), .S(out_0[3]), .A(n_161), .B(n_168), .CI(n_171));
  ADDFX1 g5675(.CO(n_171), .S(out_0[2]), .A(n_156), .B(n_159), .CI(n_162));
  ADDFX1 g5676(.CO(n_169), .S(n_170), .A(n_153), .B(n_157), .CI(n_164));
  ADDFX1 g5677(.CO(n_167), .S(n_168), .A(n_155), .B(n_154), .CI(n_158));
  ADDFX1 g5678(.CO(n_165), .S(n_166), .A(n_151), .B(n_134), .CI(n_163));
  ADDFX1 g5679(.CO(n_163), .S(n_164), .A(n_122), .B(n_147), .CI(n_152));
  ADDFX1 g5680(.CO(n_161), .S(n_162), .A(n_149), .B(n_138), .CI(n_146));
  ADDFX1 g5681(.CO(n_159), .S(out_0[1]), .A(n_141), .B(n_150), .CI(n_144));
  ADDFX1 g5682(.CO(n_157), .S(n_158), .A(n_140), .B(n_145), .CI(n_148));
  ADDFX1 g5683(.CO(n_155), .S(n_156), .A(n_111), .B(n_136), .CI(n_143));
  ADDFX1 g5684(.CO(n_153), .S(n_154), .A(n_135), .B(n_129), .CI(n_137));
  ADDFX1 g5685(.CO(n_151), .S(n_152), .A(n_125), .B(n_109), .CI(n_139));
  ADDFX1 g5686(.CO(n_149), .S(n_150), .A(n_128), .B(n_123), .CI(n_112));
  ADDFX1 g5687(.CO(n_147), .S(n_148), .A(n_131), .B(n_126), .CI(n_110));
  ADDFX1 g5688(.CO(n_145), .S(n_146), .A(n_113), .B(n_132), .CI(n_130));
  ADDFX1 g5689(.CO(n_143), .S(n_144), .A(n_114), .B(n_108), .CI(n_116));
  ADDFX1 g5690(.CO(n_141), .S(out_0[0]), .A(n_92), .B(n_78), .CI(n_124));
  ADDFX1 g5691(.CO(n_139), .S(n_140), .A(n_117), .B(in_0[3]), .CI(n_119));
  ADDFX1 g5692(.CO(n_137), .S(n_138), .A(n_118), .B(n_120), .CI(n_115));
  ADDFX1 g5693(.CO(n_135), .S(n_136), .A(n_85), .B(n_127), .CI(n_107));
  ADDFX1 g5694(.CO(n_133), .S(n_134), .A(n_25), .B(n_12), .CI(n_121));
  ADDFX1 g5695(.CO(n_131), .S(n_132), .A(n_36), .B(n_88), .CI(n_99));
  ADDFX1 g5696(.CO(n_129), .S(n_130), .A(n_96), .B(n_84), .CI(in_0[2]));
  ADDFX1 g5697(.CO(n_127), .S(n_128), .A(n_102), .B(n_94), .CI(n_105));
  ADDFX1 g5698(.CO(n_125), .S(n_126), .A(n_35), .B(n_95), .CI(n_87));
  ADDFX1 g5699(.CO(n_123), .S(n_124), .A(n_82), .B(n_106), .CI(n_80));
  ADDFX1 g5700(.CO(n_121), .S(n_122), .A(n_97), .B(n_26), .CI(in_0[4]));
  ADDFX1 g5701(.CO(n_119), .S(n_120), .A(n_93), .B(n_75), .CI(in_1[2]));
  ADDFX1 g5702(.CO(n_117), .S(n_118), .A(n_89), .B(n_103), .CI(n_101));
  ADDFX1 g5703(.CO(n_115), .S(n_116), .A(n_91), .B(n_81), .CI(in_0[1]));
  ADDFX1 g5704(.CO(n_113), .S(n_114), .A(n_104), .B(n_90), .CI(n_79));
  ADDFX1 g5705(.CO(n_111), .S(n_112), .A(n_86), .B(n_100), .CI(n_77));
  ADDFX1 g5706(.CO(n_109), .S(n_110), .A(n_83), .B(n_98), .CI(in_1[3]));
  ADDFX1 g5707(.CO(n_107), .S(n_108), .A(n_49), .B(n_76), .CI(in_1[1]));
  ADDFX1 g5708(.CO(n_105), .S(n_106), .A(n_70), .B(n_46), .CI(n_32));
  ADDFX1 g5709(.CO(n_103), .S(n_104), .A(n_47), .B(n_31), .CI(n_61));
  ADDFX1 g5710(.CO(n_101), .S(n_102), .A(n_24), .B(n_67), .CI(n_73));
  ADDFX1 g5711(.CO(n_99), .S(n_100), .A(n_72), .B(n_58), .CI(n_40));
  ADDFX1 g5712(.CO(n_97), .S(n_98), .A(n_65), .B(n_23), .CI(n_59));
  ADDFX1 g5713(.CO(n_95), .S(n_96), .A(n_57), .B(n_71), .CI(n_41));
  ADDFX1 g5714(.CO(n_93), .S(n_94), .A(n_45), .B(n_37), .CI(n_69));
  ADDFX1 g5715(.CO(n_91), .S(n_92), .A(n_68), .B(n_64), .CI(n_74));
  ADDFX1 g5716(.CO(n_89), .S(n_90), .A(n_29), .B(n_51), .CI(n_63));
  ADDFX1 g5717(.CO(n_87), .S(n_88), .A(n_22), .B(n_55), .CI(n_39));
  ADDFX1 g5718(.CO(n_85), .S(n_86), .A(n_56), .B(n_42), .CI(n_28));
  ADDFX1 g5719(.CO(n_83), .S(n_84), .A(n_60), .B(n_66), .CI(n_27));
  ADDFX1 g5720(.CO(n_81), .S(n_82), .A(n_38), .B(n_48), .CI(n_52));
  ADDFX1 g5721(.CO(n_79), .S(n_80), .A(n_54), .B(n_62), .CI(n_30));
  ADDFX1 g5722(.CO(n_77), .S(n_78), .A(n_50), .B(in_1[0]), .CI(in_0[0]));
  ADDFX1 g5723(.CO(n_75), .S(n_76), .A(in_19[1]), .B(in_13[1]), .CI(n_53));
  ADDFX1 g5724(.CO(n_73), .S(n_74), .A(in_25[0]), .B(in_36[0]), .CI(n_17));
  ADDFX1 g5725(.CO(n_71), .S(n_72), .A(in_31[0]), .B(in_7[1]), .CI(in_34[0]));
  ADDFX1 g5726(.CO(n_69), .S(n_70), .A(in_18[0]), .B(in_29[0]), .CI(in_45[0]));
  ADDFX1 g5727(.CO(n_67), .S(n_68), .A(in_5[0]), .B(in_22[0]), .CI(n_11));
  ADDFX1 g5728(.CO(n_65), .S(n_66), .A(in_42[2]), .B(n_1), .CI(n_19));
  ADDFX1 g5729(.CO(n_63), .S(n_64), .A(in_15[0]), .B(n_10), .CI(in_21[0]));
  ADDFX1 g5730(.CO(n_61), .S(n_62), .A(in_33), .B(in_49), .CI(n_4));
  INVX1 g5731(.Y(n_60), .A(n_44));
  INVX1 g5732(.Y(n_59), .A(n_43));
  INVX1 g5733(.Y(n_58), .A(n_34));
  INVX1 g5734(.Y(n_57), .A(n_33));
  ADDFX1 g5735(.CO(n_55), .S(n_56), .A(in_15[0]), .B(n_5), .CI(n_9));
  ADDFX1 g5736(.CO(n_53), .S(n_54), .A(in_9[0]), .B(in_2[0]), .CI(n_8));
  ADDFX1 g5737(.CO(n_51), .S(n_52), .A(in_10[0]), .B(in_19[0]), .CI(in_52[0]));
  ADDFX1 g5738(.CO(n_49), .S(n_50), .A(in_43[0]), .B(in_8[0]), .CI(in_17[0]));
  ADDFX1 g5739(.CO(n_47), .S(n_48), .A(n_14), .B(in_47[0]), .CI(n_16));
  ADDFX1 g5740(.CO(n_45), .S(n_46), .A(in_23[0]), .B(n_13), .CI(in_31[0]));
  ADDFX1 g5741(.CO(n_43), .S(n_44), .A(in_8[2]), .B(in_48[0]), .CI(in_13[2]));
  ADDFX1 g5742(.CO(n_41), .S(n_42), .A(in_14[1]), .B(n_6), .CI(in_38[1]));
  ADDFX1 g5743(.CO(n_39), .S(n_40), .A(in_4[1]), .B(in_10[1]), .CI(in_47[0]));
  ADDFX1 g5744(.CO(n_37), .S(n_38), .A(in_13[0]), .B(n_7), .CI(in_44[0]));
  ADDFX1 g5745(.CO(n_35), .S(n_36), .A(in_44[0]), .B(n_3), .CI(in_10[2]));
  ADDFX1 g5746(.CO(n_33), .S(n_34), .A(in_11[1]), .B(in_30[1]), .CI(in_32[1]));
  ADDFX1 g5747(.CO(n_31), .S(n_32), .A(in_34[0]), .B(n_15), .CI(n_20));
  ADDFX1 g5748(.CO(n_29), .S(n_30), .A(in_7[0]), .B(n_2), .CI(in_48[0]));
  ADDFX1 g5749(.CO(n_27), .S(n_28), .A(in_50[1]), .B(in_8[1]), .CI(n_18));
  XNOR2X1 g5750(.Y(n_26), .A(n_21), .B(in_1[4]));
  NOR2BX1 g5751(.Y(n_25), .AN(n_21), .B(in_1[4]));
  OAI21X1 g5752(.Y(n_24), .A0(in_3[1]), .A1(in_5[1]), .B0(n_22));
  OAI21X1 g5753(.Y(n_23), .A0(in_44[0]), .A1(in_10[3]), .B0(n_21));
  NAND2X1 g5754(.Y(n_22), .A(in_5[1]), .B(in_3[1]));
  NAND2X1 g5755(.Y(n_21), .A(in_44[0]), .B(in_10[3]));
  INVX1 g5756(.Y(n_20), .A(in_41[0]));
  INVX1 g5757(.Y(n_19), .A(in_53[2]));
  INVX1 g5758(.Y(n_18), .A(in_17[1]));
  INVX1 g5759(.Y(n_17), .A(in_16[0]));
  INVX1 g5760(.Y(n_16), .A(in_6[0]));
  INVX1 g5761(.Y(n_15), .A(in_37[0]));
  INVX1 g5762(.Y(n_14), .A(in_12[0]));
  INVX1 g5763(.Y(n_13), .A(in_27[0]));
  INVX1 g5764(.Y(n_12), .A(in_0[5]));
  INVX1 g5765(.Y(n_11), .A(in_46[0]));
  INVX1 g5766(.Y(n_10), .A(in_51[0]));
  INVX1 g5767(.Y(n_9), .A(in_40[1]));
  INVX1 g5768(.Y(n_8), .A(in_26[0]));
  INVX1 g5769(.Y(n_7), .A(in_20[0]));
  INVX1 g5770(.Y(n_6), .A(in_35[1]));
  INVX1 g5771(.Y(n_5), .A(in_24[1]));
  INVX1 g5772(.Y(n_4), .A(in_28[0]));
  INVX1 g5773(.Y(n_3), .A(in_19[2]));
  INVX1 g5774(.Y(n_2), .A(in_39[0]));
  INVX1 g5775(.Y(n_1), .A(in_22[0]));
endmodule

module layer1(clk, rst_n, updown, in, out);
input  clk, rst_n, updown;
input   [0:127] in;
output  [179:0] out;
wire  n_3001_danc, n_2996_danc, n_2981_danc, n_2980_danc, n_2976_danc, 
    n_2975_danc, n_2950_danc, n_2929_danc, n_2928_danc, n_2927_danc, 
    n_2926_danc, n_2925_danc, n_2871_danc, n_2870_danc, n_2867_danc, 
    n_2866_danc, n_2864_danc, n_2862_danc, n_2861_danc, n_2826_danc, 
    n_2823_danc, n_2822_danc, n_2818_danc, n_2817_danc, n_2794_danc, 
    n_2793_danc, n_2788_danc, n_2787_danc, n_2780_danc, n_2779_danc, 
    n_2773_danc, n_2772_danc, n_2757_danc, n_2667_danc, n_2631_danc, 
    n_2603_danc, n_2602_danc, n_1554, n_1553, n_1552, n_1551, n_1550, n_1549, 
    n_1548, n_1547, n_1546, n_1545, n_1544, n_1543, n_1542, n_1541, n_1540, 
    n_1539, n_1538, n_1537, n_1536, n_1535, n_1534, n_1533, n_1532, n_1531, 
    n_1530, n_1529, n_1528, n_1527, n_1526, n_1525, n_1524, n_1523, n_1522, 
    n_1521, n_1520, n_1519, n_1518, n_1517, n_1516, n_1515, n_1514, n_1513, 
    n_1512, n_1511, n_1510, n_1509, n_1508, n_1507, n_1506, n_1505, n_1504, 
    n_1503, n_1502, n_1501, n_1500, n_1499, n_1498, n_1497, n_1496, n_1495, 
    n_1494, n_1493, n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486, 
    n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478, n_1477, 
    n_1476, n_1475, n_1474, n_1473, n_1472, n_1471, n_1470, n_1469, n_1468, 
    n_1467, n_1466, n_1465, n_1464, n_1463, n_1462, n_1461, n_1460, n_1459, 
    n_1458, n_1457, n_1456, n_1455, n_1454, n_1453, n_1452, n_1451, n_1450, 
    n_1449, n_1448, n_1447, n_1446, n_1445, n_1444, n_1443, n_1442, n_1441, 
    n_1440, n_1439, n_1438, n_1437, n_1436, n_1435, n_1434, n_1433, n_1432, 
    n_1431, n_1430, n_1429, n_1428, n_1427, n_1426, n_1425, n_1424, n_1423, 
    n_1422, n_1421, n_1420, n_1419, n_1418, n_1417, n_1416, n_1415, n_1414, 
    n_1413, n_1412, n_1411, n_1410, n_1409, n_1408, n_1407, n_1406, n_1405, 
    n_1404, n_1403, n_1402, n_1401, n_1400, n_1399, n_1398, n_1397, n_1396, 
    n_1395, n_1394, n_1393, n_1392, n_1391, n_1390, n_1389, n_1388, n_1387, 
    n_1386, n_1385, n_1384, n_1383, n_1382, n_1381, n_1380, n_1379, n_1378, 
    n_1246, n_1245, n_1244, n_1243, n_1242, n_1241, n_1240, n_1239, n_1238, 
    n_1237, n_1236, n_1235, n_1234, n_1233, n_1232, n_1231, n_1230, n_1229, 
    n_1228, n_1227, n_1226, n_1225, n_1224, n_1223, n_1222, n_1221, n_1220, 
    n_1219, n_1218, n_1216, n_1215, n_1214, n_1213, n_1212, n_1211, n_1210, 
    n_1209, n_1208, n_1207, n_1206, n_1205, n_1204, n_1203, n_1202, n_1201, 
    n_1200, n_1199, n_1198, n_1197, n_1196, n_1195, n_1194, n_1193, n_1192, 
    n_1191, n_1190, n_1189, n_1188, n_1187, n_1186, n_1185, n_1184, n_1183, 
    n_1182, n_1181, n_1180, n_1179, n_1178, n_1177, n_1176, n_1175, n_1174, 
    n_1173, n_1172, n_1171, n_1170, n_1169, n_1168, n_1167, n_1166, n_1165, 
    n_1164, n_1163, n_1162, n_1161, n_1160, n_1159, n_1158, n_1157, n_1156, 
    n_1155, n_1154, n_1153, n_1152, n_1151, n_1150, n_1149, n_1148, n_1147, 
    n_1146, n_1145, n_1144, n_1143, n_1142, n_1141, n_1140, n_1139, n_1138, 
    n_1137, n_1136, n_1135, n_1134, n_1133, n_1132, n_1131, n_1130, n_1129, 
    n_1128, n_1127, n_1126, n_1125, n_1124, n_1123, n_1122, n_1121, n_1120, 
    n_1119, n_1118, n_1117, n_1116, n_1115, n_1114, n_1113, n_1112, n_1111, 
    n_1110, n_1109, n_1108, n_1107, n_1106, n_1105, n_1104, n_1103, n_1102, 
    n_1101, n_1100, n_1099, n_1098, n_1097, n_1096, n_1095, n_1094, n_1093, 
    n_1092, n_1091, n_1090, n_1089, n_1088, n_1087, n_1086, n_1085, n_1084, 
    n_1083, n_1082, n_1081, n_1080, n_1079, n_1078, n_1077, n_1076, n_1075, 
    n_1074, n_1073, n_1072, n_1071, n_1070, n_1069, n_1068, n_1067, n_1066, 
    n_1065, n_1064, n_1063, n_1062, n_1061, n_1060, n_1059, n_1058, n_1057, 
    n_1056, n_1055, n_1054, n_1053, n_1052, n_1051, n_1050, n_1049, n_1048, 
    n_1047, n_1046, n_1045, n_1044, n_1043, n_1042, n_1041, n_1040, n_1039, 
    n_1038, n_1037, n_1036, n_1035, n_1034, n_1033, n_1032, n_1031, n_1030, 
    n_1029, n_1028, n_1027, n_1026, n_1025, n_1024, n_1023, n_1022, n_1021, 
    n_1020, n_1019, n_1018, n_1017, n_1016, n_1015, n_1014, n_1013, n_1012, 
    n_1011, n_1010, n_1009, n_1008, n_1007, n_1006, n_1005, n_1004, n_1003, 
    n_1002, n_1001, n_1000, n_999, n_998, n_997, n_996, n_995, n_994, n_993, 
    n_992, n_991, n_990, n_989, n_988, n_987, n_986, n_985, n_984, n_983, 
    n_982, n_981, n_980, n_979, n_978, n_977, n_976, n_975, n_974, n_973, 
    n_972, n_971, n_970, n_969, n_968, n_967, n_966, n_965, n_964, n_963, 
    n_962, n_961, n_960, n_959, n_958, n_957, n_956, n_955, n_954, n_953, 
    n_952, n_951, n_950, n_949, n_948, n_947, n_946, n_945, n_944, n_943, 
    n_942, n_941, n_940, n_939, n_938, n_937, n_936, n_935, n_934, n_933, 
    n_932, n_931, n_930, n_929, n_928, n_927, n_926, n_925, n_924, n_923, 
    n_922, n_921, n_920, n_919, n_918, n_917, n_916, n_915, n_914, n_913, 
    n_912, n_911, n_910, n_909, n_908, n_907, n_906, n_905, n_904, n_903, 
    n_902, n_901, n_900, n_899, n_898, n_897, n_896, n_895, n_894, n_893, 
    n_892, n_891, n_890, n_889, n_888, n_887, n_886, n_885, n_884, n_883, 
    n_882, n_881, n_880, n_879, n_878, n_877, n_876, n_875, n_874, n_873, 
    n_872, n_871, n_870, n_869, n_868, n_867, n_866, n_865, n_864, n_863, 
    n_862, n_861, n_860, n_859, n_858, n_857, n_856, n_855, n_854, n_853, 
    n_852, n_851, n_850, n_849, n_848, n_847, n_846, n_845, n_844, n_843, 
    n_842, n_841, n_840, n_839, n_838, n_837, n_836, n_835, n_834, n_833, 
    n_832, n_831, n_830, n_829, n_828, n_827, n_826, n_825, n_824, n_823, 
    n_822, n_821, n_820, n_819, n_818, n_817, n_816, n_815, n_814, n_813, 
    n_812, n_811, n_810, n_809, n_808, n_807, n_806, n_805, n_804, n_803, 
    n_802, n_801, n_800, n_799, n_798, n_797, n_796, n_795, n_794, n_793, 
    n_792, n_791, n_790, n_789, n_788, n_787, n_786, n_785, n_784, n_783, 
    n_782, n_781, n_780, n_779, n_778, n_777, n_776, n_775, n_774, n_773, 
    n_772, n_771, n_770, n_769, n_768, n_767, n_766, n_765, n_764, n_763, 
    n_762, n_761, n_760, n_759, n_758, n_757, n_756, n_755, n_754, n_753, 
    n_752, n_751, n_750, n_749, n_748, n_747, n_746, n_745, n_744, n_743, 
    n_742, n_741, n_740, n_739, n_738, n_737, n_736, n_735, n_734, n_733, 
    n_732, n_731, n_730, n_729, n_728, n_727, n_726, n_725, n_724, n_723, 
    n_722, n_721, n_720, n_719, n_718, n_717, n_716, n_715, n_714, n_713, 
    n_712, n_711, n_710, n_709, n_708, n_707, n_706, n_705, n_704, n_703, 
    n_702, n_701, n_700, n_699, n_698, n_697, n_696, n_695, n_694, n_693, 
    n_692, n_691, n_690, n_689, n_688, n_687, n_686, n_685, n_684, n_683, 
    n_682, n_681, n_680, n_679, n_678, n_677, n_676, n_675, n_674, n_673, 
    n_672, n_671, n_670, n_669, n_668, n_667, n_666, n_665, n_664, n_663, 
    n_662, n_661, n_660, n_659, n_658, n_657, n_656, n_655, n_654, n_653, 
    n_652, n_651, n_650, n_649, n_648, n_647, n_646, n_645, n_644, n_643, 
    n_642, n_641, n_640, n_639, n_638, n_637, n_636, n_635, n_634, n_633, 
    n_632, n_631, n_630, n_629, n_628, n_627, n_626, n_625, n_624, n_623, 
    n_622, n_621, n_620, n_619, n_618, n_617, n_616, n_615, n_614, n_613, 
    n_612, n_611, n_610, n_609, n_608, n_607, n_606, n_605, n_604, n_603, 
    n_602, n_601, n_600, n_599, n_598, n_597, n_596, n_595, n_594, n_593, 
    n_592, n_591, n_590, n_589, n_588, n_587, n_586, n_585, n_584, n_583, 
    n_582, n_581, n_580, n_579, n_578, n_577, n_576, n_575, n_574, n_573, 
    n_572, n_571, n_570, n_569, n_568, n_567, n_566, n_565, n_564, n_563, 
    n_562, n_561, n_560, n_559, n_558, n_557, n_556, n_555, n_554, n_553, 
    n_552, n_551, n_550, n_549, n_548, n_547, n_546, n_545, n_544, n_543, 
    n_542, n_541, n_540, n_539, n_538, n_537, n_536, n_535, n_534, n_533, 
    n_532, n_531, n_530, n_529, n_528, n_527, n_526, n_525, n_524, n_523, 
    n_522, n_521, n_520, n_519, n_518, n_517, n_516, n_515, n_514, n_513, 
    n_512, n_511, n_510, n_509, n_508, n_507, n_506, n_505, n_504, n_503, 
    n_502, n_501, n_500, n_499, n_498, n_497, n_496, n_495, n_494, n_493, 
    n_492, n_491, n_490, n_489, n_488, n_487, n_486, n_485, n_484, n_483, 
    n_482, n_481, n_480, n_479, n_478, n_477, n_476, n_475, n_474, n_473, 
    n_472, n_471, n_470, n_469, n_468, n_467, n_466, n_465, n_464, n_463, 
    n_462, n_461, n_460, n_459, n_458, n_457, n_456, n_455, n_454, n_453, 
    n_452, n_451, n_450, n_449, n_448, n_447, n_446, n_445, n_444, n_443, 
    n_442, n_441, n_440, n_439, n_438, n_437, n_436, n_435, n_434, n_433, 
    n_432, n_431, n_430, n_429, n_428, n_427, n_426, n_425, n_424, n_423, 
    n_422, n_421, n_420, n_419, n_418, n_417, n_416, n_415, n_414, n_413, 
    n_412, n_411, n_410, n_409, n_408, n_407, n_406, n_405, n_404, n_403, 
    n_402, n_401, n_400, n_399, n_398, n_397, n_396, n_395, n_394, n_393, 
    n_392, n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, n_383, 
    n_382, n_381, n_380, n_379, n_378, n_377, n_376, n_375, n_374, n_373, 
    n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_365, n_364, n_363, 
    n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, 
    n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, 
    n_342, n_341, n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, 
    n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, 
    n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, 
    n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, 
    n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, 
    n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, 
    n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, 
    n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, 
    n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, 
    n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, 
    n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
    n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
    n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, 
    n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, 
    n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, 
    n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
    n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, 
    n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
    n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, 
    n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
    n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
    n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, 
    n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, 
    n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1, n_0, \level_8_sums[18][8] , \level_8_sums[18][7] , 
    \level_8_sums[18][6] , \level_8_sums[18][5] , \level_8_sums[18][4] , 
    \level_8_sums[18][3] , \level_8_sums[18][2] , \level_8_sums[18][1] , 
    \level_8_sums[16][8] , \level_8_sums[16][7] , \level_8_sums[16][6] , 
    \level_8_sums[16][5] , \level_8_sums[16][4] , \level_8_sums[16][3] , 
    \level_8_sums[16][2] , \level_8_sums[16][1] , \level_8_sums[16][0] , 
    \level_8_sums[13][8] , \level_8_sums[13][7] , \level_8_sums[13][6] , 
    \level_8_sums[13][5] , \level_8_sums[12][9] , \level_8_sums[12][7] , 
    \level_8_sums[12][6] , \level_8_sums[12][5] , \level_8_sums[12][4] , 
    \level_8_sums[12][3] , \level_8_sums[12][2] , \level_8_sums[9][9] , 
    \level_8_sums[9][8] , \level_8_sums[9][7] , \level_8_sums[9][6] , 
    \level_8_sums[9][5] , \level_8_sums[9][4] , \level_8_sums[9][3] , 
    \level_8_sums[9][2] , \level_8_sums[9][1] , \level_8_sums[3][8] , 
    \level_8_sums[3][7] , \level_8_sums[3][6] , \level_8_sums[3][5] , 
    \level_8_sums[3][4] , \level_8_sums[3][3] , \level_8_sums[3][2] , 
    \level_8_sums[3][1] , \level_8_sums[3][0] , \level_4_sums[16][10][7] , 
    \level_4_sums[16][10][3] , \level_4_sums[16][10][2] , 
    \level_4_sums[16][10][1] , \level_4_sums[16][10][0] , 
    \level_4_sums[12][11][6] , \level_4_sums[12][11][3] , 
    \level_4_sums[12][11][2] , \level_4_sums[12][11][1] , 
    \level_4_sums[12][11][0] , \level_3_sums[19][22][4] , 
    \level_3_sums[19][22][3] , \level_3_sums[19][22][2] , 
    \level_3_sums[19][22][1] , \level_3_sums[19][22][0] , 
    \level_3_sums[10][22][3] , \level_3_sums[10][22][2] , 
    \level_3_sums[10][22][1] , \level_3_sums[10][22][0] , 
    \level_3_sums[2][12][3] , \level_3_sums[2][12][2] , 
    \level_3_sums[2][12][1] , \level_3_sums[2][12][0] , 
    \level_2_sums[17][29][2] , \level_2_sums[17][29][1] , 
    \level_2_sums[17][25][4] , \level_2_sums[17][25][2] , 
    \level_2_sums[17][25][1] , \level_2_sums[17][25][0] , 
    \level_1_sums[4][37][1] , \level_1_sums[1][81][0] , \final_sums[18][0] , 
    \final_sums[13][4] , \final_sums[13][3] , \final_sums[13][2] , 
    \final_sums[13][1] , \final_sums[13][0] , \final_sums[12][1] , 
    \final_sums[12][0] , \final_sums[9][0] , 
    \dot_product_and_ReLU[19].product_terms[138][0] , 
    \dot_product_and_ReLU[19].product_terms[60][2] , 
    \dot_product_and_ReLU[19].product_terms[59][1] , 
    \dot_product_and_ReLU[19].product_terms[48][1] , 
    \dot_product_and_ReLU[19].product_terms[46][2] , 
    \dot_product_and_ReLU[19].product_terms[26][2] , 
    \dot_product_and_ReLU[19].product_terms[2][0] , 
    \dot_product_and_ReLU[18].product_terms[186][0] , 
    \dot_product_and_ReLU[18].product_terms[183][1] , 
    \dot_product_and_ReLU[18].product_terms[153][0] , 
    \dot_product_and_ReLU[17].product_terms[156][2] , 
    \dot_product_and_ReLU[17].product_terms[124][0] , 
    \dot_product_and_ReLU[17].product_terms[112][2] , 
    \dot_product_and_ReLU[17].product_terms[53][1] , 
    \dot_product_and_ReLU[16].product_terms[107][0] , 
    \dot_product_and_ReLU[16].product_terms[102][2] , 
    \dot_product_and_ReLU[16].product_terms[71][0] , 
    \dot_product_and_ReLU[16].product_terms[12][0] , 
    \dot_product_and_ReLU[15].product_terms[61][1] , 
    \dot_product_and_ReLU[14].product_terms[154][0] , 
    \dot_product_and_ReLU[14].product_terms[131][0] , 
    \dot_product_and_ReLU[14].product_terms[99][0] , 
    \dot_product_and_ReLU[14].product_terms[18][0] , 
    \dot_product_and_ReLU[13].product_terms[89][0] , 
    \dot_product_and_ReLU[12].product_terms[87][0] , 
    \dot_product_and_ReLU[11].product_terms[50][0] , 
    \dot_product_and_ReLU[10].product_terms[172][1] , 
    \dot_product_and_ReLU[10].product_terms[80][0] , 
    \dot_product_and_ReLU[10].product_terms[78][1] , 
    \dot_product_and_ReLU[9].product_terms[163][0] , 
    \dot_product_and_ReLU[9].product_terms[152][0] , 
    \dot_product_and_ReLU[9].product_terms[128][1] , 
    \dot_product_and_ReLU[8].product_terms[182][0] , 
    \dot_product_and_ReLU[8].product_terms[180][0] , 
    \dot_product_and_ReLU[8].product_terms[173][1] , 
    \dot_product_and_ReLU[8].product_terms[139][0] , 
    \dot_product_and_ReLU[8].product_terms[92][1] , 
    \dot_product_and_ReLU[8].product_terms[36][0] , 
    \dot_product_and_ReLU[8].product_terms[32][1] , 
    \dot_product_and_ReLU[7].product_terms[111][0] , 
    \dot_product_and_ReLU[7].product_terms[109][1] , 
    \dot_product_and_ReLU[7].product_terms[103][0] , 
    \dot_product_and_ReLU[7].product_terms[64][1] , 
    \dot_product_and_ReLU[7].product_terms[58][0] , 
    \dot_product_and_ReLU[7].product_terms[57][2] , 
    \dot_product_and_ReLU[7].product_terms[38][1] , 
    \dot_product_and_ReLU[7].product_terms[16][0] , 
    \dot_product_and_ReLU[7].product_terms[10][0] , 
    \dot_product_and_ReLU[7].product_terms[7][0] , 
    \dot_product_and_ReLU[6].product_terms[188][1] , 
    \dot_product_and_ReLU[6].product_terms[43][0] , 
    \dot_product_and_ReLU[6].product_terms[14][1] , 
    \dot_product_and_ReLU[6].product_terms[9][0] , 
    \dot_product_and_ReLU[5].product_terms[185][0] , 
    \dot_product_and_ReLU[5].product_terms[160][1] , 
    \dot_product_and_ReLU[5].product_terms[96][0] , 
    \dot_product_and_ReLU[5].product_terms[75][0] , 
    \dot_product_and_ReLU[5].product_terms[72][0] , 
    \dot_product_and_ReLU[5].product_terms[51][1] , 
    \dot_product_and_ReLU[4].product_terms[190][1] , 
    \dot_product_and_ReLU[4].product_terms[166][0] , 
    \dot_product_and_ReLU[4].product_terms[146][0] , 
    \dot_product_and_ReLU[4].product_terms[136][1] , 
    \dot_product_and_ReLU[4].product_terms[133][0] , 
    \dot_product_and_ReLU[4].product_terms[127][0] , 
    \dot_product_and_ReLU[4].product_terms[126][1] , 
    \dot_product_and_ReLU[4].product_terms[125][1] , 
    \dot_product_and_ReLU[4].product_terms[118][0] , 
    \dot_product_and_ReLU[4].product_terms[101][1] , 
    \dot_product_and_ReLU[4].product_terms[98][1] , 
    \dot_product_and_ReLU[4].product_terms[97][0] , 
    \dot_product_and_ReLU[4].product_terms[82][0] , 
    \dot_product_and_ReLU[4].product_terms[79][0] , 
    \dot_product_and_ReLU[4].product_terms[68][0] , 
    \dot_product_and_ReLU[4].product_terms[24][0] , 
    \dot_product_and_ReLU[4].product_terms[20][0] , 
    \dot_product_and_ReLU[4].product_terms[15][0] , 
    \dot_product_and_ReLU[4].product_terms[3][0] , 
    \dot_product_and_ReLU[4].product_terms[1][0] , 
    \dot_product_and_ReLU[3].product_terms[184][1] , 
    \dot_product_and_ReLU[3].product_terms[181][0] , 
    \dot_product_and_ReLU[3].product_terms[178][0] , 
    \dot_product_and_ReLU[3].product_terms[168][0] , 
    \dot_product_and_ReLU[3].product_terms[164][0] , 
    \dot_product_and_ReLU[3].product_terms[161][0] , 
    \dot_product_and_ReLU[3].product_terms[151][0] , 
    \dot_product_and_ReLU[3].product_terms[123][1] , 
    \dot_product_and_ReLU[3].product_terms[120][1] , 
    \dot_product_and_ReLU[3].product_terms[110][0] , 
    \dot_product_and_ReLU[3].product_terms[86][0] , 
    \dot_product_and_ReLU[3].product_terms[84][0] , 
    \dot_product_and_ReLU[3].product_terms[83][0] , 
    \dot_product_and_ReLU[3].product_terms[81][0] , 
    \dot_product_and_ReLU[3].product_terms[54][0] , 
    \dot_product_and_ReLU[3].product_terms[47][1] , 
    \dot_product_and_ReLU[3].product_terms[45][1] , 
    \dot_product_and_ReLU[3].product_terms[25][0] , 
    \dot_product_and_ReLU[2].product_terms[175][0] , 
    \dot_product_and_ReLU[2].product_terms[174][1] , 
    \dot_product_and_ReLU[2].product_terms[165][0] , 
    \dot_product_and_ReLU[2].product_terms[144][0] , 
    \dot_product_and_ReLU[2].product_terms[143][0] , 
    \dot_product_and_ReLU[2].product_terms[134][1] , 
    \dot_product_and_ReLU[2].product_terms[129][0] , 
    \dot_product_and_ReLU[2].product_terms[121][1] , 
    \dot_product_and_ReLU[2].product_terms[117][0] , 
    \dot_product_and_ReLU[2].product_terms[116][0] , 
    \dot_product_and_ReLU[2].product_terms[113][1] , 
    \dot_product_and_ReLU[2].product_terms[95][0] , 
    \dot_product_and_ReLU[2].product_terms[91][1] , 
    \dot_product_and_ReLU[2].product_terms[70][0] , 
    \dot_product_and_ReLU[2].product_terms[67][0] , 
    \dot_product_and_ReLU[2].product_terms[52][0] , 
    \dot_product_and_ReLU[2].product_terms[44][1] , 
    \dot_product_and_ReLU[2].product_terms[40][0] , 
    \dot_product_and_ReLU[2].product_terms[37][1] , 
    \dot_product_and_ReLU[2].product_terms[35][0] , 
    \dot_product_and_ReLU[2].product_terms[34][0] , 
    \dot_product_and_ReLU[2].product_terms[33][0] , 
    \dot_product_and_ReLU[2].product_terms[31][1] , 
    \dot_product_and_ReLU[2].product_terms[21][1] , 
    \dot_product_and_ReLU[2].product_terms[4][0] , 
    \dot_product_and_ReLU[1].product_terms[176][0] , 
    \dot_product_and_ReLU[1].product_terms[171][1] , 
    \dot_product_and_ReLU[1].product_terms[170][0] , 
    \dot_product_and_ReLU[1].product_terms[158][0] , 
    \dot_product_and_ReLU[1].product_terms[149][0] , 
    \dot_product_and_ReLU[1].product_terms[148][0] , 
    \dot_product_and_ReLU[1].product_terms[147][0] , 
    \dot_product_and_ReLU[1].product_terms[137][0] , 
    \dot_product_and_ReLU[1].product_terms[135][0] , 
    \dot_product_and_ReLU[1].product_terms[132][1] , 
    \dot_product_and_ReLU[1].product_terms[115][0] , 
    \dot_product_and_ReLU[1].product_terms[108][0] , 
    \dot_product_and_ReLU[1].product_terms[85][0] , 
    \dot_product_and_ReLU[1].product_terms[77][0] , 
    \dot_product_and_ReLU[1].product_terms[73][0] , 
    \dot_product_and_ReLU[1].product_terms[69][1] , 
    \dot_product_and_ReLU[1].product_terms[62][0] , 
    \dot_product_and_ReLU[1].product_terms[56][1] , 
    \dot_product_and_ReLU[1].product_terms[55][0] , 
    \dot_product_and_ReLU[1].product_terms[30][1] , 
    \dot_product_and_ReLU[1].product_terms[19][1] , 
    \dot_product_and_ReLU[1].product_terms[11][1] , 
    \dot_product_and_ReLU[0].product_terms[191][1] , 
    \dot_product_and_ReLU[0].product_terms[189][0] , 
    \dot_product_and_ReLU[0].product_terms[187][0] , 
    \dot_product_and_ReLU[0].product_terms[179][0] , 
    \dot_product_and_ReLU[0].product_terms[177][0] , 
    \dot_product_and_ReLU[0].product_terms[169][0] , 
    \dot_product_and_ReLU[0].product_terms[167][0] , 
    \dot_product_and_ReLU[0].product_terms[159][1] , 
    \dot_product_and_ReLU[0].product_terms[157][0] , 
    \dot_product_and_ReLU[0].product_terms[155][0] , 
    \dot_product_and_ReLU[0].product_terms[150][0] , 
    \dot_product_and_ReLU[0].product_terms[145][1] , 
    \dot_product_and_ReLU[0].product_terms[142][0] , 
    \dot_product_and_ReLU[0].product_terms[141][0] , 
    \dot_product_and_ReLU[0].product_terms[130][0] , 
    \dot_product_and_ReLU[0].product_terms[122][0] , 
    \dot_product_and_ReLU[0].product_terms[119][0] , 
    \dot_product_and_ReLU[0].product_terms[114][1] , 
    \dot_product_and_ReLU[0].product_terms[106][0] , 
    \dot_product_and_ReLU[0].product_terms[105][0] , 
    \dot_product_and_ReLU[0].product_terms[100][0] , 
    \dot_product_and_ReLU[0].product_terms[94][1] , 
    \dot_product_and_ReLU[0].product_terms[93][0] , 
    \dot_product_and_ReLU[0].product_terms[90][0] , 
    \dot_product_and_ReLU[0].product_terms[88][1] , 
    \dot_product_and_ReLU[0].product_terms[76][0] , 
    \dot_product_and_ReLU[0].product_terms[66][0] , 
    \dot_product_and_ReLU[0].product_terms[65][0] , 
    \dot_product_and_ReLU[0].product_terms[63][1] , 
    \dot_product_and_ReLU[0].product_terms[49][0] , 
    \dot_product_and_ReLU[0].product_terms[42][1] , 
    \dot_product_and_ReLU[0].product_terms[41][0] , 
    \dot_product_and_ReLU[0].product_terms[39][0] , 
    \dot_product_and_ReLU[0].product_terms[29][0] , 
    \dot_product_and_ReLU[0].product_terms[28][0] , 
    \dot_product_and_ReLU[0].product_terms[27][0] , 
    \dot_product_and_ReLU[0].product_terms[23][0] , 
    \dot_product_and_ReLU[0].product_terms[22][0] , 
    \dot_product_and_ReLU[0].product_terms[17][1] , 
    \dot_product_and_ReLU[0].product_terms[13][0] , 
    \dot_product_and_ReLU[0].product_terms[8][0] , 
    \dot_product_and_ReLU[0].product_terms[6][2] , 
    \dot_product_and_ReLU[0].product_terms[5][0] , 
    \dot_product_and_ReLU[0].product_terms[0][0] , UNCONNECTED358, 
    UNCONNECTED357, UNCONNECTED356, UNCONNECTED355, UNCONNECTED354, 
    UNCONNECTED353, UNCONNECTED352, UNCONNECTED351, UNCONNECTED350, 
    UNCONNECTED349, UNCONNECTED348, UNCONNECTED347, UNCONNECTED346, 
    UNCONNECTED345, UNCONNECTED344, UNCONNECTED343, UNCONNECTED342, 
    UNCONNECTED341, UNCONNECTED340, UNCONNECTED339, UNCONNECTED338, 
    UNCONNECTED337, UNCONNECTED336, UNCONNECTED335, UNCONNECTED334, 
    UNCONNECTED333, UNCONNECTED332, UNCONNECTED331, UNCONNECTED330, 
    UNCONNECTED329, UNCONNECTED328, UNCONNECTED327, UNCONNECTED326, 
    UNCONNECTED325, UNCONNECTED324, UNCONNECTED323, UNCONNECTED322, 
    UNCONNECTED321, UNCONNECTED320, UNCONNECTED319, UNCONNECTED318, 
    UNCONNECTED317, UNCONNECTED316, UNCONNECTED315, UNCONNECTED314, 
    UNCONNECTED313, UNCONNECTED312, UNCONNECTED311, UNCONNECTED310, 
    UNCONNECTED309, UNCONNECTED308, UNCONNECTED307, UNCONNECTED306, 
    UNCONNECTED305, UNCONNECTED304, UNCONNECTED303, UNCONNECTED302, 
    UNCONNECTED301, UNCONNECTED300, UNCONNECTED299, UNCONNECTED298, 
    UNCONNECTED297, UNCONNECTED296, UNCONNECTED295, UNCONNECTED294, 
    UNCONNECTED293, UNCONNECTED292, UNCONNECTED291, UNCONNECTED290, 
    UNCONNECTED289, UNCONNECTED288, UNCONNECTED287, UNCONNECTED286, 
    UNCONNECTED285, UNCONNECTED284, UNCONNECTED283, UNCONNECTED282, 
    UNCONNECTED281, UNCONNECTED280, UNCONNECTED279, UNCONNECTED278, 
    UNCONNECTED277, UNCONNECTED276, UNCONNECTED275, UNCONNECTED274, 
    UNCONNECTED273, UNCONNECTED272, UNCONNECTED271, UNCONNECTED270, 
    UNCONNECTED269, UNCONNECTED268, UNCONNECTED267, UNCONNECTED266, 
    UNCONNECTED265, UNCONNECTED264, UNCONNECTED263, UNCONNECTED262, 
    UNCONNECTED261, UNCONNECTED260, UNCONNECTED259, UNCONNECTED258, 
    UNCONNECTED257, UNCONNECTED256, UNCONNECTED255, UNCONNECTED254, 
    UNCONNECTED253, UNCONNECTED252, UNCONNECTED251, UNCONNECTED250, 
    UNCONNECTED249, UNCONNECTED248, UNCONNECTED247, UNCONNECTED246, 
    UNCONNECTED245, UNCONNECTED244, UNCONNECTED243, UNCONNECTED242, 
    UNCONNECTED241, UNCONNECTED240, UNCONNECTED239, UNCONNECTED238, 
    UNCONNECTED237, UNCONNECTED236, UNCONNECTED235, UNCONNECTED234, 
    UNCONNECTED233, UNCONNECTED232, UNCONNECTED231, UNCONNECTED230, 
    UNCONNECTED229, UNCONNECTED228, UNCONNECTED227, UNCONNECTED226, 
    UNCONNECTED225, UNCONNECTED224, UNCONNECTED223, UNCONNECTED222, 
    UNCONNECTED221, UNCONNECTED220, UNCONNECTED219, UNCONNECTED218, 
    UNCONNECTED217, UNCONNECTED216, UNCONNECTED215, UNCONNECTED214, 
    UNCONNECTED213, UNCONNECTED212, UNCONNECTED211, UNCONNECTED210, 
    UNCONNECTED209, UNCONNECTED208, UNCONNECTED207, UNCONNECTED206, 
    UNCONNECTED205, UNCONNECTED204, UNCONNECTED203, UNCONNECTED202, 
    UNCONNECTED201, UNCONNECTED200, UNCONNECTED199, UNCONNECTED198, 
    UNCONNECTED197, UNCONNECTED196, UNCONNECTED195, UNCONNECTED194, 
    UNCONNECTED193, UNCONNECTED192, UNCONNECTED191, UNCONNECTED190, 
    UNCONNECTED189, UNCONNECTED188, UNCONNECTED187, UNCONNECTED186, 
    UNCONNECTED185, UNCONNECTED184, UNCONNECTED183, UNCONNECTED182, 
    UNCONNECTED181, UNCONNECTED180, UNCONNECTED179, UNCONNECTED178, 
    UNCONNECTED177, UNCONNECTED176, UNCONNECTED175, UNCONNECTED174, 
    UNCONNECTED173, UNCONNECTED172, UNCONNECTED171, UNCONNECTED170, 
    UNCONNECTED169, UNCONNECTED168, UNCONNECTED167, UNCONNECTED166, 
    UNCONNECTED165, UNCONNECTED164, UNCONNECTED163, UNCONNECTED162, 
    UNCONNECTED161, UNCONNECTED160, UNCONNECTED159, UNCONNECTED158, 
    UNCONNECTED157, UNCONNECTED156, UNCONNECTED155, UNCONNECTED154, 
    UNCONNECTED153, UNCONNECTED152, UNCONNECTED151, UNCONNECTED150, 
    UNCONNECTED149, UNCONNECTED148, UNCONNECTED147, UNCONNECTED146, 
    UNCONNECTED145, UNCONNECTED144, UNCONNECTED143, UNCONNECTED142, 
    UNCONNECTED141, UNCONNECTED140, UNCONNECTED139, UNCONNECTED138, 
    UNCONNECTED137, UNCONNECTED136, UNCONNECTED135, UNCONNECTED134, 
    UNCONNECTED133, UNCONNECTED132, UNCONNECTED131, UNCONNECTED130, 
    UNCONNECTED129, UNCONNECTED128, UNCONNECTED127, UNCONNECTED126, 
    UNCONNECTED125, UNCONNECTED124, UNCONNECTED123, UNCONNECTED122, 
    UNCONNECTED121, UNCONNECTED120, UNCONNECTED119, UNCONNECTED118, 
    UNCONNECTED117, UNCONNECTED116, UNCONNECTED115, UNCONNECTED114, 
    UNCONNECTED113, UNCONNECTED112, UNCONNECTED111, UNCONNECTED110, 
    UNCONNECTED109, UNCONNECTED108, UNCONNECTED107, UNCONNECTED106, 
    UNCONNECTED105, UNCONNECTED104, UNCONNECTED103, UNCONNECTED102, 
    UNCONNECTED101, UNCONNECTED100, UNCONNECTED99, UNCONNECTED98, 
    UNCONNECTED97, UNCONNECTED96, UNCONNECTED95, UNCONNECTED94, UNCONNECTED93, 
    UNCONNECTED92, UNCONNECTED91, UNCONNECTED90, UNCONNECTED89, UNCONNECTED88, 
    UNCONNECTED87, UNCONNECTED86, UNCONNECTED85, UNCONNECTED84, UNCONNECTED83, 
    UNCONNECTED82, UNCONNECTED81, UNCONNECTED80, UNCONNECTED79, UNCONNECTED78, 
    UNCONNECTED77, UNCONNECTED76, UNCONNECTED75, UNCONNECTED74, UNCONNECTED73, 
    UNCONNECTED72, UNCONNECTED71, UNCONNECTED70, UNCONNECTED69, UNCONNECTED68, 
    UNCONNECTED67, UNCONNECTED66, UNCONNECTED65, UNCONNECTED64, UNCONNECTED63, 
    UNCONNECTED62, UNCONNECTED61, UNCONNECTED60, UNCONNECTED59, UNCONNECTED58, 
    UNCONNECTED57, UNCONNECTED56, UNCONNECTED55, UNCONNECTED54, UNCONNECTED53, 
    UNCONNECTED52, UNCONNECTED51, UNCONNECTED50, UNCONNECTED49, UNCONNECTED48, 
    UNCONNECTED47, UNCONNECTED46, UNCONNECTED45, UNCONNECTED44, UNCONNECTED43, 
    UNCONNECTED42, UNCONNECTED41, UNCONNECTED40, UNCONNECTED39, UNCONNECTED38, 
    UNCONNECTED37, UNCONNECTED36, UNCONNECTED35, UNCONNECTED34, UNCONNECTED33, 
    UNCONNECTED32, UNCONNECTED31, UNCONNECTED30, UNCONNECTED29, UNCONNECTED28, 
    UNCONNECTED27, UNCONNECTED26, UNCONNECTED25, UNCONNECTED24, UNCONNECTED23, 
    UNCONNECTED22, UNCONNECTED21, UNCONNECTED20, UNCONNECTED19, UNCONNECTED18, 
    UNCONNECTED17, UNCONNECTED16, UNCONNECTED15, UNCONNECTED14, UNCONNECTED13, 
    UNCONNECTED12, UNCONNECTED11, UNCONNECTED10, UNCONNECTED9, UNCONNECTED8, 
    UNCONNECTED7, UNCONNECTED6, UNCONNECTED5, UNCONNECTED4, UNCONNECTED3, 
    UNCONNECTED2, UNCONNECTED1, UNCONNECTED0, UNCONNECTED, updown, rst_n, clk;
wire   [8:0] \level_4_sums[14][6] ;
wire   [9:0] \level_5_sums[14][2] ;
wire   [9:0] \level_8_sums[0] ;
wire   [9:0] \level_8_sums[7] ;
wire   [9:0] \level_6_sums[0][0] ;
wire   [8:0] \level_4_sums[9][10] ;
wire   [9:0] \level_6_sums[7][3] ;
wire   [9:0] \level_6_sums[18][2] ;
wire   [9:0] \level_6_sums[7][0] ;
wire   [9:0] \level_6_sums[19][2] ;
wire   [9:0] \level_8_sums[6] ;
wire   [9:0] \final_sums[5] ;
wire   [9:0] \level_6_sums[5][2] ;
wire   [9:0] \final_sums[4] ;
wire   [9:0] \level_8_sums[10] ;
wire   [6:0] \level_2_sums[10][29] ;
wire   [7:0] \level_3_sums[10][12] ;
wire   [7:0] \level_3_sums[18][10] ;
wire   [8:0] \level_4_sums[18][4] ;
wire   [9:0] \level_7_sums[18][1] ;
wire   [9:0] \level_8_sums[19] ;
wire   [7:0] \level_3_sums[19][8] ;
wire   [7:0] \level_3_sums[19][14] ;
wire   [9:0] \level_7_sums[19][1] ;
wire   [7:0] \level_3_sums[9][8] ;
wire   [9:0] \level_7_sums[9][1] ;
wire   [9:0] \level_6_sums[5][0] ;
wire   [9:0] \level_7_sums[6][1] ;
wire   [9:0] \level_6_sums[13][2] ;
wire   [9:0] \level_6_sums[13][3] ;
wire   [9:0] \level_8_sums[8] ;
wire   [7:0] \level_3_sums[16][15] ;
wire   [9:0] \level_6_sums[16][3] ;
wire   [9:0] \level_6_sums[16][0] ;
wire   [9:0] \level_6_sums[0][3] ;
wire   [9:0] \final_sums[17] ;
wire   [9:0] \level_6_sums[17][2] ;
wire   [9:0] \level_7_sums[17][0] ;
wire   [9:0] \final_sums[14] ;
wire   [9:0] \level_6_sums[14][2] ;
wire   [9:0] \level_7_sums[14][0] ;
wire   [9:0] \level_7_sums[4][0] ;
wire   [9:0] \final_sums[2] ;
wire   [5:0] \level_1_sums[12][95] ;
wire   [6:0] \level_2_sums[2][32] ;
wire   [6:0] \level_2_sums[2][41] ;
wire   [6:0] \level_2_sums[2][45] ;
wire   [7:0] \level_3_sums[2][17] ;
wire   [7:0] \level_3_sums[2][21] ;
wire   [9:0] \level_6_sums[2][1] ;
wire   [9:0] \level_5_sums[9][4] ;
wire   [9:0] \level_7_sums[10][1] ;
wire   [9:0] \level_6_sums[10][2] ;
wire   [9:0] \level_8_sums[11] ;
wire   [8:0] \level_4_sums[11][5] ;
wire   [9:0] \level_6_sums[11][2] ;
wire   [9:0] \level_6_sums[11][3] ;
wire   [9:0] \level_8_sums[15] ;
wire   [9:0] \level_6_sums[15][3] ;
wire   [9:0] \level_6_sums[15][0] ;
wire   [9:0] \level_6_sums[4][2] ;
wire   [5:0] \level_1_sums[16][87] ;
wire   [9:0] \level_6_sums[4][1] ;
wire   [9:0] \level_7_sums[8][1] ;
wire   [9:0] \level_6_sums[8][2] ;
wire   [0:255] B;
wire   [9:0] \level_6_sums[6][2] ;
wire   [9:0] \level_6_sums[5][1] ;
wire   [9:0] \level_6_sums[17][1] ;
wire   [9:0] \level_6_sums[2][0] ;
wire   [9:0] \level_8_sums[1] ;
wire   [9:0] \level_5_sums[1][3] ;
wire   [9:0] \level_6_sums[1][2] ;
wire   [9:0] \level_6_sums[1][3] ;
wire   [5:0] \level_1_sums[12][86] ;
wire   [7:0] \level_3_sums[12][19] ;
wire   [8:0] \level_4_sums[12][8] ;
wire   [8:0] \level_4_sums[12][6] ;
wire   [9:0] \level_6_sums[12][3] ;
wire   [9:0] \level_5_sums[6][3] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[104] ;
wire   [5:0] \level_1_sums[2][73] ;
wire   [5:0] \level_1_sums[7][92] ;
wire   [5:0] \level_1_sums[3][46] ;
wire   [5:0] \level_1_sums[8][55] ;
wire   [9:0] \level_6_sums[3][3] ;
wire   [9:0] \level_6_sums[3][0] ;
wire   [179:0] out;
wire   [0:127] in;
  assign out[179] = 1'b0;
  assign out[170] = 1'b0;
  assign out[152] = 1'b0;
  assign out[143] = 1'b0;
  assign out[134] = 1'b0;
  assign out[125] = 1'b0;
  assign out[116] = 1'b0;
  assign out[107] = 1'b0;
  assign out[98] = 1'b0;
  assign out[71] = 1'b0;
  assign out[53] = 1'b0;
  assign out[44] = 1'b0;
  assign out[35] = 1'b0;
  assign out[17] = 1'b0;
  assign out[8] = 1'b0;
  WALLACE_CSA_DUMMY_OP4_group_359292 WALLACE_CSA_DUMMY_OP4_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] }), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }),
     .in_2({1'b0, 1'b0, 1'b0, \level_6_sums[3][0] [9],  \level_6_sums[3][0] [5:0] }), .in_3({1'b0, 1'b0, 
    1'b0, \level_6_sums[3][3] [9],  \level_6_sums[3][3] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[179][0] , 
    \dot_product_and_ReLU[3].product_terms[178][0] }), .in_5({1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }), .in_7({1'b0, 
    1'b0, 1'b0, \level_1_sums[8][55] [4], n_1422, \level_1_sums[8][55] [0]}),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] , 1'b0}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[102][2] , 1'b0}),
     .in_10({1'b0, 1'b0, 1'b0, n_1421, n_1420, 
    \dot_product_and_ReLU[4].product_terms[101][1] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[96][0] }), .in_12({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[95][0] }), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, \level_1_sums[3][46] [4], \level_1_sums[3][46] [0]}), .in_14({1'b0, 
    1'b0, 1'b0, 1'b0, n_1419, n_1418}), .in_15({1'b0, 1'b0, 1'b0, n_1417, 
    n_1416, \dot_product_and_ReLU[3].product_terms[84][0] }), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }),
     .in_17({1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] , 1'b0, 1'b0}), .in_18({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] }), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[65][0] , 
    \dot_product_and_ReLU[7].product_terms[64][1] }), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] }), .in_21({
    1'b0, 1'b0, 1'b0, n_1415, \level_1_sums[7][92] [0], 
    \dot_product_and_ReLU[5].product_terms[185][0] }), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[180][0] , 
    \dot_product_and_ReLU[3].product_terms[181][0] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[172][1] }),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[170][0] }), .in_25({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[168][0] }),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[1][81][0] }), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, n_1449, n_1448}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[152][0] }), .in_29({1'b0, 
    1'b0, 1'b0, 1'b0, \level_1_sums[2][73] [2], \level_1_sums[2][73] [0]}),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[142][0] }), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[135][0] , 1'b0}),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[132][1] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[130][0] , 1'b0}),
     .in_34({1'b0, \dot_product_and_ReLU[3].product_terms[123][1] , 1'b0}),
     .in_35({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[120][1] , 
    1'b0}), .in_36({1'b0, \dot_product_and_ReLU[2].product_terms[121][1] }),
     .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[119][0] }), .in_38({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] }), .in_39({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }),
     .in_40({1'b0, \dot_product_and_ReLU[2].product_terms[113][1] }), .in_41({
    \dot_product_and_ReLU[1].product_terms[108][0] , 1'b0, 1'b0}), .in_42({1'b0, 
    \dot_product_and_ReLU[7].product_terms[109][1] }), .in_43({1'b0, 
    \dot_product_and_ReLU[2].product_terms[104] [1]}), .in_44({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[105][0] }), .in_45({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[98][1] }),
     .in_46({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[99][0] }), .in_47(
    \dot_product_and_ReLU[0].product_terms[90][0] ), .in_48({
    \dot_product_and_ReLU[2].product_terms[91][1] , 1'b0}), .in_49({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 1'b0}), .in_50({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[80][0] }),
     .in_51({1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }), .in_52({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] , 1'b0}),
     .in_53({1'b0, \dot_product_and_ReLU[4].product_terms[79][0] , 1'b0}),
     .in_54({\dot_product_and_ReLU[0].product_terms[76][0] , 1'b0}), .in_55(
    \dot_product_and_ReLU[1].product_terms[77][0] ), .in_56({1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[72][0] }), .in_57({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[73][0] , 1'b0}), .in_58(
    \dot_product_and_ReLU[4].product_terms[68][0] ), .in_59({
    \dot_product_and_ReLU[1].product_terms[69][1] , 1'b0}), .in_60({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[191][1] , 1'b0}), .in_61({
    \dot_product_and_ReLU[18].product_terms[186][0] , 1'b0}), .in_62({
    \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_63({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[183][1] }), .in_64({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[174][1] , 1'b0}),
     .in_65({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[175][0] }), .in_66({1'b0, 
    \dot_product_and_ReLU[3].product_terms[164][0] }), .in_67({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[165][0] }), .in_68({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[160][1] }),
     .in_69({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[161][0] }), .in_70({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[158][0] , 1'b0}), .in_71({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0}),
     .in_72({1'b0, \dot_product_and_ReLU[14].product_terms[154][0] , 1'b0}),
     .in_73({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[155][0] }), .in_74({1'b0, 
    \dot_product_and_ReLU[0].product_terms[150][0] , 1'b0}), .in_75({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }),
     .in_76(\dot_product_and_ReLU[1].product_terms[148][0] ), .in_77({1'b0, 
    \dot_product_and_ReLU[1].product_terms[149][0] }), .in_78({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[144][0] , 1'b0}), .in_79({
    1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 1'b0}), .in_80({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 1'b0}),
     .in_81({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[141][0] , 
    1'b0}), .in_82({1'b0, \dot_product_and_ReLU[8].product_terms[139][0] }),
     .in_83({\dot_product_and_ReLU[4].product_terms[136][1] , 1'b0}), .in_84(
    \dot_product_and_ReLU[1].product_terms[137][0] ), .in_85({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }), .in_86({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}),
     .out_0({\level_8_sums[3][8] , UNCONNECTED, \level_8_sums[3][7] , 
    \level_8_sums[3][6] , \level_8_sums[3][5] , \level_8_sums[3][4] , 
    \level_8_sums[3][3] , \level_8_sums[3][2] , \level_8_sums[3][1] , 
    \level_8_sums[3][0] }));
  WALLACE_CSA_DUMMY_OP8_group_359302 WALLACE_CSA_DUMMY_OP8_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[122][0] , 
    1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[117][0] , 1'b0}), .in_3({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[102][2] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] }), .in_5({1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] , 1'b0}), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[120][1] }), .in_7({1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[121][1] }), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }), .in_9({1'b0, 
    \dot_product_and_ReLU[0].product_terms[119][0] }), .in_10({1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] }), .in_11(
    \dot_product_and_ReLU[1].product_terms[115][0] ), .in_12(
    \dot_product_and_ReLU[17].product_terms[112][2] ), .in_13({
    \dot_product_and_ReLU[2].product_terms[113][1] , 1'b0}), .in_14({
    \dot_product_and_ReLU[3].product_terms[110][0] , 1'b0}), .in_15(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .in_16({1'b0, 
    \dot_product_and_ReLU[7].product_terms[109][1] , 1'b0}), .in_17(
    \dot_product_and_ReLU[0].product_terms[106][0] ), .in_18({
    \dot_product_and_ReLU[16].product_terms[107][0] , 1'b0}), .in_19({1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[105][0] }), .in_20({
    \dot_product_and_ReLU[0].product_terms[100][0] , 1'b0}), .in_21(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .in_22({1'b0, 
    \dot_product_and_ReLU[4].product_terms[98][1] , 1'b0}), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] }), .in_24({
    \dot_product_and_ReLU[5].product_terms[96][0] , 1'b0}), .in_25(
    \dot_product_and_ReLU[4].product_terms[97][0] ), .out_0({
    \level_5_sums[6][3] [9], UNCONNECTED2, UNCONNECTED1, UNCONNECTED0,  \level_5_sums[6][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP12_group_106221 WALLACE_CSA_DUMMY_OP12_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }), .in_1({
    1'b0, 1'b0, 1'b0, \level_6_sums[12][3] [9],  \level_6_sums[12][3] [5:0] }), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[12][6] [8],  \level_4_sums[12][6] [3:0] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[12][11][6] , \level_4_sums[12][11][3] , 
    \level_4_sums[12][11][2] , \level_4_sums[12][11][1] , 
    \level_4_sums[12][11][0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[12][8] [8],  \level_4_sums[12][8] [3:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0,  \level_3_sums[12][19] [3:0] }), .in_6({1'b0, 
    1'b0, 1'b0, n_1425, n_1424, n_1423}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[120][1] , 
    \dot_product_and_ReLU[2].product_terms[121][1] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[88][1] }),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[72][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] }), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[64][1] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[60][2] }), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, n_1465, n_2773_danc}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[56][1] , 1'b0}), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] }), .in_17({
    1'b0, 1'b0, 1'b0, 1'b0, n_1413, n_2823_danc}), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, n_2975_danc, n_2976_danc}), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, n_2826_danc, n_1443}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[21][1] }), .in_22({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }), .in_23({
    1'b0, 1'b0, 1'b0, 1'b0, n_1482, n_2788_danc}), .in_24({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[13][0] , 1'b0}), .in_25({1'b0, 
    1'b0, 1'b0, n_2980_danc, n_2981_danc, 
    \dot_product_and_ReLU[1].product_terms[11][1] }), .in_26({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0}), .in_27({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[2][0] , 1'b0}),
     .in_28({1'b0, 1'b0, 1'b0, 1'b0,  \level_1_sums[12][86] [1:0] }), .in_29({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[170][0] , 1'b0}), .in_30({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[168][0] }),
     .in_31({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[160][1] }), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[148][0] }),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[144][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_35({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] , 1'b0}),
     .in_36({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[124][0] , 
    1'b0}), .in_37({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[125][1] , 1'b0}), .in_38({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[116][0] }),
     .in_39({1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }), .in_40({
    1'b0, \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}), .in_41({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] , 1'b0}),
     .in_42(\dot_product_and_ReLU[17].product_terms[112][2] ), .in_43({
    \dot_product_and_ReLU[2].product_terms[113][1] , 1'b0}), .in_44({1'b0, 
    \dot_product_and_ReLU[0].product_terms[94][1] }), .in_45({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[95][0] }), .in_46({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[92][1] , 1'b0}), .in_47({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[93][0] }), .in_48({
    1'b0, \dot_product_and_ReLU[0].product_terms[90][0] }), .in_49({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_50({1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] }), .in_51({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[12].product_terms[87][0] }), .in_52({1'b0, 
    \dot_product_and_ReLU[3].product_terms[84][0] }), .in_53({
    \dot_product_and_ReLU[1].product_terms[85][0] , 1'b0}), .in_54({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_55({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}), .in_56({
    1'b0, \dot_product_and_ReLU[10].product_terms[80][0] }), .in_57({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[81][0] , 1'b0}), .in_58({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] , 1'b0}),
     .in_59({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[79][0] }), .in_60({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[76][0] }), .in_61({1'b0, 
    \dot_product_and_ReLU[1].product_terms[77][0] }), .in_62({1'b0, 1'b0, 1'b0, 
    1'b0, \level_1_sums[4][37][1] }), .in_63({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_64({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] , 1'b0}), .in_65({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[71][0] }), .in_66(
    \dot_product_and_ReLU[4].product_terms[68][0] ), .in_67({1'b0, 
    \dot_product_and_ReLU[1].product_terms[69][1] }), .in_68({
    \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}), .in_69(
    \dot_product_and_ReLU[0].product_terms[63][1] ), .in_70({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_71({1'b0, 
    \dot_product_and_ReLU[1].product_terms[55][0] }), .in_72(
    \dot_product_and_ReLU[2].product_terms[52][0] ), .in_73({1'b0, 
    \dot_product_and_ReLU[17].product_terms[53][1] }), .in_74({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] }), .in_75({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}),
     .in_76({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[48][1] }), .in_77({1'b0, 
    \dot_product_and_ReLU[0].product_terms[49][0] }), .in_78({1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] , 1'b0}), .in_79({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[47][1] }), .in_80({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[40][0] }),
     .in_81({1'b0, \dot_product_and_ReLU[0].product_terms[41][0] }), .in_82(
    \dot_product_and_ReLU[8].product_terms[32][1] ), .in_83(
    \dot_product_and_ReLU[2].product_terms[33][0] ), .in_84({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0}), .in_85({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[31][1] , 1'b0}), .in_86({1'b0, 
    \dot_product_and_ReLU[0].product_terms[29][0] }), .in_87({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[25][0] }), .in_88({1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] }), .in_89({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[15][0] }), .in_90({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_91({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[9][0] }), .in_92(
    \dot_product_and_ReLU[2].product_terms[4][0] ), .in_93({
    \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}), .in_94({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] }), .in_95({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[1][0] , 1'b0}), .in_96({1'b0, 
    \dot_product_and_ReLU[0].product_terms[167][0] , 1'b0}), .in_97({
    \dot_product_and_ReLU[3].product_terms[164][0] , 1'b0}), .in_98({
    \dot_product_and_ReLU[2].product_terms[165][0] , 1'b0}), .in_99({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[163][0] , 1'b0}), .in_100({
    \dot_product_and_ReLU[0].product_terms[150][0] , 1'b0, 1'b0}), .in_101({
    1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }), .in_102(
    \dot_product_and_ReLU[4].product_terms[146][0] ), .in_103(
    \dot_product_and_ReLU[1].product_terms[147][0] ), .out_0({
    \level_8_sums[12][9] , UNCONNECTED3, \level_8_sums[12][7] , 
    \level_8_sums[12][6] , \level_8_sums[12][5] , \level_8_sums[12][4] , 
    \level_8_sums[12][3] , \level_8_sums[12][2] , \final_sums[12][1] , 
    \final_sums[12][0] }));
  WALLACE_CSA_DUMMY_OP17_group_106212 WALLACE_CSA_DUMMY_OP17_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }), .in_1({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[21][1] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[1][3] [9],  \level_6_sums[1][3] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 
    \level_6_sums[1][2] [9],  \level_6_sums[1][2] [5:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_5_sums[1][3] [9],  \level_5_sums[1][3] [4:0] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[39][0] }), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[65][0] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[62][0] }),
     .in_9({1'b0, 1'b0, 1'b0, n_2772_danc, n_2773_danc, 
    \dot_product_and_ReLU[7].product_terms[58][0] }), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[56][1] , 1'b0}), .in_11({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }),
     .in_12({1'b0, 1'b0, 1'b0, n_1490, n_1491, n_1489}), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, n_1485, n_2818_danc}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0}), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, n_1484, n_1483}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[26][2] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] }), .in_18({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[23][0] , 
    1'b0}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[19][1] , 1'b0}), .in_20({1'b0, 1'b0, 
    1'b0, 1'b0, n_1482, n_2788_danc}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] }), .in_22({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_23({1'b0, 
    1'b0, 1'b0, 1'b0, n_1481, n_1480}), .in_24({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_25({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[94][1] }), .in_26({1'b0, 
    \dot_product_and_ReLU[2].product_terms[95][0] , 1'b0}), .in_27({1'b0, 
    \dot_product_and_ReLU[0].product_terms[93][0] }), .in_28(
    \dot_product_and_ReLU[0].product_terms[90][0] ), .in_29(
    \dot_product_and_ReLU[2].product_terms[91][1] ), .in_30({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[88][1] }), .in_31({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 1'b0}), .in_32({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}),
     .in_33({1'b0, \dot_product_and_ReLU[1].product_terms[85][0] }), .in_34({
    1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}), .in_36({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }), .in_37({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }),
     .in_38({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[79][0] }), .in_39({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[76][0] , 1'b0}), .in_40({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[77][0] }), .in_41({1'b0, 
    1'b0, 1'b0, \level_1_sums[4][37][1] , 1'b0}), .in_42({1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_43({1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] }), .in_44({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[71][0] , 1'b0}), .in_45({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[68][0] }), .in_46({
    1'b0, \dot_product_and_ReLU[1].product_terms[69][1] , 1'b0}), .in_47({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] , 1'b0}), .in_48({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] , 1'b0}),
     .in_49({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[60][2] }), .in_50({1'b0, 
    \dot_product_and_ReLU[15].product_terms[61][1] }), .in_51({1'b0, 
    \dot_product_and_ReLU[3].product_terms[54][0] }), .in_52({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[55][0] }), .in_53({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] }), .in_54({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] }),
     .in_55({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[40][0] , 
    1'b0}), .in_56({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[41][0] }), .in_57({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[32][1] , 1'b0}), .in_58({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }), .in_59({1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] }), .in_60({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_61({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[10][0] , 1'b0}), .in_62({
    1'b0, \dot_product_and_ReLU[1].product_terms[11][1] , 1'b0}), .in_63({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0}), .in_64({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[1][0] , 1'b0}), .out_0({
    \level_8_sums[1] [8], UNCONNECTED4,  \level_8_sums[1] [7:0] }));
  WALLACE_CSA_DUMMY_OP22_group_106194 WALLACE_CSA_DUMMY_OP22_groupi(.in_0({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0}), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, n_1478, n_1477, n_1476}), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }), .in_3({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[48][1] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_5({1'b0, 1'b0, 
    n_1485, n_2818_danc, \dot_product_and_ReLU[2].product_terms[44][1] , 
    \dot_product_and_ReLU[3].product_terms[45][1] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[40][0] }), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, n_1475, n_1474}), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_10({1'b0, 
    1'b0, 1'b0, n_1473, n_1472, \dot_product_and_ReLU[1].product_terms[19][1] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1482, n_2788_danc}), .in_12({1'b0, 1'b0, 
    1'b0, n_1471, n_1470, n_1469}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[58][0] }), .in_16({
    1'b0, \dot_product_and_ReLU[19].product_terms[59][1] , 1'b0}), .in_17({1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] }), .in_18(
    \dot_product_and_ReLU[3].product_terms[54][0] ), .in_19(
    \dot_product_and_ReLU[1].product_terms[55][0] ), .in_20({1'b0, 
    \dot_product_and_ReLU[11].product_terms[50][0] }), .in_21({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] }), .in_22({1'b0, 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_23({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[43][0] }), .in_24({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[37][1] , 1'b0}), .in_25({1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[32][1] , 1'b0, 1'b0}), .in_26({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }),
     .in_27({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] }), .in_28({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[31][1] , 1'b0}), .in_29({1'b0, 
    \dot_product_and_ReLU[0].product_terms[29][0] , 1'b0}), .in_30({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[27][0] , 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[20][0] }), .in_32({
    1'b0, \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[14][1] }), .in_34({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[15][0] }),
     .in_35({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] }), .in_36({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_37({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[10][0] , 1'b0}), .in_38({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[11][1] , 1'b0}),
     .in_39({1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_40({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[9][0] , 1'b0}),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[6][2] }), .in_42({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }), .out_0({
    \level_6_sums[2][0] [9], UNCONNECTED6, UNCONNECTED5,  \level_6_sums[2][0] [6:0] }));
  WALLACE_CSA_DUMMY_OP40_group_359279 WALLACE_CSA_DUMMY_OP40_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, \level_2_sums[17][29][2] , 
    \level_2_sums[17][29][1] , \dot_product_and_ReLU[4].product_terms[118][0] }),
     .in_2({1'b0, 1'b0, 1'b0, \level_2_sums[17][25][4] , 
    \level_2_sums[17][25][2] , \level_2_sums[17][25][1] , 
    \level_2_sums[17][25][0] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[122][0] }), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[110][0] , 1'b0}), .in_5({1'b0, 
    1'b0, 1'b0, n_1438, n_1437, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_6({1'b0, 
    \dot_product_and_ReLU[4].product_terms[98][1] , 1'b0}), .in_7({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[14].product_terms[99][0] , 1'b0}), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[94][1] , 1'b0}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[84][0] , 
    \dot_product_and_ReLU[1].product_terms[85][0] }), .in_10({1'b0, 1'b0, 1'b0, 
    n_2862_danc, n_1436, \dot_product_and_ReLU[10].product_terms[80][0] }),
     .in_11({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] , 
    1'b0, 1'b0}), .in_12({1'b0, 1'b0, 1'b0, n_2866_danc, n_1215, n_2867_danc}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] , 1'b0}), .in_14({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}),
     .in_15({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] , 
    1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[124][0] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }), .in_18({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[120][1] }),
     .in_19({1'b0, \dot_product_and_ReLU[2].product_terms[121][1] }), .in_20({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }),
     .in_21({1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[112][2] , 1'b0, 
    1'b0}), .in_22({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[113][1] , 1'b0}), .in_23({1'b0, 
    \dot_product_and_ReLU[1].product_terms[108][0] , 1'b0}), .in_24({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[109][1] , 1'b0}),
     .in_25({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[92][1] , 
    1'b0}), .in_26({1'b0, \dot_product_and_ReLU[0].product_terms[93][0] }),
     .in_27({\dot_product_and_ReLU[0].product_terms[88][1] , 1'b0, 1'b0}),
     .in_28(\dot_product_and_ReLU[13].product_terms[89][0] ), .in_29({1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] }), .in_30({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[12].product_terms[87][0] }), .in_31({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[72][0] , 1'b0}), .in_32({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }),
     .in_33(\dot_product_and_ReLU[2].product_terms[70][0] ), .in_34(
    \dot_product_and_ReLU[16].product_terms[71][0] ), .in_35({1'b0, 
    \dot_product_and_ReLU[1].product_terms[69][1] }), .in_36({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[66][0] }), .in_37({1'b0, 
    \dot_product_and_ReLU[2].product_terms[67][0] , 1'b0}), .in_38({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] , 1'b0, 1'b0}), .out_0({
    \level_6_sums[17][1] [9], UNCONNECTED8, UNCONNECTED7,  \level_6_sums[17][1] [6:0] }));
  WALLACE_CSA_DUMMY_OP43_group_359277 WALLACE_CSA_DUMMY_OP43_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[95][0] }), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[118][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    n_1238, n_1237, n_1236, n_1235}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[113][1] }), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[108][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[107][0] , 1'b0}), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[96][0] }),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[92][1] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 
    \dot_product_and_ReLU[0].product_terms[88][1] }), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, n_1419, n_1418}), .in_11({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[82][0] , 1'b0}), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }), .in_13({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_15({1'b0, 1'b0, 1'b0, 
    n_1407, n_1406, \dot_product_and_ReLU[5].product_terms[72][0] }), .in_16({
    1'b0, 1'b0, 1'b0, 1'b0, n_2870_danc, n_2871_danc}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }), .in_18({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[126][1] }),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] }), .in_20({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0}), .in_21({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[120][1] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[121][1] }), .in_24({
    1'b0, \dot_product_and_ReLU[3].product_terms[110][0] }), .in_25(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .in_26({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[98][1] }), .in_27({1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[99][0] }), .in_28({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[90][0] , 1'b0}), .in_29({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] , 1'b0}), .in_30({
    \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}), .in_31(
    \dot_product_and_ReLU[1].product_terms[85][0] ), .in_32({1'b0, 1'b0, 
    \level_1_sums[4][37][1] }), .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_34({1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] }), .in_35({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[71][0] , 1'b0}), .in_36({1'b0, 
    \dot_product_and_ReLU[7].product_terms[64][1] , 1'b0}), .in_37({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[65][0] }), .out_0({
    \level_6_sums[5][1] [9], UNCONNECTED11, UNCONNECTED10, UNCONNECTED9,  \level_6_sums[5][1] [5:0] }));
  WALLACE_CSA_DUMMY_OP50_group_359285 WALLACE_CSA_DUMMY_OP50_groupi(.in_0({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[135][0] , 1'b0}), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] , 
    \dot_product_and_ReLU[0].product_terms[189][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] , 1'b0, 1'b0}), .in_3({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[175][0] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[168][0] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[164][0] , 
    \dot_product_and_ReLU[2].product_terms[165][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, n_1393, n_1392}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[157][0] , 
    \dot_product_and_ReLU[17].product_terms[156][2] }), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, n_1391, n_1390}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[148][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[143][0] , 
    \dot_product_and_ReLU[0].product_terms[142][0] }), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 1'b0}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[136][1] }), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[131][0] }),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_16({1'b0, 
    \dot_product_and_ReLU[0].product_terms[191][1] }), .in_17({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_18(
    \dot_product_and_ReLU[3].product_terms[184][1] ), .in_19({
    \dot_product_and_ReLU[5].product_terms[185][0] , 1'b0}), .in_20({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[182][0] , 1'b0}), .in_21({
    1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[183][1] , 1'b0, 1'b0}),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[178][0] }), .in_23({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[179][0] , 1'b0, 1'b0}), .in_24({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[177][0] }),
     .in_25({1'b0, \dot_product_and_ReLU[10].product_terms[172][1] }), .in_26({
    \dot_product_and_ReLU[8].product_terms[173][1] , 1'b0}), .in_27({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[170][0] }), .in_28({
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[171][1] }), .in_29({1'b0, 
    \dot_product_and_ReLU[0].product_terms[167][0] }), .in_30({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[163][0] }), .in_31({
    1'b0, \dot_product_and_ReLU[5].product_terms[160][1] }), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] }), .in_33(
    \dot_product_and_ReLU[14].product_terms[154][0] ), .in_34({
    \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[18].product_terms[153][0] , 1'b0}), .in_36({
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }), .in_37({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] }),
     .in_38({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[138][0] , 
    1'b0}), .in_39({1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 
    1'b0}), .in_40({1'b0, \dot_product_and_ReLU[1].product_terms[132][1] , 
    1'b0}), .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }), .in_43({
    1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}), .out_0({
    \level_6_sums[6][2] [9], UNCONNECTED14, UNCONNECTED13, UNCONNECTED12,  \level_6_sums[6][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP58_group_109825_6338 WALLACE_CSA_DUMMY_OP58_groupi(.in_0({
    1'b0, 1'b0, 1'b0, B[238], 1'b0}), .in_1({1'b0, B[239], 1'b0}), .in_2({1'b0, 
    1'b0, \level_6_sums[8][2] [9],  \level_6_sums[8][2] [6:0] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  B[250:251] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[215]}), .in_5({1'b0, B[247], 
    1'b0}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, n_1499, n_1498}), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, n_1515, n_1549}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, n_2667_danc, 
    n_1547}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_1514, n_1513}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, B[218]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, B[216]}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1530, n_1529}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[203]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0,  B[200:201] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, n_1540, n_1539}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, B[252]}),
     .in_17({1'b0, B[253], 1'b0, 1'b0}), .in_18({1'b0, 1'b0, 1'b0, B[243], 1'b0}),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_20({1'b0, B[241]}), .in_21({
    1'b0, B[234]}), .in_22({1'b0, 1'b0, 1'b0, B[235], 1'b0}), .in_23({1'b0, 
    1'b0, B[230]}), .in_24({1'b0, 1'b0, 1'b0, B[231], 1'b0}), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, B[228]}), .in_26({1'b0, B[229]}), .in_27(B[226]), .in_28(
    B[227]), .in_29({1'b0, 1'b0, 1'b0, 1'b0, B[222]}), .in_30({1'b0, 1'b0, 1'b0, 
    1'b0, B[223]}), .in_31({B[208], 1'b0, 1'b0}), .in_32(B[209]), .in_33({1'b0, 
    1'b0, 1'b0, 1'b0, B[206]}), .in_34({1'b0, B[207]}), .in_35({1'b0, B[204], 
    1'b0}), .in_36({1'b0, 1'b0, 1'b0, B[205], 1'b0}), .in_37({1'b0, 1'b0, 
    B[198]}), .in_38({1'b0, 1'b0, 1'b0, 1'b0, B[199]}), .in_39({1'b0, 1'b0, 
    B[195]}), .in_40(B[192]), .in_41({B[193], 1'b0, 1'b0}), .out_0({
    \level_7_sums[8][1] [9], UNCONNECTED15,  \level_7_sums[8][1] [7:0] }));
  WALLACE_CSA_DUMMY_OP58_group_109825 WALLACE_CSA_DUMMY_OP58_groupi4211(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[84][0] }), .in_2({1'b0, 
    \dot_product_and_ReLU[1].product_terms[85][0] , 1'b0}), .in_3({1'b0, 1'b0, 
    1'b0, 1'b0, \level_1_sums[8][55] [4], n_1422, \level_1_sums[8][55] [0]}),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[91][1] , 1'b0}), .in_5({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_6({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] }), .in_7({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0}),
     .in_8({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] , 
    1'b0}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_1412, n_1411}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1447, n_1446}), .in_12({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[106][0] , 1'b0}), .in_13({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[104] [1]}), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[98][1] , 1'b0}), .in_15({
    1'b0, 1'b0, 1'b0, n_1435, n_2928_danc, 
    \dot_product_and_ReLU[2].product_terms[95][0] }), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[92][1] }), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] , 1'b0}), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, n_1410, n_2871_danc}), .in_19({1'b0, 
    \dot_product_and_ReLU[2].product_terms[116][0] }), .in_20(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .in_21({1'b0, 
    \dot_product_and_ReLU[16].product_terms[102][2] }), .in_22({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[103][0] , 1'b0}), .in_23({
    1'b0, \dot_product_and_ReLU[4].product_terms[101][1] , 1'b0}), .in_24({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[96][0] }), .in_25({
    1'b0, \dot_product_and_ReLU[4].product_terms[97][0] }), .in_26({1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] }), .in_27(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .in_28({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_29({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }), .in_30({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[80][0] , 1'b0}),
     .in_31({1'b0, \dot_product_and_ReLU[3].product_terms[81][0] , 1'b0}),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[10].product_terms[78][1] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[79][0] }), .in_34({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[76][0] , 1'b0}), .in_35({
    1'b0, \dot_product_and_ReLU[1].product_terms[77][0] }), .in_36({1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] , 1'b0, 1'b0}), .in_37({1'b0, 
    \dot_product_and_ReLU[16].product_terms[71][0] , 1'b0}), .in_38({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] , 1'b0}), .in_39({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] , 1'b0}),
     .in_40({\dot_product_and_ReLU[7].product_terms[64][1] , 1'b0}), .in_41(
    \dot_product_and_ReLU[0].product_terms[65][0] ), .out_0({
    \level_6_sums[4][1] [9], UNCONNECTED18, UNCONNECTED17, UNCONNECTED16,  \level_6_sums[4][1] [5:0] }));
  WALLACE_CSA_DUMMY_OP61_group_359287 WALLACE_CSA_DUMMY_OP61_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[157][0] }), .in_1({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] , 
    \dot_product_and_ReLU[0].product_terms[191][1] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] }), .in_3(
    \dot_product_and_ReLU[18].product_terms[186][0] ), .in_4(
    \dot_product_and_ReLU[0].product_terms[187][0] ), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[180][0] }), .in_6({1'b0, 
    1'b0, 1'b0, 1'b0,  \level_1_sums[16][87] [2:1] }), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[171][1] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[164][0] , 1'b0}), .in_9({1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_10({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_11({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[150][0] }), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, n_1409, n_1408}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 1'b0}), .in_15({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[138][0] }), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] , 1'b0}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] }), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[183][1] }), .in_19({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[178][0] }),
     .in_20({1'b0, \dot_product_and_ReLU[0].product_terms[179][0] }), .in_21(
    \dot_product_and_ReLU[1].product_terms[176][0] ), .in_22({1'b0, 
    \dot_product_and_ReLU[0].product_terms[177][0] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[172][1] }), .in_24({
    1'b0, \dot_product_and_ReLU[8].product_terms[173][1] , 1'b0}), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[168][0] }),
     .in_26({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[169][0] , 
    1'b0}), .in_27({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] }), .in_28({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[167][0] , 1'b0}), .in_29({
    \level_1_sums[1][81][0] , 1'b0}), .in_30({
    \dot_product_and_ReLU[9].product_terms[163][0] , 1'b0}), .in_31({
    \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}), .in_32(
    \dot_product_and_ReLU[3].product_terms[161][0] ), .in_33({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[158][0] , 1'b0}), .in_34({1'b0, 
    \dot_product_and_ReLU[0].product_terms[159][1] }), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[148][0] , 1'b0}), .in_36({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[149][0] }),
     .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[144][0] }), .in_38({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] }), .in_39({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[136][1] , 1'b0}),
     .in_40({1'b0, \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}),
     .in_41({1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] }),
     .in_42({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_43({1'b0, 
    \dot_product_and_ReLU[14].product_terms[131][0] , 1'b0, 1'b0}), .in_44({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}),
     .out_0({\level_6_sums[4][2] [9], UNCONNECTED21, UNCONNECTED20, 
    UNCONNECTED19,  \level_6_sums[4][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP62_group_359293 WALLACE_CSA_DUMMY_OP62_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[72][0] }), .in_1({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] , 1'b0}),
     .in_2({1'b0, 1'b0, 1'b0, \level_6_sums[15][0] [9],  \level_6_sums[15][0] [5:0] }), .in_3({1'b0, 1'b0, 
    1'b0, \level_6_sums[15][3] [9],  \level_6_sums[15][3] [5:0] }), .in_4({
    \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_5(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[113][1] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[94][1] }), .in_10({1'b0, 
    \dot_product_and_ReLU[2].product_terms[91][1] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[86][0] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[69][1] }), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] , 1'b0}), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[186][0] }),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] }), .in_19({1'b0, 1'b0, 
    1'b0, n_1400, n_1399, \dot_product_and_ReLU[1].product_terms[176][0] }),
     .in_20({1'b0, 1'b0, 1'b0, 1'b0,  \level_1_sums[16][87] [2:1] }), .in_21({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[170][0] , 1'b0}), .in_22({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[166][0] }),
     .in_23({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[165][0] }), .in_24({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[160][1] }),
     .in_25({1'b0, 1'b0, 1'b0, 1'b0, n_1393, n_1392}), .in_26({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[156][2] , 1'b0, 1'b0}), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_28({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[148][0] }),
     .in_29({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[146][0] }), .in_30({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 1'b0}),
     .in_31({1'b0, 1'b0, 1'b0, n_1378, n_1404, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, n_1381, n_1440}), .in_33({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[128][1] }), .in_34({1'b0, 
    \dot_product_and_ReLU[4].product_terms[118][0] }), .in_35({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[119][0] }), .in_36({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] }),
     .in_37({1'b0, \dot_product_and_ReLU[1].product_terms[115][0] , 1'b0}),
     .in_38({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[111][0] , 
    1'b0}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[108][0] }), .in_40({1'b0, 
    \dot_product_and_ReLU[7].product_terms[109][1] }), .in_41({1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[107][0] }), .in_43({
    1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}), .in_44({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[105][0] , 1'b0}), .in_45({
    1'b0, \dot_product_and_ReLU[16].product_terms[102][2] }), .in_46({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[103][0] }),
     .in_47({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[100][0] }), .in_48({1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[101][1] }), .in_49(
    \dot_product_and_ReLU[4].product_terms[98][1] ), .in_50({1'b0, 
    \dot_product_and_ReLU[14].product_terms[99][0] }), .in_51({1'b0, 
    \dot_product_and_ReLU[5].product_terms[96][0] }), .in_52({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[97][0] }), .in_53({1'b0, 
    \dot_product_and_ReLU[8].product_terms[92][1] }), .in_54({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_55({1'b0, 
    \dot_product_and_ReLU[1].product_terms[85][0] , 1'b0}), .in_56({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}), .in_57({1'b0, 
    \dot_product_and_ReLU[10].product_terms[80][0] }), .in_58({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }), .in_59({1'b0, 
    1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] }), .in_60({1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_61({
    \dot_product_and_ReLU[2].product_terms[70][0] , 1'b0}), .in_62({
    \dot_product_and_ReLU[16].product_terms[71][0] , 1'b0}), .in_63({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[64][1] }), .in_64({1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] }), .in_65({1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] }), .in_66({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }), .in_67(
    \dot_product_and_ReLU[3].product_terms[184][1] ), .in_68(
    \dot_product_and_ReLU[5].product_terms[185][0] ), .in_69({1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] }), .in_70({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[181][0] , 1'b0}), .in_71({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[178][0] , 1'b0}),
     .in_72({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[179][0] }), .in_73({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[172][1] , 1'b0}), .in_74({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] }),
     .in_75({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[169][0] }), .in_76({1'b0, 1'b0, 
    1'b0, 1'b0, \level_1_sums[1][81][0] }), .in_77({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] }), .in_78({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[152][0] , 1'b0}), .in_79({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }),
     .in_80({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[151][0] }), .in_81({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }), .in_82({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 1'b0}),
     .in_83({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[143][0] , 
    1'b0}), .in_84({1'b0, \dot_product_and_ReLU[17].product_terms[140] [0]}),
     .in_85(\dot_product_and_ReLU[0].product_terms[141][0] ), .in_86({1'b0, 
    \dot_product_and_ReLU[1].product_terms[137][0] }), .in_87({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[134][1] , 1'b0}), .in_88({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[135][0] , 1'b0}),
     .out_0({\level_8_sums[15] [8], UNCONNECTED22,  \level_8_sums[15] [7:0] }));
  WALLACE_CSA_DUMMY_OP70_group_106217 WALLACE_CSA_DUMMY_OP70_groupi(.in_0({1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0}), .in_1({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[31][1] }), .in_2({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[11][1] }), .in_3({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] , 1'b0}),
     .in_4({1'b0, 1'b0, 1'b0, \level_6_sums[11][3] [9],  \level_6_sums[11][3] [5:0] }), .in_5({1'b0, 1'b0, 
    \level_6_sums[11][2] [9],  \level_6_sums[11][2] [6:0] }), .in_6({1'b0, 1'b0, 1'b0, 
    \level_4_sums[11][5] [8],  \level_4_sums[11][5] [4:0] }), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1427, n_1426, 
    1'b0}), .in_8({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0, 1'b0}), .in_9({
    1'b0, 1'b0, 1'b0, 1'b0, n_2925_danc, n_2926_danc}), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[112][2] }), .in_12({1'b0, 1'b0, 
    n_2866_danc, n_2867_danc, \dot_product_and_ReLU[1].product_terms[77][0] , 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] }), .in_14({1'b0, 
    1'b0, 1'b0, 1'b0, n_1465, n_2773_danc}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] }),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[49][0] }), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[46][2] }), .in_19({
    1'b0, 1'b0, 1'b0, n_2950_danc, n_1414, 
    \dot_product_and_ReLU[8].product_terms[36][0] }), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[29][0] }), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[27][0] , 1'b0}),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[18][0] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }), .in_24({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[14][1] , 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_25({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[16].product_terms[12][0] , 
    \dot_product_and_ReLU[0].product_terms[13][0] }), .in_26({1'b0, 1'b0, 1'b0, 
    n_1471, n_1470, n_1469}), .in_27({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_28({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[126][1] }), .in_29({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] , 1'b0}),
     .in_30({1'b0, \dot_product_and_ReLU[0].product_terms[122][0] }), .in_31({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[123][1] }),
     .in_32(\dot_product_and_ReLU[2].product_terms[116][0] ), .in_33(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .in_34(
    \dot_product_and_ReLU[0].product_terms[114][1] ), .in_35({
    \dot_product_and_ReLU[1].product_terms[115][0] , 1'b0}), .in_36({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[107][0] }), .in_37({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}),
     .in_38({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_39({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[16].product_terms[102][2] , 1'b0}), .in_40({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[103][0] }),
     .in_41({1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[100][0] }),
     .in_42({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[101][1] }), .in_43({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[98][1] , 1'b0}), .in_44({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] }),
     .in_45({\dot_product_and_ReLU[5].product_terms[96][0] , 1'b0}), .in_46({
    \dot_product_and_ReLU[4].product_terms[97][0] , 1'b0}), .in_47({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }), .in_48({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[79][0] , 1'b0}),
     .in_49({1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] , 1'b0}), .in_50({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[75][0] , 1'b0}), .in_51({
    1'b0, \dot_product_and_ReLU[1].product_terms[73][0] , 1'b0, 1'b0}), .in_52({
    1'b0, \dot_product_and_ReLU[2].product_terms[70][0] }), .in_53({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[71][0] }), .in_54({
    \dot_product_and_ReLU[4].product_terms[68][0] , 1'b0}), .in_55({
    \dot_product_and_ReLU[1].product_terms[69][1] , 1'b0}), .in_56({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[65][0] , 1'b0}), .in_57({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}), .in_58({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[63][1] }),
     .in_59({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[60][2] }), .in_60({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[15].product_terms[61][1] }), .in_61({
    \dot_product_and_ReLU[1].product_terms[56][1] , 1'b0}), .in_62(
    \dot_product_and_ReLU[7].product_terms[57][2] ), .in_63({
    \dot_product_and_ReLU[2].product_terms[44][1] , 1'b0}), .in_64(
    \dot_product_and_ReLU[3].product_terms[45][1] ), .in_65({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[40][0] , 1'b0}), .in_66({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[41][0] , 1'b0}), .in_67({1'b0, 
    \dot_product_and_ReLU[2].product_terms[34][0] }), .in_68({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[35][0] }), .in_69({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[32][1] , 1'b0}), .in_70({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }), .in_71({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] }),
     .in_72({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[25][0] }), .in_73({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] }), .in_74({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_75({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[20][0] }), .in_76({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }),
     .in_77({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] }), .in_78({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[9][0] , 1'b0}), .in_79({1'b0, 
    \dot_product_and_ReLU[7].product_terms[7][0] }), .in_80({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0, 1'b0}), .in_81({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[1][0] , 1'b0}), .out_0({ \level_8_sums[11] [9:0] }));
  WALLACE_CSA_DUMMY_OP74_group_109823 WALLACE_CSA_DUMMY_OP74_groupi(.in_0({1'b0, 
    B[228], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_2({1'b0, 1'b0, 
    1'b0, \level_6_sums[10][2] [9],  \level_6_sums[10][2] [5:0] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, n_1503, 
    n_1525}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, B[248], 1'b0}), .in_5({1'b0, 1'b0, 
    1'b0, 1'b0, n_1496, n_1495}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[244]}),
     .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1488, n_1553}), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[236]}), .in_9({1'b0, 1'b0, 1'b0, n_1550, n_1549, 1'b0}),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[224]}), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, B[223], 1'b0}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, B[219], 1'b0}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, B[216], 1'b0}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, n_1504, n_1529}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[204]}),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[200]}), .in_17({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[198]}), .in_18({1'b0, 1'b0, 1'b0, n_1486, n_1539, 1'b0}),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, n_1508, n_1527}), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[193]}), .in_21({1'b0, B[252]}), .in_22({1'b0, 1'b0, 1'b0, 
    1'b0, B[253]}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_24({1'b0, 
    B[241]}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, B[239]}), .in_26({1'b0, B[230]}),
     .in_27({1'b0, 1'b0, 1'b0, 1'b0, B[231]}), .in_28({1'b0, B[226], 1'b0}),
     .in_29({1'b0, 1'b0, 1'b0, 1'b0, B[227]}), .in_30({1'b0, 1'b0, B[220]}),
     .in_31({1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_32({1'b0, B[215], 1'b0}),
     .in_33({1'b0, B[212], 1'b0}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[213]}),
     .in_35({1'b0, B[208]}), .in_36({1'b0, 1'b0, 1'b0, B[209], 1'b0}), .in_37(
    B[206]), .in_38(B[207]), .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[202]}), .in_40({
    1'b0, B[203]}), .out_0({\level_7_sums[10][1] [9], UNCONNECTED24, 
    UNCONNECTED23,  \level_7_sums[10][1] [6:0] }));
  WALLACE_CSA_DUMMY_OP75_group_109813_6325 WALLACE_CSA_DUMMY_OP75_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[205]}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[251], 1'b0}), .in_2({1'b0, 1'b0, 1'b0, n_1518, n_1534, B[255]}), .in_3({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[252]}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    n_1496, n_1495}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1531, n_1553}), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_7({1'b0, 1'b0, 1'b0, B[239], 1'b0}),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[235]}), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[233]}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, B[230], 1'b0}),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1214, n_1547}), .in_12({1'b0, 1'b0, 1'b0, 
    n_1487, n_2602_danc, n_2603_danc}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, n_1497, 
    n_1513}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, B[218], 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, n_1530, n_1529}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[207]}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, B[202], 1'b0}), .in_18({1'b0, 
    1'b0, 1'b0, 1'b0, B[200], 1'b0}), .in_19({1'b0, 1'b0, 1'b0, n_1528, n_1508, 
    n_1527}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[193]}), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, B[244]}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, B[245]}),
     .in_23({1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_24({1'b0, 1'b0, 1'b0, 1'b0, 
    B[241]}), .in_25({1'b0, 1'b0, B[229]}), .in_26({1'b0, 1'b0, 1'b0, B[226], 
    1'b0}), .in_27({1'b0, 1'b0, 1'b0, 1'b0, B[227]}), .in_28({1'b0, 1'b0, 1'b0, 
    1'b0, B[216]}), .in_29({1'b0, B[217]}), .in_30({1'b0, B[215]}), .in_31({
    1'b0, 1'b0, B[212], 1'b0, 1'b0}), .in_32({1'b0, 1'b0, 1'b0, 1'b0, B[213]}),
     .in_33({1'b0, B[208]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[209]}), .in_35({
    1'b0, 1'b0, 1'b0, B[198], 1'b0}), .in_36({1'b0, 1'b0, B[199]}), .in_37(
    B[196]), .in_38({B[197], 1'b0}), .out_0({\level_6_sums[11][3] [9], 
    UNCONNECTED27, UNCONNECTED26, UNCONNECTED25,  \level_6_sums[11][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP75_group_109813 WALLACE_CSA_DUMMY_OP75_groupi4121(.in_0({
    1'b0, \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[7][0] }), .in_3({1'b0, 1'b0, 1'b0, 
    1'b0, n_1216, n_1492}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[11].product_terms[50][0] , 1'b0}), .in_5({1'b0, 1'b0, 
    1'b0, 1'b0, n_1485, n_2818_danc}), .in_6({1'b0, 1'b0, n_2822_danc, 
    n_2823_danc, \dot_product_and_ReLU[6].product_terms[43][0] , 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, n_2929_danc, n_2780_danc}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[38][1] , 1'b0}), .in_9({1'b0, 1'b0, 
    1'b0, n_1405, n_1414, \dot_product_and_ReLU[2].product_terms[37][1] }),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[32][1] , 
    \dot_product_and_ReLU[2].product_terms[33][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[28][0] , 
    \dot_product_and_ReLU[0].product_terms[29][0] }), .in_12({1'b0, 1'b0, 1'b0, 
    n_2996_danc, n_2976_danc, \dot_product_and_ReLU[0].product_terms[27][0] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[24][0] }), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, n_1482, n_2788_danc}), .in_16({1'b0, 1'b0, 1'b0, 
    n_2980_danc, n_2981_danc, \dot_product_and_ReLU[1].product_terms[11][1] }),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[9][0] }), .in_18({1'b0, 
    \dot_product_and_ReLU[19].product_terms[60][2] }), .in_19({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[15].product_terms[61][1] , 1'b0}), .in_20({
    1'b0, \dot_product_and_ReLU[7].product_terms[58][0] , 1'b0, 1'b0}), .in_21({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[59][1] }),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] }), .in_23({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[53][1] }), .in_24({1'b0, 
    \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}), .in_25({1'b0, 
    \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0}), .in_26({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[34][0] , 1'b0}), .in_27({1'b0, 
    \dot_product_and_ReLU[2].product_terms[35][0] }), .in_28({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[31][1] }), .in_29({1'b0, 
    \dot_product_and_ReLU[4].product_terms[20][0] }), .in_30({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }), .in_32({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_34({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[16].product_terms[12][0] }), .in_35({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] , 1'b0}), .in_36({
    1'b0, \dot_product_and_ReLU[19].product_terms[2][0] , 1'b0}), .in_37({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[3][0] , 1'b0}), .in_38({
    1'b0, \dot_product_and_ReLU[4].product_terms[1][0] , 1'b0}), .out_0({
    \level_6_sums[15][0] [9], UNCONNECTED30, UNCONNECTED29, UNCONNECTED28,  \level_6_sums[15][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP78_group_359273 WALLACE_CSA_DUMMY_OP78_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[175][0] }), .in_1({
    \level_1_sums[1][81][0] , 1'b0}), .in_2({1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] }), .in_3({1'b0, 1'b0, 1'b0, 
    1'b0, \level_3_sums[10][22][3] , \level_3_sums[10][22][2] , 
    \level_3_sums[10][22][1] , \level_3_sums[10][22][0] }), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] }), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[186][0] }),
     .in_6({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 
    1'b0}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[10].product_terms[172][1] , 1'b0}), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, n_1453, n_1452}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[168][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[155][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[152][0] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[149][0] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[2][73] [2], 
    \level_1_sums[2][73] [0]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[142][0] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 1'b0}),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[136][1] , 1'b0}), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[133][0] }),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[131][0] }), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }),
     .in_20(\dot_product_and_ReLU[6].product_terms[188][1] ), .in_21(
    \dot_product_and_ReLU[0].product_terms[189][0] ), .in_22({
    \dot_product_and_ReLU[4].product_terms[166][0] , 1'b0}), .in_23(
    \dot_product_and_ReLU[0].product_terms[167][0] ), .in_24({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[165][0] }), .in_25({1'b0, 
    \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0}), .in_26({1'b0, 
    \dot_product_and_ReLU[0].product_terms[157][0] , 1'b0}), .in_27({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[150][0] }),
     .in_28({1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }), .in_29({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[145][1] }), .in_31({1'b0, 
    \dot_product_and_ReLU[8].product_terms[139][0] , 1'b0}), .in_32({1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[135][0] }), .out_0({
    \level_6_sums[10][2] [9], UNCONNECTED33, UNCONNECTED32, UNCONNECTED31,  \level_6_sums[10][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP82_group_359272 WALLACE_CSA_DUMMY_OP82_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[152][0] }), .in_1({
    1'b0, \dot_product_and_ReLU[18].product_terms[153][0] , 1'b0}), .in_2({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[146][0] }), .in_3({1'b0, 1'b0, 1'b0, 
    1'b0, n_1387, n_1390}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[143][0] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, n_1441, n_1440}), .in_6({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[159][1] }), .in_7({1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[156][2] }), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[157][0] }), .in_9(
    \dot_product_and_ReLU[14].product_terms[154][0] ), .in_10(
    \dot_product_and_ReLU[0].product_terms[155][0] ), .in_11({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[148][0] , 1'b0}), .in_12({1'b0, 
    \dot_product_and_ReLU[1].product_terms[149][0] , 1'b0}), .in_13({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0]}),
     .in_14({1'b0, \dot_product_and_ReLU[0].product_terms[141][0] }), .in_15(
    \dot_product_and_ReLU[19].product_terms[138][0] ), .in_16(
    \dot_product_and_ReLU[8].product_terms[139][0] ), .in_17({1'b0, 
    \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}), .in_18({1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] , 1'b0}), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[135][0] }),
     .in_20({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_21({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[128][1] , 1'b0}), .in_22({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}),
     .out_0({\level_5_sums[9][4] [9], UNCONNECTED37, UNCONNECTED36, 
    UNCONNECTED35, UNCONNECTED34,  \level_5_sums[9][4] [4:0] }));
  WALLACE_CSA_DUMMY_OP86_group_109840 WALLACE_CSA_DUMMY_OP86_groupi(.in_0({1'b0, 
    1'b0, 1'b0, B[210], 1'b0}), .in_1({1'b0, B[211], 1'b0}), .in_2({1'b0, 1'b0, 
    1'b0, \level_6_sums[2][1] [9],  \level_6_sums[2][1] [5:0] }), .in_3({1'b0, 1'b0, 
    \level_6_sums[2][0] [9],  \level_6_sums[2][0] [6:0] }), .in_4({1'b0, 1'b0, 1'b0, 
    \level_3_sums[2][21] [7],  \level_3_sums[2][21] [3:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0,  \level_3_sums[2][17] [3:0] }), .in_6({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[251], B[250]}), .in_7({1'b0, 1'b0, 1'b0, 
    \level_2_sums[2][45] [6],  \level_2_sums[2][45] [2:1] , \level_3_sums[19][22][0] }), .in_8({1'b0, 1'b0, 
    1'b0, \level_2_sums[2][41] [6],  \level_2_sums[2][41] [2:0] }), .in_9({1'b0, 1'b0, 1'b0, 
    \level_2_sums[2][32] [6],  \level_2_sums[2][32] [2:0] }), .in_10({1'b0, 1'b0, 1'b0, 1'b0, B[254], 1'b0}),
     .in_11({1'b0, 1'b0, n_1554, n_1553,  B[242:243] }), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[240]}), .in_13({1'b0, 1'b0, 1'b0, B[236], 1'b0, 1'b0}), .in_14({1'b0, 
    1'b0, n_1552, n_1551, 1'b0, B[235]}), .in_15({1'b0, 1'b0, 1'b0, n_1550, 
    n_1549, B[232]}), .in_16({1'b0, 1'b0, 1'b0, B[228], 1'b0, 1'b0}), .in_17({
    1'b0, 1'b0, 1'b0, 1'b0, n_1548, n_1547}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, B[222]}), .in_19({1'b0, 1'b0, 1'b0, n_1546, n_1545, B[218]}), .in_20({
    1'b0, 1'b0, 1'b0, n_1544, n_1543, B[216]}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, B[209]}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, n_1542, n_1541}), .in_23({
    1'b0, 1'b0, 1'b0, n_1540, n_1539}), .in_24({1'b0, 1'b0, 1'b0, 1'b0, n_1538, 
    \level_1_sums[12][95] [0]}), .in_25(
    \dot_product_and_ReLU[18].product_terms[186][0] ), .in_26(
    \dot_product_and_ReLU[0].product_terms[187][0] ), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, n_1537, n_1536}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[156][2] }), .in_29({1'b0, 1'b0, 
    1'b0,  \level_1_sums[2][73] [2:0] }), .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] , 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] }),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, B[252]}), .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    B[253]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[247]}), .in_35({1'b0, 1'b0, 
    B[244], 1'b0, 1'b0}), .in_36({1'b0, 1'b0, 1'b0, 1'b0, B[245]}), .in_37({
    1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_38({1'b0, B[239]}), .in_39({1'b0, 
    1'b0, 1'b0, 1'b0, B[230]}), .in_40({1'b0, 1'b0, 1'b0, B[231], 1'b0}),
     .in_41({1'b0, B[226]}), .in_42({1'b0, 1'b0, 1'b0, 1'b0, B[227]}), .in_43({
    1'b0, B[220]}), .in_44(B[221]), .in_45({1'b0, 1'b0, 1'b0, 1'b0, B[214]}),
     .in_46({1'b0, 1'b0, 1'b0, B[215], 1'b0}), .in_47({1'b0, 1'b0, 1'b0, 1'b0, 
    B[213]}), .in_48({1'b0, B[206]}), .in_49({1'b0, 1'b0, 1'b0, 1'b0, B[207]}),
     .in_50({1'b0, 1'b0, B[203]}), .in_51({1'b0, 1'b0, 1'b0, B[200], 1'b0}),
     .in_52({1'b0, 1'b0, B[201]}), .in_53({B[194], 1'b0}), .in_54({B[195], 1'b0}),
     .in_55({1'b0, B[192], 1'b0}), .in_56({1'b0, 1'b0, 1'b0, 1'b0, B[193]}),
     .in_57({1'b0, \dot_product_and_ReLU[6].product_terms[188][1] }), .in_58({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }),
     .in_59({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[176][0] }), .in_60({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[177][0] , 1'b0}), .in_61({
    1'b0, \dot_product_and_ReLU[9].product_terms[163][0] }), .in_62({1'b0, 
    \dot_product_and_ReLU[3].product_terms[161][0] , 1'b0, 1'b0}), .in_63({
    1'b0, \dot_product_and_ReLU[1].product_terms[158][0] , 1'b0}), .in_64({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[159][1] }),
     .in_65(\dot_product_and_ReLU[14].product_terms[154][0] ), .in_66({
    \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_67({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }), .in_68({
    \dot_product_and_ReLU[1].product_terms[148][0] , 1'b0}), .in_69(
    \dot_product_and_ReLU[1].product_terms[149][0] ), .in_70({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }), .in_71({1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[145][1] }), .out_0({ \final_sums[2] [9:0] }));
  WALLACE_CSA_DUMMY_OP89_group_106209 WALLACE_CSA_DUMMY_OP89_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }), .in_1({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[19][1] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[4][1] [9],  \level_6_sums[4][1] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_1467, 
    n_1466}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[62][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, n_1465, n_2773_danc}), .in_7({1'b0, 1'b0, 1'b0, n_1216, n_1468, 
    n_1492}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_9({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[44][1] , 1'b0, 1'b0}), .in_10({1'b0, 
    1'b0, n_2822_danc, n_2823_danc, 
    \dot_product_and_ReLU[6].product_terms[43][0] , 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[40][0] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[26][2] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, n_1464, n_1463}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }), .in_15({1'b0, 
    1'b0, 1'b0, n_1462, n_1480, \dot_product_and_ReLU[7].product_terms[7][0] }),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, n_1461, n_2757_danc}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[60][2] }), .in_18({
    1'b0, \dot_product_and_ReLU[15].product_terms[61][1] , 1'b0}), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[54][0] }), .in_20({
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] , 1'b0, 1'b0}),
     .in_21({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] , 
    1'b0}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[53][1] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] }), .in_24({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[48][1] }),
     .in_25({1'b0, \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[37][1] }), .in_27({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[34][0] , 1'b0}), .in_28({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[35][0] }), .in_29({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] , 1'b0}), .in_30({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] , 1'b0}),
     .in_31({1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[31][1] }), .in_33({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[28][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[0].product_terms[29][0] , 1'b0}), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[23][0] , 1'b0}), .in_36({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[20][0] }), .in_37({
    1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }), .in_38({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[10][0] }), .in_39({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[11][1] }), .in_40({
    1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_41({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[9][0] }), .in_42({1'b0, 
    \dot_product_and_ReLU[4].product_terms[3][0] }), .out_0({
    \level_7_sums[4][0] [9], UNCONNECTED39, UNCONNECTED38,  \level_7_sums[4][0] [6:0] }));
  WALLACE_CSA_DUMMY_OP91_group_109814 WALLACE_CSA_DUMMY_OP91_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, B[227]}), .in_1({1'b0, 1'b0, 1'b0, B[193], 1'b0}), .in_2({
    1'b0, 1'b0, \level_7_sums[14][0] [9],  \level_7_sums[14][0] [6:0] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[14][2] [9],  \level_6_sums[14][2] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[246]}), .in_5({1'b0, 1'b0, 1'b0, n_1209, n_1518, n_1534}), .in_6({1'b0, 
    1'b0, 1'b0, 1'b0, B[243], 1'b0}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1517, 
    n_1516}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[236]}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, n_1515, n_1549}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, n_1524, 
    n_1523}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, n_1514, n_1513}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[216]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[214]}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[210]}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, n_1512, 
    n_1511}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, n_1542, n_1541}), .in_18({1'b0, 
    1'b0, 1'b0, n_1510, n_1509, B[201]}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    B[198]}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, B[196]}), .in_21({1'b0, 1'b0, 
    1'b0, n_1508, n_1507, n_1527}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, B[252]}),
     .in_23({1'b0, B[253], 1'b0}), .in_24({1'b0, B[250]}), .in_25({1'b0, 1'b0, 
    1'b0, 1'b0, B[251]}), .in_26({1'b0, 1'b0, 1'b0, B[248], 1'b0}), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, B[249]}), .in_28({1'b0, B[240]}), .in_29({1'b0, 
    1'b0, 1'b0, B[241], 1'b0}), .in_30({1'b0, B[234]}), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, B[235]}), .in_32(B[228]), .in_33(B[229]), .in_34({1'b0, 1'b0, 
    1'b0, 1'b0, B[224]}), .in_35({1'b0, 1'b0, 1'b0, 1'b0, B[225]}), .in_36({
    B[218], 1'b0}), .in_37(B[219]), .in_38({1'b0, 1'b0, 1'b0, 1'b0, B[213]}),
     .in_39({1'b0, 1'b0, B[208]}), .in_40({1'b0, 1'b0, 1'b0, 1'b0, B[209]}),
     .in_41(B[202]), .in_42({1'b0, B[203]}), .out_0({ \final_sums[14] [9:0] }));
  WALLACE_CSA_DUMMY_OP93_group_109834 WALLACE_CSA_DUMMY_OP93_groupi(.in_0({1'b0, 
    \level_7_sums[17][0] [9],  \level_7_sums[17][0] [7:0] }), .in_1({1'b0, 1'b0, 1'b0, 
    \level_6_sums[17][2] [9],  \level_6_sums[17][2] [5:0] }), .in_2({1'b0, 1'b0, 1'b0, 1'b0, n_1506, n_1534}),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, B[246], 1'b0}), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[245]}), .in_5({1'b0, 1'b0, 1'b0, 1'b0,  B[240:241] }), .in_6({1'b0, 1'b0, 
    B[219]}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[215]}), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[207]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, B[204], 1'b0}),
     .in_10({1'b0, 1'b0, 1'b0, n_1510, n_1509, B[201]}), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[196]}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1508, n_1527}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[192]}), .in_14(B[252]), .in_15({
    B[253], 1'b0}), .in_16({B[250], 1'b0}), .in_17({1'b0, B[251]}), .in_18({
    1'b0, 1'b0, 1'b0, B[248], 1'b0}), .in_19({1'b0, 1'b0, B[249], 1'b0, 1'b0}),
     .in_20({1'b0, 1'b0, 1'b0, B[238], 1'b0}), .in_21({1'b0, B[239]}), .in_22(
    B[236]), .in_23({B[237], 1'b0, 1'b0}), .in_24(B[234]), .in_25({B[235], 1'b0}),
     .in_26(B[232]), .in_27({B[233], 1'b0}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, 
    B[230]}), .in_29({1'b0, B[231]}), .in_30({1'b0, B[229], 1'b0}), .in_31({
    1'b0, B[224]}), .in_32({1'b0, 1'b0, 1'b0, B[225], 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, B[222]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_35({
    1'b0, 1'b0, 1'b0, B[220], 1'b0}), .in_36({1'b0, B[221]}), .in_37({1'b0, 
    B[212], 1'b0}), .in_38({1'b0, 1'b0, 1'b0, B[213], 1'b0}), .in_39({1'b0, 
    1'b0, 1'b0, 1'b0, B[211]}), .in_40({1'b0, 1'b0, 1'b0, B[208]}), .in_41({
    1'b0, 1'b0, 1'b0, 1'b0, B[209]}), .in_42({1'b0, B[203], 1'b0}), .in_43({
    1'b0, 1'b0, 1'b0, 1'b0, B[199]}), .out_0({ \final_sums[17] [9:0] }));
  WALLACE_CSA_DUMMY_OP95_group_109821 WALLACE_CSA_DUMMY_OP95_groupi(.in_0({1'b0, 
    1'b0, 1'b0, B[193], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[241]}), .in_2({
    1'b0, 1'b0, 1'b0, n_1518, n_1534, B[255]}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, B[250]}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[248]}), .in_5({1'b0, 
    1'b0, 1'b0, 1'b0,  B[244:245] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, B[239], B[238]}), .in_7({
    1'b0, 1'b0, 1'b0, 1'b0, B[237], 1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0,  B[234:235] }),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[230]}), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[228]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1505, n_1521}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[224]}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[222]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[220]}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[216]}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, n_1504, n_1529}), .in_17({1'b0, 1'b0, 1'b0, n_1520, n_1519, B[208]}),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0,  B[200:201] }), .in_19({1'b0, 1'b0, 1'b0, B[252], 1'b0}),
     .in_20({1'b0, B[253]}), .in_21({B[246], 1'b0}), .in_22(B[247]), .in_23({
    1'b0, 1'b0, 1'b0, 1'b0, B[242]}), .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[243]}),
     .in_25({1'b0, 1'b0, 1'b0, B[232], 1'b0}), .in_26({1'b0, B[233]}), .in_27({
    1'b0, B[219]}), .in_28({1'b0, B[212]}), .in_29({1'b0, 1'b0, 1'b0, B[213], 
    1'b0}), .in_30({1'b0, B[204]}), .in_31({1'b0, 1'b0, 1'b0, B[205], 1'b0}),
     .in_32(B[202]), .in_33(B[203]), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[199]}),
     .in_35({1'b0, B[196]}), .in_36({1'b0, 1'b0, B[197], 1'b0, 1'b0}), .in_37({
    1'b0, 1'b0, 1'b0, B[194], 1'b0}), .in_38({1'b0, 1'b0, 1'b0, 1'b0, B[195]}),
     .out_0({\level_6_sums[0][3] [9], UNCONNECTED42, UNCONNECTED41, 
    UNCONNECTED40,  \level_6_sums[0][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP98_group_359290 WALLACE_CSA_DUMMY_OP98_groupi(.in_0({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[71][0] }), .in_1({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] , 1'b0}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[69][1] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[16][0] [9],  \level_6_sums[16][0] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 
    \level_6_sums[16][3] [9],  \level_6_sums[16][3] [5:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[16][10][7] , \level_4_sums[16][10][3] , 
    \level_4_sums[16][10][2] , \level_4_sums[16][10][1] , 
    \level_4_sums[16][10][0] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0,  \level_3_sums[16][15] [3:0] }), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 
    1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[118][0] , 1'b0}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[117][0] , 1'b0}),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }), .in_12({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[111][0] , 
    \dot_product_and_ReLU[3].product_terms[110][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[94][1] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 
    \dot_product_and_ReLU[0].product_terms[88][1] }), .in_16({1'b0, 1'b0, 1'b0, 
    n_2866_danc, n_1215, n_2867_danc}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \level_1_sums[4][37][1] }), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[73][0] }), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }), .in_20({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[186][0] }), .in_21({1'b0, 1'b0, 
    1'b0, n_1415, \level_1_sums[7][92] [0], 
    \dot_product_and_ReLU[5].product_terms[185][0] }), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[182][0] }),
     .in_23({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[155][0] }), .in_24({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] , 
    \dot_product_and_ReLU[9].product_terms[152][0] }), .in_25({1'b0, 
    \dot_product_and_ReLU[0].product_terms[150][0] }), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, n_1389, n_1408}), .in_28({1'b0, 1'b0, 1'b0, n_1380, 
    n_1379, \dot_product_and_ReLU[17].product_terms[140] [0]}), .in_29({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] }),
     .in_30(\dot_product_and_ReLU[1].product_terms[108][0] ), .in_31(
    \dot_product_and_ReLU[7].product_terms[109][1] ), .in_32({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] , 1'b0}), .in_33({1'b0, 
    1'b0, \dot_product_and_ReLU[16].product_terms[107][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_35({1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[102][2] , 1'b0, 1'b0}), .in_36({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[103][0] }),
     .in_37(\dot_product_and_ReLU[0].product_terms[100][0] ), .in_38({
    \dot_product_and_ReLU[4].product_terms[101][1] , 1'b0}), .in_39(
    \dot_product_and_ReLU[5].product_terms[96][0] ), .in_40(
    \dot_product_and_ReLU[4].product_terms[97][0] ), .in_41({
    \dot_product_and_ReLU[8].product_terms[92][1] , 1'b0}), .in_42(
    \dot_product_and_ReLU[0].product_terms[93][0] ), .in_43({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[86][0] }), .in_44({1'b0, 
    \dot_product_and_ReLU[12].product_terms[87][0] , 1'b0}), .in_45({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] }), .in_46({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[85][0] }),
     .in_47({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[82][0] }), .in_48({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }), .in_49({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[80][0] , 1'b0}), .in_50({
    1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }), .in_51({1'b0, 
    \dot_product_and_ReLU[10].product_terms[78][1] }), .in_52({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[79][0] }), .in_53({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[66][0] , 1'b0}), .in_54({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }),
     .in_55({1'b0, \dot_product_and_ReLU[7].product_terms[64][1] }), .in_56({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[65][0] , 1'b0}),
     .in_57({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] , 
    1'b0}), .in_58({1'b0, \dot_product_and_ReLU[0].product_terms[191][1] }),
     .in_59({1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[181][0] }),
     .in_60({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[178][0] , 
    1'b0}), .in_61({1'b0, \dot_product_and_ReLU[0].product_terms[179][0] }),
     .in_62(\dot_product_and_ReLU[1].product_terms[176][0] ), .in_63({
    \dot_product_and_ReLU[0].product_terms[177][0] , 1'b0}), .in_64({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[158][0] }), .in_65({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0}),
     .in_66({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[156][2] }), .in_67({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[157][0] , 1'b0}), .in_68({
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[147][0] }), .in_69({1'b0, 
    \dot_product_and_ReLU[0].product_terms[145][1] }), .in_70({1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] }), .in_71({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[135][0] , 1'b0}), .in_72({
    1'b0, \dot_product_and_ReLU[0].product_terms[130][0] , 1'b0}), .in_73({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[131][0] }),
     .in_74({1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}),
     .out_0({\level_8_sums[16][8] , UNCONNECTED43, \level_8_sums[16][7] , 
    \level_8_sums[16][6] , \level_8_sums[16][5] , \level_8_sums[16][4] , 
    \level_8_sums[16][3] , \level_8_sums[16][2] , \level_8_sums[16][1] , 
    \level_8_sums[16][0] }));
  WALLACE_CSA_DUMMY_OP99_group_106220 WALLACE_CSA_DUMMY_OP99_groupi(.in_0({1'b0, 
    \dot_product_and_ReLU[0].product_terms[28][0] , 1'b0}), .in_1({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[29][0] , 1'b0}), .in_2({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[27][0] }), .in_3({
    1'b0, \level_7_sums[8][1] [9],  \level_7_sums[8][1] [7:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[125][1] , 
    \dot_product_and_ReLU[17].product_terms[124][0] }), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[122][0] }), .in_7({
    1'b0, 1'b0, 1'b0, \level_1_sums[8][55] [4],  \level_1_sums[8][55] [1:0] }), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[106][0] }), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[100][0] }),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[98][1] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[86][0] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] }),
     .in_13({1'b0, 1'b0, 1'b0, n_2862_danc, n_1436, 1'b0}), .in_14({1'b0, 1'b0, 
    n_2866_danc, n_2867_danc, \dot_product_and_ReLU[1].product_terms[77][0] , 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, n_2870_danc, n_2871_danc}), .in_16({1'b0, 1'b0, 1'b0, n_2772_danc, 
    n_2773_danc, \dot_product_and_ReLU[7].product_terms[58][0] }), .in_17({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] , n_1433, 
    n_1432}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[42][1] }), .in_20({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[34][0] }), .in_21({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[32][1] , 1'b0}), .in_22({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }),
     .in_23({1'b0, 1'b0, 1'b0, 1'b0, n_1464, n_1463}), .in_24({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[19][1] , 1'b0}), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] }), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[13][0] , 1'b0}), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, n_1431, n_1430}), .in_29({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[4][0] }), .in_30({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[120][1] , 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[121][1] }),
     .in_32({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] , 
    1'b0}), .in_33({1'b0, \dot_product_and_ReLU[0].product_terms[119][0] }),
     .in_34({1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }), .in_35({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}),
     .in_36({1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }), .in_37({
    1'b0, \dot_product_and_ReLU[17].product_terms[112][2] }), .in_38({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[113][1] , 1'b0}),
     .in_39({1'b0, \dot_product_and_ReLU[7].product_terms[109][1] }), .in_40({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1], 1'b0}),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[103][0] }), .in_43({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[96][0] , 1'b0}),
     .in_44({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[97][0] , 
    1'b0}), .in_45({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[94][1] }), .in_46({1'b0, 
    \dot_product_and_ReLU[2].product_terms[95][0] }), .in_47({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[92][1] , 1'b0}), .in_48({1'b0, 
    \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_49({1'b0, 
    \dot_product_and_ReLU[0].product_terms[90][0] }), .in_50({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_51({1'b0, 
    \dot_product_and_ReLU[0].product_terms[88][1] }), .in_52({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] }), .in_53({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[82][0] , 1'b0}), .in_54({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}),
     .in_55({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[78][1] , 
    1'b0}), .in_56({1'b0, \dot_product_and_ReLU[4].product_terms[79][0] }),
     .in_57({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_58({1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[72][0] , 1'b0, 1'b0}), .in_59({1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[73][0] , 1'b0, 1'b0}), .in_60({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[71][0] }),
     .in_61({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[67][0] }), .in_62({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[64][1] }), .in_63({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] }), .in_64({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}), .in_65({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[63][1] , 1'b0}), .in_66({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[15].product_terms[61][1] }),
     .in_67({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[56][1] }), .in_68({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0}), .in_69({1'b0, 
    \dot_product_and_ReLU[17].product_terms[53][1] , 1'b0}), .in_70({1'b0, 
    \dot_product_and_ReLU[19].product_terms[48][1] }), .in_71({
    \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}), .in_72({1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_73({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[47][1] }), .in_74({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] }), .in_75({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[45][1] }),
     .in_76({1'b0, \dot_product_and_ReLU[2].product_terms[40][0] }), .in_77({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[41][0] }),
     .in_78(\dot_product_and_ReLU[7].product_terms[38][1] ), .in_79(
    \dot_product_and_ReLU[0].product_terms[39][0] ), .in_80(
    \dot_product_and_ReLU[8].product_terms[36][0] ), .in_81(
    \dot_product_and_ReLU[2].product_terms[37][1] ), .in_82({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_83({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_84({1'b0, 
    \dot_product_and_ReLU[4].product_terms[20][0] , 1'b0}), .in_85({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}), .in_86({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[10][0] , 1'b0}), .in_87({
    1'b0, \dot_product_and_ReLU[1].product_terms[11][1] }), .in_88({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[7][0] , 1'b0}), .in_89({1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] , 1'b0}), .in_90({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[3][0] }), .in_91({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] }), .in_92(
    \dot_product_and_ReLU[4].product_terms[1][0] ), .out_0({ \level_8_sums[8] [9:0] }));
  WALLACE_CSA_DUMMY_OP102_group_106219 WALLACE_CSA_DUMMY_OP102_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }),
     .in_1({1'b0, 1'b0, 1'b0, \level_6_sums[13][3] [9],  \level_6_sums[13][3] [5:0] }), .in_2({1'b0, 1'b0, 
    1'b0, \level_6_sums[13][2] [9],  \level_6_sums[13][2] [5:0] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    n_2996_danc, n_2976_danc, \dot_product_and_ReLU[0].product_terms[27][0] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[125][1] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[123][1] }), .in_6({1'b0, 
    1'b0, 1'b0, 1'b0, n_3001_danc, n_2926_danc}), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_2927_danc, n_2928_danc}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[75][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] }), .in_12({1'b0, 1'b0, 1'b0, 
    1'b0, n_2870_danc, n_2871_danc}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] , 1'b0}), .in_15({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[48][1] , 
    1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] }), .in_18({
    1'b0, 1'b0, 1'b0, 1'b0, n_1413, n_2823_danc}), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[28][0] , 1'b0}), .in_20({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[22][0] }),
     .in_21({1'b0, 1'b0, 1'b0, 1'b0, n_1467, n_1466}), .in_22({1'b0, 1'b0, 1'b0, 
    1'b0, n_1431, n_1430}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, n_1481, n_1480}),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] }), .in_25({1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] }), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }), .in_27({
    1'b0, \dot_product_and_ReLU[0].product_terms[119][0] }), .in_28({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }), .in_29({
    1'b0, \dot_product_and_ReLU[17].product_terms[112][2] }), .in_30({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[113][1] }),
     .in_31({1'b0, \dot_product_and_ReLU[1].product_terms[108][0] }), .in_32({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[109][1] }),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[16].product_terms[107][0] }), .in_35({1'b0, 
    \dot_product_and_ReLU[16].product_terms[102][2] }), .in_36({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[103][0] , 1'b0}), .in_37({
    1'b0, \dot_product_and_ReLU[4].product_terms[101][1] }), .in_38(
    \dot_product_and_ReLU[4].product_terms[98][1] ), .in_39({
    \dot_product_and_ReLU[14].product_terms[99][0] , 1'b0}), .in_40({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[97][0] }), .in_41({
    \dot_product_and_ReLU[8].product_terms[92][1] , 1'b0}), .in_42({
    \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_43({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[90][0] , 1'b0}), .in_44({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_45(
    \dot_product_and_ReLU[0].product_terms[88][1] ), .in_46(
    \dot_product_and_ReLU[13].product_terms[89][0] ), .in_47({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[12].product_terms[87][0] , 1'b0}), .in_48({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}), .in_49({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[85][0] , 1'b0}),
     .in_50({1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_51(
    \dot_product_and_ReLU[3].product_terms[83][0] ), .in_52({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }), .in_53({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[79][0] , 1'b0}), .in_54({1'b0, 
    \dot_product_and_ReLU[1].product_terms[77][0] }), .in_55({1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[72][0] }), .in_56({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }), .in_57({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[67][0] , 1'b0}), .in_58(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .in_59(
    \dot_product_and_ReLU[0].product_terms[65][0] ), .in_60(
    \dot_product_and_ReLU[1].product_terms[62][0] ), .in_61({1'b0, 
    \dot_product_and_ReLU[0].product_terms[63][1] }), .in_62({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[60][2] }), .in_63({1'b0, 
    \dot_product_and_ReLU[15].product_terms[61][1] }), .in_64({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[59][1] , 1'b0}), .in_65({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[56][1] }),
     .in_66({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] }), .in_67(
    \dot_product_and_ReLU[11].product_terms[50][0] ), .in_68({1'b0, 
    \dot_product_and_ReLU[5].product_terms[51][1] }), .in_69({1'b0, 
    \dot_product_and_ReLU[0].product_terms[41][0] }), .in_70({1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[36][0] , 1'b0, 1'b0}), .in_71({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_72({
    1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }), .in_73(
    \dot_product_and_ReLU[2].product_terms[33][0] ), .in_74(
    \dot_product_and_ReLU[1].product_terms[30][1] ), .in_75(
    \dot_product_and_ReLU[2].product_terms[31][1] ), .in_76({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[20][0] , 1'b0}), .in_77({1'b0, 
    \dot_product_and_ReLU[2].product_terms[21][1] }), .in_78({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[16][0] , 1'b0}), .in_79({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[17][1] , 1'b0}), .in_80({1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] }), .in_81({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_82({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[11][1] }), .in_83({
    1'b0, \dot_product_and_ReLU[2].product_terms[4][0] , 1'b0, 1'b0}), .in_84({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}),
     .in_85({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_86({1'b0, 
    \dot_product_and_ReLU[4].product_terms[3][0] }), .in_87({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({
    \level_8_sums[13][8] , UNCONNECTED44, \level_8_sums[13][7] , 
    \level_8_sums[13][6] , \level_8_sums[13][5] , \final_sums[13][4] , 
    \final_sums[13][3] , \final_sums[13][2] , \final_sums[13][1] , 
    \final_sums[13][0] }));
  WALLACE_CSA_DUMMY_OP106_group_109836_6302 WALLACE_CSA_DUMMY_OP106_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[210]}), .in_1({1'b0, B[211], 1'b0}), .in_2({1'b0, 
    1'b0, 1'b0, B[237], 1'b0}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, B[233]}), .in_4({
    1'b0, 1'b0, 1'b0, 1'b0, B[217]}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, B[203]}),
     .in_6({1'b0, 1'b0, 1'b0, \level_6_sums[6][2] [9],  \level_6_sums[6][2] [5:0] }), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[251], B[250]}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[244]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_1488, n_1553}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[234]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1522, 
    n_1521}), .in_12({1'b0, 1'b0, 1'b0, n_1487, n_2602_danc, n_2603_danc}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[218]}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, B[213], 1'b0}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, B[198], 1'b0}),
     .in_16({1'b0, 1'b0, 1'b0, n_1486, n_1539, 1'b0}), .in_17({1'b0, 1'b0, 1'b0, 
    1'b0, B[254]}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, B[255]}), .in_19({1'b0, 
    1'b0, 1'b0, B[252], 1'b0}), .in_20({1'b0, B[253], 1'b0}), .in_21({1'b0, 
    1'b0, B[246]}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, B[247]}), .in_23(B[240]),
     .in_24(B[241]), .in_25({1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_26({1'b0, 
    1'b0, 1'b0, B[239], 1'b0}), .in_27({1'b0, B[230]}), .in_28({1'b0, 1'b0, 
    1'b0, 1'b0, B[231]}), .in_29({1'b0, 1'b0, 1'b0, 1'b0, B[228]}), .in_30({
    1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_31({1'b0, B[225]}), .in_32({1'b0, 
    B[220]}), .in_33({1'b0, 1'b0, 1'b0, B[221], 1'b0}), .in_34({1'b0, 1'b0, 
    1'b0, B[215], 1'b0}), .in_35(B[208]), .in_36(B[209]), .in_37(B[206]),
     .in_38({B[207], 1'b0}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[204]}), .in_40({
    1'b0, 1'b0, 1'b0, B[205], 1'b0}), .in_41({1'b0, B[200]}), .in_42({1'b0, 
    1'b0, 1'b0, 1'b0, B[201]}), .in_43({1'b0, 1'b0, 1'b0, 1'b0, B[194]}),
     .in_44({1'b0, B[195]}), .in_45({1'b0, 1'b0, 1'b0, 1'b0, B[193]}), .out_0({
    \level_7_sums[6][1] [9], UNCONNECTED46, UNCONNECTED45,  \level_7_sums[6][1] [6:0] }));
  WALLACE_CSA_DUMMY_OP106_group_109836 WALLACE_CSA_DUMMY_OP106_groupi4118(.in_0({
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }),
     .in_3({1'b0, \dot_product_and_ReLU[1].product_terms[19][1] , 1'b0}), .in_4({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[49][0] }),
     .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[29][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, n_2772_danc, n_2773_danc}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[63][1] , 
    \dot_product_and_ReLU[1].product_terms[62][0] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[60][2] , 1'b0}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}),
     .in_10({1'b0, 1'b0, 1'b0, n_2779_danc, n_2780_danc, 
    \dot_product_and_ReLU[2].product_terms[40][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[34][0] }), .in_13({
    1'b0, \dot_product_and_ReLU[2].product_terms[35][0] }), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[26][2] }),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[20][0] }), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, n_2787_danc, n_2788_danc}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    n_2980_danc, n_2981_danc}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] }), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, n_2793_danc, n_2794_danc}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0}), .in_21({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }), .in_22({1'b0, 
    \dot_product_and_ReLU[17].product_terms[53][1] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] }), .in_24({
    1'b0, \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] }), .in_26({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[45][1] , 1'b0}),
     .in_27({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_28({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[43][0] , 1'b0}), .in_29({
    \dot_product_and_ReLU[7].product_terms[38][1] , 1'b0}), .in_30({1'b0, 
    \dot_product_and_ReLU[0].product_terms[39][0] }), .in_31({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[31][1] }), .in_33({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] , 1'b0}), .in_34({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[25][0] }),
     .in_35({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] }), .in_36({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] , 1'b0}), .in_37({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[12][0] }), .in_38({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }),
     .in_39({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[6][2] }), .in_40({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }), .in_41({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] }), .out_0({
    \level_6_sums[5][0] [9], UNCONNECTED49, UNCONNECTED48, UNCONNECTED47,  \level_6_sums[5][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP109_group_109822_6312 WALLACE_CSA_DUMMY_OP109_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_1({1'b0, 1'b0, 1'b0, B[251], 1'b0}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, B[210]}), .in_3({1'b0, B[211], 1'b0}),
     .in_4({1'b0, 1'b0, 1'b0, B[194], 1'b0}), .in_5({1'b0, B[195], 1'b0}),
     .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_1517, n_1516}), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, B[255]}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, n_1496, n_1495}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, B[244], 1'b0}), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, B[240], 1'b0}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[235]}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, B[230], 1'b0}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[226]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, n_1214, n_1547}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, n_1514, n_1513}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, B[216], 1'b0}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[212]}),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0, B[206], 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[198]}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[192]}),
     .in_21({1'b0, 1'b0, 1'b0, 1'b0, B[248]}), .in_22({1'b0, B[249]}), .in_23({
    1'b0, 1'b0, 1'b0, 1'b0, B[242]}), .in_24({1'b0, B[243], 1'b0}), .in_25({
    1'b0, B[233]}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, B[222]}), .in_27({1'b0, 
    B[223]}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, B[218]}), .in_29({1'b0, 1'b0, 
    1'b0, 1'b0, B[219]}), .in_30({1'b0, 1'b0, 1'b0, B[214], 1'b0}), .in_31({
    1'b0, 1'b0, 1'b0, 1'b0, B[215]}), .in_32({1'b0, 1'b0, 1'b0, 1'b0, B[209]}),
     .in_33({1'b0, B[204]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[205]}), .in_35({
    1'b0, 1'b0, 1'b0, B[203], 1'b0}), .in_36({1'b0, 1'b0, 1'b0, 1'b0, B[200]}),
     .in_37({1'b0, B[201]}), .in_38({1'b0, B[197], 1'b0}), .out_0({
    \level_6_sums[3][3] [9], UNCONNECTED52, UNCONNECTED51, UNCONNECTED50,  \level_6_sums[3][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP109_group_109822 WALLACE_CSA_DUMMY_OP109_groupi4120(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }),
     .in_1({1'b0, \dot_product_and_ReLU[2].product_terms[33][0] , 1'b0}), .in_2({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0}),
     .in_3({\dot_product_and_ReLU[19].product_terms[46][2] , 1'b0}), .in_4({
    \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0}), .in_5({1'b0, 
    \level_7_sums[9][1] [9],  \level_7_sums[9][1] [7:0] }), .in_6({1'b0, 1'b0, 1'b0, 
    \level_3_sums[9][8] [7],  \level_3_sums[9][8] [3:0] }), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1427, n_1426, 
    1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[124][0] }), .in_10({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[120][1] , 
    \dot_product_and_ReLU[2].product_terms[121][1] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[116][0] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[106][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[98][1] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[88][1] }), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[82][0] }), .in_18({1'b0, 1'b0, 1'b0, 
    n_2862_danc, n_1436, 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[72][0] }), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[58][0] }),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] , 1'b0}), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] , 1'b0}),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_25({1'b0, 
    \dot_product_and_ReLU[6].product_terms[43][0] , 1'b0}), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[36][0] }), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[34][0] }), .in_28({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0, 1'b0}), .in_29({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[26][2] }),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[22][0] }), .in_31({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }), .in_32({1'b0, 
    1'b0, 1'b0, 1'b0, n_1442, n_2981_danc}), .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_34({1'b0, 1'b0, 
    1'b0, n_1470, n_1469, \dot_product_and_ReLU[2].product_terms[4][0] }),
     .in_35({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[0][0] , 
    1'b0, 1'b0}), .in_36({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_37({1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] }), .in_38({1'b0, 
    \dot_product_and_ReLU[3].product_terms[123][1] , 1'b0}), .in_39(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .in_40(
    \dot_product_and_ReLU[0].product_terms[119][0] ), .in_41({1'b0, 
    \dot_product_and_ReLU[2].product_terms[113][1] , 1'b0}), .in_42({1'b0, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_43(
    \dot_product_and_ReLU[16].product_terms[102][2] ), .in_44(
    \dot_product_and_ReLU[7].product_terms[103][0] ), .in_45({
    \dot_product_and_ReLU[0].product_terms[100][0] , 1'b0}), .in_46({
    \dot_product_and_ReLU[4].product_terms[101][1] , 1'b0}), .in_47({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[97][0] , 1'b0}), .in_48({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[94][1] , 1'b0}), .in_49({
    1'b0, \dot_product_and_ReLU[2].product_terms[95][0] }), .in_50({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_51({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_52({
    \dot_product_and_ReLU[3].product_terms[86][0] , 1'b0}), .in_53(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .in_54({1'b0, 
    \dot_product_and_ReLU[4].product_terms[79][0] }), .in_55({1'b0, 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_56({
    \dot_product_and_ReLU[1].product_terms[77][0] , 1'b0}), .in_57({1'b0, 
    \level_1_sums[4][37][1] }), .in_58(
    \dot_product_and_ReLU[5].product_terms[75][0] ), .in_59({
    \dot_product_and_ReLU[19].product_terms[60][2] , 1'b0}), .in_60(
    \dot_product_and_ReLU[15].product_terms[61][1] ), .in_61({
    \dot_product_and_ReLU[1].product_terms[56][1] , 1'b0}), .in_62({
    \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0}), .in_63({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[54][0] }), .in_64({1'b0, 
    \dot_product_and_ReLU[1].product_terms[55][0] }), .in_65({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[48][1] }), .in_66({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}), .in_67({
    1'b0, \dot_product_and_ReLU[3].product_terms[45][1] , 1'b0}), .in_68({
    \dot_product_and_ReLU[7].product_terms[38][1] , 1'b0}), .in_69({
    \dot_product_and_ReLU[0].product_terms[39][0] , 1'b0}), .in_70({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[29][0] , 1'b0}), .in_71({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] , 1'b0}),
     .in_72({1'b0, \dot_product_and_ReLU[1].product_terms[19][1] , 1'b0}),
     .in_73({\dot_product_and_ReLU[7].product_terms[16][0] , 1'b0}), .in_74({
    \dot_product_and_ReLU[0].product_terms[17][1] , 1'b0}), .in_75({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0}), .in_76({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }), .in_77({
    \dot_product_and_ReLU[19].product_terms[2][0] , 1'b0}), .in_78({1'b0, 
    \dot_product_and_ReLU[4].product_terms[3][0] }), .out_0({
    \level_8_sums[9][9] , \level_8_sums[9][8] , \level_8_sums[9][7] , 
    \level_8_sums[9][6] , \level_8_sums[9][5] , \level_8_sums[9][4] , 
    \level_8_sums[9][3] , \level_8_sums[9][2] , \level_8_sums[9][1] , 
    \final_sums[9][0] }));
  WALLACE_CSA_DUMMY_OP125_group_106193 WALLACE_CSA_DUMMY_OP125_groupi(.in_0({
    1'b0, \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, n_1478, n_1477, n_1476}), .in_3({1'b0, 1'b0, 1'b0, 
    1'b0, n_2772_danc, n_2773_danc}), .in_4(
    \dot_product_and_ReLU[11].product_terms[50][0] ), .in_5({
    \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }), .in_7({
    1'b0, 1'b0, 1'b0, n_1405, n_1414, 
    \dot_product_and_ReLU[2].product_terms[37][1] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[28][0] }),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, n_2975_danc, n_2976_danc}), .in_11({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[16][0] }), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[10][0] }), .in_14({1'b0, 
    1'b0, 1'b0, n_1462, n_1480, \dot_product_and_ReLU[7].product_terms[7][0] }),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_16({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[3][0] , 1'b0}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[56][1] }), .in_18({1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] }), .in_19({1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] }), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[53][1] }), .in_21({1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] , 1'b0}), .in_22({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0}), .in_23({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] , 1'b0}),
     .in_24({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[45][1] , 
    1'b0}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[42][1] }), .in_26({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[43][0] , 1'b0}), .in_27({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[41][0] , 1'b0}), .in_28({1'b0, 
    \dot_product_and_ReLU[2].product_terms[33][0] }), .in_29({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] }), .in_30({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[23][0] , 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[20][0] }), .in_32({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[18][0] }), .in_34({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }), .in_35({1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[14][1] , 1'b0, 1'b0}), .in_36({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[15][0] , 1'b0}),
     .in_37({1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[12][0] }),
     .in_38({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] , 
    1'b0}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] }), .in_40({1'b0, 
    \dot_product_and_ReLU[6].product_terms[9][0] , 1'b0}), .in_41({1'b0, 
    \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}), .out_0({
    \level_6_sums[16][0] [9], UNCONNECTED55, UNCONNECTED54, UNCONNECTED53,  \level_6_sums[16][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP127_group_109819 WALLACE_CSA_DUMMY_OP127_groupi(.in_0({
    1'b0, B[198], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[199]}), .in_2({1'b0, 
    1'b0, 1'b0, B[239], 1'b0}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_4({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[210]}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    B[244]}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0,  B[234:235] }), .in_8({1'b0, 1'b0, 1'b0, B[232], n_2861_danc, n_1549}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_1505, n_1521}), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, n_2667_danc, n_1547}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[217]}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_2864_danc, n_1434}), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[200]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[196]}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, n_1528, n_1527}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, B[192], 1'b0}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, B[252]}), .in_18({
    1'b0, 1'b0, 1'b0, B[253], 1'b0}), .in_19({B[250], 1'b0}), .in_20({B[251], 
    1'b0, 1'b0}), .in_21({1'b0, 1'b0, 1'b0, B[249], 1'b0}), .in_22({B[242], 
    1'b0}), .in_23(B[243]), .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[236]}), .in_25({
    1'b0, 1'b0, 1'b0, B[237], 1'b0}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, B[231]}),
     .in_27({1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_28({B[220], 1'b0}), .in_29({
    1'b0, B[221]}), .in_30({1'b0, 1'b0, 1'b0, B[218], 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, B[219]}), .in_32({1'b0, B[214]}), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, B[215]}), .in_34({1'b0, 1'b0, 1'b0, B[213], 1'b0}), .in_35({
    1'b0, 1'b0, 1'b0, 1'b0, B[206]}), .in_36({1'b0, 1'b0, B[207]}), .in_37({
    1'b0, 1'b0, 1'b0, B[205], 1'b0}), .out_0({\level_6_sums[12][3] [9], 
    UNCONNECTED58, UNCONNECTED57, UNCONNECTED56,  \level_6_sums[12][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP130_group_109827 WALLACE_CSA_DUMMY_OP130_groupi(.in_0({
    1'b0, B[234], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[235]}), .in_2({1'b0, 
    1'b0, 1'b0, B[194], 1'b0}), .in_3({1'b0, B[195], 1'b0}), .in_4({B[230], 
    1'b0}), .in_5(B[231]), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[254]}),
     .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_2631_danc, n_1495}), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[236]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[220]}),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, B[218], 1'b0}), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[209]}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[206]}),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, B[200], 1'b0}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, B[196], 1'b0}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[192]}),
     .in_16({B[252], 1'b0}), .in_17(B[253]), .in_18({1'b0, B[251], 1'b0}),
     .in_19({1'b0, B[249], 1'b0}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, B[244]}),
     .in_21({1'b0, 1'b0, 1'b0, B[245], 1'b0}), .in_22({1'b0, 1'b0, 1'b0, B[242], 
    1'b0}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, B[243]}), .in_24({1'b0, 1'b0, 1'b0, 
    B[241], 1'b0}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, B[239]}), .in_26({1'b0, 
    1'b0, 1'b0, B[233], 1'b0}), .in_27({1'b0, 1'b0, 1'b0, 1'b0, B[222]}),
     .in_28({1'b0, 1'b0, 1'b0, B[223], 1'b0}), .in_29({1'b0, 1'b0, 1'b0, B[216], 
    1'b0}), .in_30({1'b0, 1'b0, 1'b0, 1'b0, B[217]}), .in_31({B[214], 1'b0}),
     .in_32(B[215]), .in_33({1'b0, B[212]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, 
    B[213]}), .in_35({1'b0, B[211], 1'b0}), .in_36({1'b0, 1'b0, 1'b0, B[204], 
    1'b0}), .in_37({1'b0, 1'b0, 1'b0, 1'b0, B[205]}), .in_38({1'b0, 1'b0, 1'b0, 
    1'b0, B[202]}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[203]}), .in_40({1'b0, 
    1'b0, 1'b0, 1'b0, B[198]}), .in_41({1'b0, B[199]}), .out_0({
    \level_6_sums[16][3] [9], UNCONNECTED61, UNCONNECTED60, UNCONNECTED59,  \level_6_sums[16][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP131_group_106210 WALLACE_CSA_DUMMY_OP131_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }),
     .in_1({1'b0, \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0}), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[31][1] }),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[11][1] }), .in_4({1'b0, 1'b0, 
    \level_6_sums[17][1] [9],  \level_6_sums[17][1] [6:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1241, n_1240, 
    \dot_product_and_ReLU[0].product_terms[41][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, n_1213, n_1479}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1494, n_2773_danc}),
     .in_8({1'b0, 1'b0, 1'b0, n_1491, n_1490, n_1489}), .in_9({1'b0, 1'b0, 1'b0, 
    n_1405, n_1414, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_10({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[28][0] , 
    \dot_product_and_ReLU[0].product_terms[29][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }), .in_12({1'b0, 
    \dot_product_and_ReLU[14].product_terms[18][0] , 1'b0}), .in_13({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }), .in_14({
    \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}), .in_15({1'b0, 
    \dot_product_and_ReLU[0].product_terms[63][1] }), .in_16({1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[54][0] }), .in_18({1'b0, 
    \dot_product_and_ReLU[1].product_terms[55][0] , 1'b0, 1'b0}), .in_19({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] , 1'b0}), .in_20({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[53][1] , 1'b0}),
     .in_21({1'b0, \dot_product_and_ReLU[11].product_terms[50][0] }), .in_22({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}),
     .in_23(\dot_product_and_ReLU[19].product_terms[46][2] ), .in_24({1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[47][1] }), .in_25({1'b0, 
    \dot_product_and_ReLU[2].product_terms[44][1] }), .in_26({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[45][1] }), .in_27({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[35][0] }), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }), .in_29({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }),
     .in_30(\dot_product_and_ReLU[19].product_terms[26][2] ), .in_31({
    \dot_product_and_ReLU[0].product_terms[27][0] , 1'b0}), .in_32({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[24][0] , 1'b0}), .in_33({1'b0, 
    \dot_product_and_ReLU[3].product_terms[25][0] }), .in_34({
    \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_35(
    \dot_product_and_ReLU[0].product_terms[23][0] ), .in_36({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] , 1'b0}), .in_37({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[15][0] }), .in_38({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[12][0] }),
     .in_39({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[13][0] }), .in_40({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[9][0] , 1'b0}), .in_41({
    \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0}), .in_42({1'b0, 
    \dot_product_and_ReLU[7].product_terms[7][0] , 1'b0}), .in_43({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[4][0] }), .in_44({1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0, 1'b0}), .in_45({
    \dot_product_and_ReLU[19].product_terms[2][0] , 1'b0}), .in_46(
    \dot_product_and_ReLU[4].product_terms[3][0] ), .in_47({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[0][0] }), .in_48({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({
    \level_7_sums[17][0] [9], UNCONNECTED62,  \level_7_sums[17][0] [7:0] }));
  WALLACE_CSA_DUMMY_OP140_group_106218 WALLACE_CSA_DUMMY_OP140_groupi(.in_0({
    1'b0, \dot_product_and_ReLU[0].product_terms[22][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[41][0] }),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[123][1] }), .in_4({1'b0, 1'b0, 
    \level_7_sums[19][1] [9],  \level_7_sums[19][1] [6:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  \level_3_sums[19][14] [2:0] }), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, \level_3_sums[19][8] [7],  \level_3_sums[19][8] [2:0] }), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[120][1] , 1'b0}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[108][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[106][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[104] [1]}), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[102][2] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[100][0] , 1'b0}), .in_14({1'b0, 
    1'b0, 1'b0, 1'b0, n_1395, n_1394}), .in_15({1'b0, 1'b0, 1'b0, 
    \level_1_sums[3][46] [4], \level_1_sums[3][46] [0], 
    \dot_product_and_ReLU[8].product_terms[92][1] }), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[88][1] }), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[62][0] , 1'b0}),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }), .in_20({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[34][0] }), .in_21({1'b0, 1'b0, 1'b0, 
    1'b0, n_1484, n_1483}), .in_22({1'b0, 
    \dot_product_and_ReLU[1].product_terms[11][1] , 1'b0}), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] }), .in_24({
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[110][0] , 1'b0, 1'b0}),
     .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[111][0] }), .in_26({1'b0, 
    \dot_product_and_ReLU[0].product_terms[94][1] , 1'b0, 1'b0, 1'b0}), .in_27({
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[95][0] , 1'b0, 1'b0}),
     .in_28({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[90][0] }), .in_29({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[91][1] , 1'b0}), .in_30({1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] , 1'b0}), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[12].product_terms[87][0] }), .in_32({
    1'b0, \dot_product_and_ReLU[3].product_terms[84][0] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[85][0] }), .in_34({1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[82][0] , 1'b0, 1'b0}), .in_35({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}),
     .in_36({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[80][0] , 
    1'b0}), .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[81][0] }), .in_38({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }), .in_39({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[79][0] }), .in_40({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[76][0] }),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[77][0] }), .in_42({1'b0, 
    \level_1_sums[4][37][1] , 1'b0}), .in_43({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] }), .in_44({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[5].product_terms[72][0] }), .in_45({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }), .in_46({1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[60][2] , 1'b0, 1'b0}),
     .in_47({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[15].product_terms[61][1] , 
    1'b0}), .in_48({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[58][0] , 1'b0}), .in_49({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[59][1] , 1'b0}), .in_50({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[56][1] }),
     .in_51({1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0, 
    1'b0}), .in_52({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[48][1] , 1'b0}), .in_53({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}), .in_54({
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[46][2] , 1'b0, 1'b0}),
     .in_55({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[47][1] , 
    1'b0}), .in_56({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[44][1] }), .in_57({1'b0, 
    \dot_product_and_ReLU[3].product_terms[45][1] , 1'b0}), .in_58({1'b0, 
    \dot_product_and_ReLU[0].product_terms[39][0] , 1'b0, 1'b0}), .in_59({1'b0, 
    \dot_product_and_ReLU[8].product_terms[36][0] }), .in_60({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_61({1'b0, 
    \dot_product_and_ReLU[8].product_terms[32][1] }), .in_62({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }), .in_63({1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] }), .in_64({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[31][1] }), .in_65({1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[26][2] , 1'b0, 1'b0}), .in_66({
    1'b0, \dot_product_and_ReLU[0].product_terms[27][0] , 1'b0}), .in_67(
    \dot_product_and_ReLU[4].product_terms[24][0] ), .in_68({
    \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0}), .in_69({1'b0, 
    \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}), .in_70(
    \dot_product_and_ReLU[14].product_terms[18][0] ), .in_71(
    \dot_product_and_ReLU[1].product_terms[19][1] ), .in_72({1'b0, 
    \dot_product_and_ReLU[7].product_terms[16][0] }), .in_73({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[17][1] , 1'b0}), .in_74({1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] , 1'b0, 1'b0}), .in_75({1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] }), .in_76(
    \dot_product_and_ReLU[0].product_terms[13][0] ), .in_77({
    \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0, 1'b0}), .in_78({
    \dot_product_and_ReLU[7].product_terms[7][0] , 1'b0}), .in_79({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[4][0] }), .in_80({1'b0, 
    \dot_product_and_ReLU[0].product_terms[5][0] }), .in_81({1'b0, 
    \dot_product_and_ReLU[19].product_terms[2][0] }), .in_82(
    \dot_product_and_ReLU[4].product_terms[3][0] ), .in_83({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0, 1'b0}), .in_84({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({ \level_8_sums[19] [9:0] }));
  WALLACE_CSA_DUMMY_OP144_group_106215 WALLACE_CSA_DUMMY_OP144_groupi(.in_0({
    1'b0, \dot_product_and_ReLU[16].product_terms[12][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }),
     .in_3({1'b0, \dot_product_and_ReLU[1].product_terms[19][1] , 1'b0}), .in_4({
    1'b0, 1'b0, \level_7_sums[18][1] [9],  \level_7_sums[18][1] [6:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[18][4] [8],  \level_4_sums[18][4] [3:0] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  \level_3_sums[18][10] [2:0] }), .in_7({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[7][0] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[122][0] }), .in_9({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[123][1] , 1'b0}), .in_10({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[118][0] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[108][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[106][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[100][0] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, n_1395, n_1394}), .in_16({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[58][0] , 1'b0, 1'b0}), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, n_1216, n_1492}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] }), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[48][1] }), .in_20({
    1'b0, 1'b0, 1'b0, 1'b0, n_2817_danc, n_2818_danc}), .in_21({1'b0, 1'b0, 
    1'b0, n_2779_danc, n_2780_danc, 
    \dot_product_and_ReLU[2].product_terms[40][0] }), .in_22({1'b0, 1'b0, 1'b0, 
    1'b0, n_1475, n_1474}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[28][0] }), .in_24({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[22][0] }), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[14][1] , 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[10][0] , 1'b0}), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[9][0] }),
     .in_29({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[126][1] }),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[127][0] }), .in_31({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0}), .in_32({
    1'b0, \dot_product_and_ReLU[4].product_terms[125][1] , 1'b0}), .in_33({1'b0, 
    \dot_product_and_ReLU[2].product_terms[116][0] }), .in_34({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[117][0] , 1'b0}), .in_35({
    1'b0, \dot_product_and_ReLU[17].product_terms[112][2] }), .in_36(
    \dot_product_and_ReLU[2].product_terms[113][1] ), .in_37({1'b0, 
    \dot_product_and_ReLU[3].product_terms[110][0] }), .in_38(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .in_39({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[104] [1], 1'b0}), .in_40({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[105][0] , 1'b0}),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[103][0] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[98][1] }), .in_43({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] , 1'b0}),
     .in_44({1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[95][0] }),
     .in_45({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[92][1] , 
    1'b0}), .in_46({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_47({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[90][0] }), .in_48({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_49({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[88][1] , 1'b0}),
     .in_50({1'b0, 1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 1'b0, 
    1'b0}), .in_51(\dot_product_and_ReLU[1].product_terms[62][0] ), .in_52(
    \dot_product_and_ReLU[0].product_terms[63][1] ), .in_53(
    \dot_product_and_ReLU[19].product_terms[60][2] ), .in_54(
    \dot_product_and_ReLU[15].product_terms[61][1] ), .in_55({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[54][0] , 1'b0}), .in_56({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] }), .in_57({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[11].product_terms[50][0] , 1'b0}),
     .in_58({1'b0, \dot_product_and_ReLU[5].product_terms[51][1] }), .in_59({
    1'b0, \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0, 1'b0}), .in_60({
    \dot_product_and_ReLU[0].product_terms[42][1] , 1'b0}), .in_61({
    \dot_product_and_ReLU[6].product_terms[43][0] , 1'b0}), .in_62({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[36][0] , 1'b0}), .in_63({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_64({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }),
     .in_65({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[33][0] }), .in_66({1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0, 1'b0}), .in_67({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[31][1] , 1'b0}), .in_68({
    \dot_product_and_ReLU[4].product_terms[24][0] , 1'b0}), .in_69({1'b0, 
    \dot_product_and_ReLU[3].product_terms[25][0] }), .in_70({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }), .in_71({1'b0, 
    \dot_product_and_ReLU[0].product_terms[17][1] , 1'b0}), .in_72(
    \dot_product_and_ReLU[19].product_terms[2][0] ), .in_73(
    \dot_product_and_ReLU[4].product_terms[3][0] ), .in_74(
    \dot_product_and_ReLU[0].product_terms[0][0] ), .in_75({1'b0, 
    \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({
    \level_8_sums[18][8] , UNCONNECTED63, \level_8_sums[18][7] , 
    \level_8_sums[18][6] , \level_8_sums[18][5] , \level_8_sums[18][4] , 
    \level_8_sums[18][3] , \level_8_sums[18][2] , \level_8_sums[18][1] , 
    \final_sums[18][0] }));
  WALLACE_CSA_DUMMY_OP146_group_106214 WALLACE_CSA_DUMMY_OP146_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[27][0] }),
     .in_1({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[55][0] , 
    1'b0}), .in_2({1'b0, 1'b0, \level_7_sums[10][1] [9],  \level_7_sums[10][1] [6:0] }), .in_3({1'b0, 1'b0, 
    1'b0, \level_3_sums[10][12] [7],  \level_3_sums[10][12] [3:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0,  \level_2_sums[10][29] [2:0] }), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[70][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    n_1425, n_1424, n_1423}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_2925_danc, 
    n_2926_danc}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[112][2] , 1'b0}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[110][0] }),
     .in_10({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[106][0] , 
    1'b0}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[107][0] }), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, n_2927_danc, n_2928_danc}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[92][1] }), .in_14({1'b0, 
    \dot_product_and_ReLU[2].product_terms[91][1] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[86][0] }), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[80][0] }),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[76][0] }), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[65][0] }), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, n_1213, n_1479}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_21({1'b0, 1'b0, 
    1'b0, 1'b0, n_1491, n_1489}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[44][1] }), .in_24({
    1'b0, 1'b0, 1'b0, n_2822_danc, n_2823_danc, 
    \dot_product_and_ReLU[6].product_terms[43][0] }), .in_25({1'b0, 1'b0, 1'b0, 
    1'b0, n_2929_danc, n_2780_danc}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[32][1] , 
    \dot_product_and_ReLU[2].product_terms[33][0] }), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }), .in_28({1'b0, 
    1'b0, 1'b0, n_1473, n_1472, \dot_product_and_ReLU[1].product_terms[19][1] }),
     .in_29({1'b0, 1'b0, 1'b0, 1'b0, n_2787_danc, n_2788_danc}), .in_30({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[12][0] }),
     .in_31({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[10][0] }), .in_32({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[8][0] , 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, 1'b0, n_2793_danc, n_2794_danc}), .in_34(
    \dot_product_and_ReLU[4].product_terms[126][1] ), .in_35(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .in_36({
    \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0}), .in_37(
    \dot_product_and_ReLU[4].product_terms[125][1] ), .in_38({1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] }), .in_39({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }), .in_40({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[108][0] }),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[109][1] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] }), .in_43({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[85][0] , 1'b0}), .in_44({
    1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_45({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[83][0] }), .in_46({
    \dot_product_and_ReLU[10].product_terms[78][1] , 1'b0}), .in_47(
    \dot_product_and_ReLU[4].product_terms[79][0] ), .in_48({1'b0, 
    \dot_product_and_ReLU[5].product_terms[75][0] , 1'b0}), .in_49({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[72][0] }), .in_50({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] , 1'b0}), .in_51({
    1'b0, \dot_product_and_ReLU[0].product_terms[66][0] }), .in_52({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }), .in_53({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[63][1] , 1'b0}), .in_54({
    1'b0, \dot_product_and_ReLU[1].product_terms[56][1] }), .in_55({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[57][2] }), .in_56({
    \dot_product_and_ReLU[2].product_terms[52][0] , 1'b0}), .in_57({
    \dot_product_and_ReLU[17].product_terms[53][1] , 1'b0}), .in_58({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[38][1] , 1'b0}), .in_59({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] , 1'b0}), .in_60({
    1'b0, \dot_product_and_ReLU[2].product_terms[37][1] , 1'b0}), .in_61({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[35][0] , 1'b0}), .in_62({
    1'b0, \dot_product_and_ReLU[0].product_terms[28][0] }), .in_63({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[29][0] }), .in_64({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] }), .in_65({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0}),
     .in_66({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[23][0] }), .in_67({
    \dot_product_and_ReLU[4].product_terms[20][0] , 1'b0}), .in_68(
    \dot_product_and_ReLU[2].product_terms[21][1] ), .in_69({1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_70({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[6][2] }), .in_71({1'b0, 
    \dot_product_and_ReLU[7].product_terms[7][0] }), .in_72({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[4][0] , 1'b0}), .in_73({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] }), .in_74({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0}), .in_75({
    1'b0, \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({
    \level_8_sums[10] [8], UNCONNECTED64,  \level_8_sums[10] [7:0] }));
  WALLACE_CSA_DUMMY_OP149_group_109835 WALLACE_CSA_DUMMY_OP149_groupi(.in_0({
    1'b0, B[228], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_2({1'b0, 
    1'b0, 1'b0, B[238], 1'b0}), .in_3({1'b0, B[239], 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, B[218]}), .in_5({1'b0, B[219], 1'b0}), .in_6({1'b0, 1'b0, 
    \level_7_sums[4][0] [9],  \level_7_sums[4][0] [6:0] }), .in_7({1'b0, 1'b0, 1'b0, 
    \level_6_sums[4][2] [9],  \level_6_sums[4][2] [5:0] }), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[202]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, n_1535, n_1534}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, n_1533, n_1532}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1531, 
    n_1553}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_13({1'b0, 
    1'b0, 1'b0, n_1550, n_1549, B[232]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[230]}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[226]}), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, n_1548, n_1547}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, B[223], 
    1'b0}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[212]}), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, n_1530, n_1529}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, n_1528, 
    n_1527}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, B[192], 1'b0}), .in_22(B[252]),
     .in_23(B[253]), .in_24({1'b0, B[251]}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    B[248]}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, B[249]}), .in_27(B[246]), .in_28({
    1'b0, B[247]}), .in_29({1'b0, B[237]}), .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    B[234]}), .in_31({1'b0, B[235]}), .in_32({1'b0, B[220], 1'b0}), .in_33({
    1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_34({1'b0, 1'b0, B[217]}), .in_35({
    1'b0, 1'b0, 1'b0, 1'b0, B[214]}), .in_36({1'b0, 1'b0, 1'b0, 1'b0, B[215]}),
     .in_37({1'b0, B[208]}), .in_38({1'b0, 1'b0, 1'b0, 1'b0, B[209]}), .in_39({
    1'b0, B[207], 1'b0}), .in_40({1'b0, 1'b0, 1'b0, 1'b0, B[204]}), .in_41({
    1'b0, 1'b0, B[205]}), .in_42({1'b0, B[199], 1'b0}), .in_43({1'b0, 1'b0, 
    1'b0, B[196], 1'b0}), .in_44({1'b0, 1'b0, 1'b0, 1'b0, B[197]}), .out_0({
    \final_sums[4] [9], UNCONNECTED65,  \final_sums[4] [7:0] }));
  WALLACE_CSA_DUMMY_OP150_group_109838_6295 WALLACE_CSA_DUMMY_OP150_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[205]}), .in_1({1'b0, 1'b0, 1'b0, 
    \level_6_sums[5][1] [9],  \level_6_sums[5][1] [5:0] }), .in_2({1'b0, 1'b0, 1'b0, 
    \level_6_sums[5][0] [9],  \level_6_sums[5][0] [5:0] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[5][2] [9],  \level_6_sums[5][2] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[252]}),
     .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1526, n_1525}), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[248]}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[246]}), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    n_1524, n_1523}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[228]}), .in_11({
    1'b0, 1'b0, 1'b0, 1'b0, n_1522, n_1521}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    n_1214, n_1547}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, B[219], 1'b0}), .in_14({
    1'b0, 1'b0, 1'b0, B[212], 1'b0, 1'b0}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    B[210], 1'b0}), .in_16({1'b0, 1'b0, 1'b0, n_1520, n_1519, B[208]}), .in_17({
    1'b0, 1'b0, 1'b0, 1'b0, B[206], 1'b0}), .in_18({1'b0, 1'b0, 1'b0, 1'b0,  B[202:203] }),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[198]}), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, B[254]}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, B[255]}), .in_22({1'b0, 
    B[244]}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, B[245]}), .in_24({1'b0, 1'b0, 
    1'b0, B[242], 1'b0}), .in_25({1'b0, 1'b0, 1'b0, B[243], 1'b0}), .in_26({
    1'b0, 1'b0, 1'b0, 1'b0, B[240]}), .in_27({1'b0, 1'b0, 1'b0, B[241], 1'b0}),
     .in_28({1'b0, 1'b0, 1'b0, B[236], 1'b0}), .in_29({1'b0, 1'b0, 1'b0, 1'b0, 
    B[237]}), .in_30({1'b0, B[234], 1'b0}), .in_31({1'b0, 1'b0, 1'b0, B[235], 
    1'b0}), .in_32(B[232]), .in_33({1'b0, B[233]}), .in_34({1'b0, B[222]}),
     .in_35({1'b0, 1'b0, 1'b0, B[223], 1'b0}), .in_36({1'b0, 1'b0, 1'b0, B[221], 
    1'b0}), .in_37({1'b0, 1'b0, 1'b0, B[216], 1'b0}), .in_38({1'b0, B[217]}),
     .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[214]}), .in_40({1'b0, B[215]}), .in_41(
    B[200]), .in_42(B[201]), .in_43({1'b0, B[196]}), .in_44(B[197]), .in_45({
    1'b0, 1'b0, B[192], 1'b0, 1'b0}), .in_46({1'b0, B[193]}), .out_0({
    \final_sums[5] [9], UNCONNECTED66,  \final_sums[5] [7:0] }));
  WALLACE_CSA_DUMMY_OP150_group_109838 WALLACE_CSA_DUMMY_OP150_groupi4117(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[41][0] }),
     .in_1({1'b0, \dot_product_and_ReLU[0].product_terms[28][0] , 1'b0}), .in_2({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[29][0] , 1'b0}),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[58][0] }), .in_4({1'b0, 1'b0, 1'b0, 
    n_1216, n_1468, n_1492}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[11].product_terms[50][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, n_1491, n_1489}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1475, n_1474}),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[31][1] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[26][2] , 1'b0}), .in_10({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[20][0] , 
    1'b0}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[18][0] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, n_2980_danc, n_2981_danc}), .in_14({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[2][0] }),
     .in_15({1'b0, \dot_product_and_ReLU[15].product_terms[61][1] }), .in_16({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[54][0] }),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[55][0] }), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[52][0] }), .in_19({1'b0, 
    \dot_product_and_ReLU[17].product_terms[53][1] , 1'b0}), .in_20({1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_21({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0}), .in_22(
    \dot_product_and_ReLU[2].product_terms[44][1] ), .in_23({
    \dot_product_and_ReLU[3].product_terms[45][1] , 1'b0}), .in_24({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[43][0] }), .in_25({1'b0, 
    \dot_product_and_ReLU[7].product_terms[38][1] }), .in_26({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[39][0] , 1'b0}), .in_27({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[36][0] }), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_29({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] , 1'b0}),
     .in_30({1'b0, \dot_product_and_ReLU[3].product_terms[25][0] }), .in_31({
    \dot_product_and_ReLU[6].product_terms[14][1] , 1'b0}), .in_32({1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_33({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] , 1'b0}), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[9][0] , 1'b0}), .in_36({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[6][2] }), .in_37({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }),
     .in_38({1'b0, \dot_product_and_ReLU[2].product_terms[4][0] }), .in_39({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[5][0] , 1'b0}),
     .in_40({1'b0, \dot_product_and_ReLU[4].product_terms[1][0] }), .out_0({
    \level_6_sums[3][0] [9], UNCONNECTED69, UNCONNECTED68, UNCONNECTED67,  \level_6_sums[3][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP154_group_109832 WALLACE_CSA_DUMMY_OP154_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[207]}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[241]}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, B[228]}), .in_3({1'b0, B[229], 1'b0}),
     .in_4({1'b0, 1'b0, 1'b0, B[239], 1'b0}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, n_1429, n_1428}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[254]}),
     .in_7({1'b0, 1'b0, 1'b0, 1'b0, n_1526, n_1525}), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0,  B[244:245] }), .in_9({1'b0, 1'b0, 1'b0, 1'b0, B[242], 1'b0}), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, B[235]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, B[226], 1'b0}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[220]}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[215]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, B[213], 1'b0}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, B[208], 1'b0}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, n_2864_danc, n_1434}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[201]}),
     .in_18({1'b0, 1'b0, 1'b0, B[252], 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    B[253]}), .in_20({1'b0, B[248]}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, B[249]}),
     .in_22({1'b0, B[246], 1'b0}), .in_23({1'b0, 1'b0, 1'b0, B[247], 1'b0}),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[236]}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    B[237]}), .in_26({1'b0, 1'b0, B[233]}), .in_27({B[230], 1'b0}), .in_28({
    1'b0, B[231]}), .in_29({1'b0, B[224], 1'b0}), .in_30({1'b0, 1'b0, 1'b0, 
    1'b0, B[225]}), .in_31({1'b0, 1'b0, 1'b0, 1'b0, B[222]}), .in_32({1'b0, 
    1'b0, 1'b0, 1'b0, B[223]}), .in_33({1'b0, 1'b0, 1'b0, 1'b0, B[216]}),
     .in_34({1'b0, 1'b0, B[217]}), .in_35({1'b0, B[210], 1'b0}), .in_36({1'b0, 
    1'b0, 1'b0, 1'b0, B[211]}), .in_37(B[204]), .in_38({1'b0, B[205]}), .in_39(
    B[194]), .in_40({B[195], 1'b0}), .in_41({1'b0, 1'b0, B[192]}), .in_42({1'b0, 
    1'b0, 1'b0, B[193], 1'b0}), .out_0({\level_6_sums[13][3] [9], 
    UNCONNECTED72, UNCONNECTED71, UNCONNECTED70,  \level_6_sums[13][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP155_group_106213 WALLACE_CSA_DUMMY_OP155_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[32][1] }), .in_2({1'b0, 
    \dot_product_and_ReLU[2].product_terms[33][0] , 1'b0}), .in_3({1'b0, 1'b0, 
    \level_7_sums[6][1] [9],  \level_7_sums[6][1] [6:0] }), .in_4({1'b0, 1'b0, 1'b0, 
    \level_5_sums[6][3] [9],  \level_5_sums[6][3] [5:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[94][1] }), .in_6({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[90][0] , 1'b0}), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[75][0] }),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[63][1] , 1'b0}), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, n_2772_danc, n_2773_danc}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    n_1493, n_1492}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_13({1'b0, 1'b0, 
    1'b0, n_1490, n_1491, n_1489}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[37][1] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[28][0] }), .in_16({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[26][2] , 1'b0, 1'b0}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[23][0] , 1'b0}), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }), .in_19({
    1'b0, 1'b0, 1'b0, 1'b0, n_2787_danc, n_2788_danc}), .in_20({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[2][0] }),
     .in_22(\dot_product_and_ReLU[8].product_terms[92][1] ), .in_23({
    \dot_product_and_ReLU[0].product_terms[93][0] , 1'b0}), .in_24({1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] }), .in_25({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[12].product_terms[87][0] , 1'b0}), .in_26({
    \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}), .in_27({1'b0, 
    \dot_product_and_ReLU[1].product_terms[85][0] }), .in_28({
    \dot_product_and_ReLU[4].product_terms[82][0] , 1'b0}), .in_29(
    \dot_product_and_ReLU[3].product_terms[83][0] ), .in_30({1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[81][0] }), .in_31({1'b0, 
    \dot_product_and_ReLU[4].product_terms[79][0] , 1'b0, 1'b0}), .in_32(
    \dot_product_and_ReLU[0].product_terms[76][0] ), .in_33(
    \dot_product_and_ReLU[1].product_terms[77][0] ), .in_34({1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[71][0] }), .in_35({1'b0, 
    \dot_product_and_ReLU[1].product_terms[69][1] }), .in_36({1'b0, 
    \dot_product_and_ReLU[0].product_terms[66][0] }), .in_37(
    \dot_product_and_ReLU[2].product_terms[67][0] ), .in_38(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .in_39({1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] }), .in_40({1'b0, 
    \dot_product_and_ReLU[19].product_terms[60][2] }), .in_41(
    \dot_product_and_ReLU[15].product_terms[61][1] ), .in_42(
    \dot_product_and_ReLU[2].product_terms[52][0] ), .in_43(
    \dot_product_and_ReLU[17].product_terms[53][1] ), .in_44({1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] }), .in_45({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[47][1] }), .in_46({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[45][1] }), .in_47({
    1'b0, \dot_product_and_ReLU[6].product_terms[43][0] }), .in_48({1'b0, 
    \dot_product_and_ReLU[2].product_terms[40][0] }), .in_49({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[41][0] }), .in_50(
    \dot_product_and_ReLU[2].product_terms[34][0] ), .in_51(
    \dot_product_and_ReLU[2].product_terms[35][0] ), .in_52({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[30][1] }), .in_53({1'b0, 
    \dot_product_and_ReLU[2].product_terms[31][1] }), .in_54({1'b0, 
    \dot_product_and_ReLU[4].product_terms[24][0] }), .in_55({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0}), .in_56({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[14][1] , 1'b0}), .in_57({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[15][0] , 1'b0}), .in_58({
    1'b0, \dot_product_and_ReLU[16].product_terms[12][0] , 1'b0}), .in_59({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] , 1'b0}), .in_60({
    1'b0, \dot_product_and_ReLU[7].product_terms[10][0] }), .in_61({1'b0, 
    \dot_product_and_ReLU[1].product_terms[11][1] }), .in_62({1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] }), .in_63(
    \dot_product_and_ReLU[6].product_terms[9][0] ), .in_64({
    \dot_product_and_ReLU[0].product_terms[0][0] , 1'b0}), .in_65(
    \dot_product_and_ReLU[4].product_terms[1][0] ), .out_0({ \level_8_sums[6] [9:0] }));
  WALLACE_CSA_DUMMY_OP157_group_109824 WALLACE_CSA_DUMMY_OP157_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[245]}),
     .in_2({1'b0, 1'b0, 1'b0, 1'b0, B[195]}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    n_1506, n_1534}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[252]}), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0,  B[250:251] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[248]}),
     .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[246]}), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0,  B[240:241] }), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, B[237], 1'b0}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[234]}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1515, n_1549}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[210]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[209]}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[206]}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, B[202], 1'b0}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[200]}),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[196]}), .in_19({1'b0, B[242], 1'b0}),
     .in_20({1'b0, 1'b0, 1'b0, B[243], 1'b0}), .in_21({1'b0, B[227], 1'b0}),
     .in_22({1'b0, 1'b0, B[225]}), .in_23({1'b0, 1'b0, 1'b0, B[222], 1'b0}),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_25({1'b0, 1'b0, 1'b0, B[220], 
    1'b0}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, B[218]}), .in_28({1'b0, B[219]}), .in_29(B[216]), .in_30(B[217]),
     .in_31({1'b0, B[214], 1'b0}), .in_32({1'b0, 1'b0, 1'b0, 1'b0, B[215]}),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, B[212]}), .in_34({1'b0, 1'b0, 1'b0, B[213], 
    1'b0}), .in_35({1'b0, 1'b0, 1'b0, 1'b0, B[204]}), .in_36({1'b0, 1'b0, 1'b0, 
    1'b0, B[205]}), .in_37({1'b0, 1'b0, 1'b0, B[198], 1'b0}), .in_38({1'b0, 
    1'b0, 1'b0, 1'b0, B[199]}), .in_39(B[192]), .in_40(B[193]), .out_0({
    \level_6_sums[15][3] [9], UNCONNECTED75, UNCONNECTED74, UNCONNECTED73,  \level_6_sums[15][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP162_group_109829_6307 WALLACE_CSA_DUMMY_OP162_groupi(.in_0({
    1'b0, B[234], 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[235]}), .in_2({1'b0, 
    1'b0, 1'b0, B[210], 1'b0}), .in_3({1'b0, B[211], 1'b0}), .in_4({1'b0, 
    B[198], 1'b0}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, B[199]}), .in_6({1'b0, 1'b0, 
    1'b0, \level_6_sums[19][2] [9],  \level_6_sums[19][2] [5:0] }), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[242], 1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[254]}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[250]}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[248]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[246]}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, B[244], 1'b0}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[238]}), .in_14({1'b0, 1'b0, 1'b0, B[232], n_2861_danc, n_1549}), .in_15({
    1'b0, 1'b0, 1'b0, 1'b0, B[224], 1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, B[222]}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_18({
    1'b0, 1'b0, 1'b0, n_1546, n_1545, B[218]}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, B[217]}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[208]}), .in_21({
    1'b0, 1'b0, 1'b0, 1'b0, B[202], 1'b0}), .in_22({1'b0, B[252]}), .in_23({
    1'b0, 1'b0, 1'b0, B[253], 1'b0}), .in_24(B[236]), .in_25(B[237]), .in_26({
    1'b0, B[231], 1'b0}), .in_27({1'b0, 1'b0, 1'b0, B[229], 1'b0}), .in_28({
    1'b0, 1'b0, B[227]}), .in_29({1'b0, 1'b0, 1'b0, B[214], 1'b0}), .in_30({
    1'b0, 1'b0, B[215]}), .in_31(B[212]), .in_32(B[213]), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, B[206]}), .in_34({1'b0, B[207], 1'b0}), .in_35(B[204]), .in_36({
    B[205], 1'b0}), .in_37({1'b0, 1'b0, B[201], 1'b0, 1'b0}), .in_38({1'b0, 
    1'b0, 1'b0, 1'b0, B[197]}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[195]}),
     .in_40({B[192], 1'b0}), .in_41(B[193]), .out_0({\level_7_sums[19][1] [9], 
    UNCONNECTED77, UNCONNECTED76,  \level_7_sums[19][1] [6:0] }));
  WALLACE_CSA_DUMMY_OP162_group_109829 WALLACE_CSA_DUMMY_OP162_groupi4119(.in_0({
    1'b0, \dot_product_and_ReLU[16].product_terms[12][0] , 1'b0}), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[13][0] }), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[62][0] }),
     .in_3({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[63][1] , 
    1'b0}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, n_2817_danc, n_2818_danc}), .in_6({1'b0, 1'b0, 1'b0, n_2822_danc, 
    n_2823_danc, \dot_product_and_ReLU[6].product_terms[43][0] }), .in_7({1'b0, 
    1'b0, 1'b0, n_2779_danc, n_2780_danc, 
    \dot_product_and_ReLU[2].product_terms[40][0] }), .in_8({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[38][1] , 1'b0}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }), .in_10({1'b0, 
    \dot_product_and_ReLU[2].product_terms[35][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[26][2] }), .in_12({
    1'b0, 1'b0, 1'b0, 1'b0, n_2826_danc, n_1443}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[14].product_terms[18][0] , 1'b0}), .in_14({
    1'b0, 1'b0, 1'b0, 1'b0, n_1442, n_2981_danc}), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[4][0] , 1'b0}), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, n_1461, n_2757_danc}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[58][0] }), .in_18({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[59][1] , 1'b0}), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[56][1] }), .in_20({
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0, 1'b0}),
     .in_21({1'b0, \dot_product_and_ReLU[1].product_terms[55][0] }), .in_22({
    1'b0, \dot_product_and_ReLU[11].product_terms[50][0] , 1'b0}), .in_23({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[51][1] }), .in_24({
    1'b0, \dot_product_and_ReLU[19].product_terms[48][1] }), .in_25({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[49][0] , 1'b0}), .in_26({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[46][2] }),
     .in_27({1'b0, \dot_product_and_ReLU[3].product_terms[47][1] }), .in_28({
    1'b0, \dot_product_and_ReLU[2].product_terms[31][1] , 1'b0}), .in_29({1'b0, 
    \dot_product_and_ReLU[0].product_terms[28][0] }), .in_30({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[29][0] }), .in_31(
    \dot_product_and_ReLU[4].product_terms[24][0] ), .in_32({
    \dot_product_and_ReLU[3].product_terms[25][0] , 1'b0, 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] , 1'b0}), .in_34(
    \dot_product_and_ReLU[7].product_terms[16][0] ), .in_35(
    \dot_product_and_ReLU[0].product_terms[17][1] ), .in_36({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[14][1] }), .in_37({1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] , 1'b0}), .in_38({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[8][0] , 1'b0}), .in_39({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[9][0] }), .in_40({
    \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0}), .in_41(
    \dot_product_and_ReLU[7].product_terms[7][0] ), .out_0({
    \level_6_sums[7][0] [9], UNCONNECTED80, UNCONNECTED79, UNCONNECTED78,  \level_6_sums[7][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP258_group_359288 WALLACE_CSA_DUMMY_OP258_groupi(.in_0({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 1'b0}),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[185][0] }), .in_2({
    \level_1_sums[1][81][0] , 1'b0}), .in_3({1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] }), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[191][1] , 1'b0}), .in_5({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] , 
    \dot_product_and_ReLU[0].product_terms[189][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[178][0] }), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, n_1454, \level_1_sums[16][87] [1]}), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[172][1] , 1'b0}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[140] [0]}), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] }),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, n_1441, n_1440}), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[18].product_terms[186][0] }), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[187][0] }),
     .in_18({1'b0, \dot_product_and_ReLU[8].product_terms[182][0] }), .in_19(
    \dot_product_and_ReLU[18].product_terms[183][1] ), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[180][0] }), .in_21({1'b0, 
    \dot_product_and_ReLU[3].product_terms[181][0] }), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[177][0] }), .in_23({
    1'b0, \dot_product_and_ReLU[1].product_terms[170][0] }), .in_24({1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[171][1] , 1'b0, 1'b0}), .in_25({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[168][0] , 1'b0}),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[169][0] }), .in_27(
    \dot_product_and_ReLU[3].product_terms[164][0] ), .in_28({
    \dot_product_and_ReLU[2].product_terms[165][0] , 1'b0}), .in_29({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[158][0] , 1'b0}), .in_30({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[159][1] }),
     .in_31({1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[156][2] , 1'b0, 
    1'b0}), .in_32({1'b0, \dot_product_and_ReLU[0].product_terms[157][0] }),
     .in_33({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[152][0] , 
    1'b0}), .in_34({1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }),
     .in_35(\dot_product_and_ReLU[0].product_terms[150][0] ), .in_36({
    \dot_product_and_ReLU[3].product_terms[151][0] , 1'b0}), .in_37({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[148][0] }), .in_38({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[149][0] }),
     .in_39({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 
    1'b0}), .in_40({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[142][0] }), .in_41({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[143][0] , 1'b0}), .in_42({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[136][1] }),
     .in_43({1'b0, \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}),
     .in_44({1'b0, \dot_product_and_ReLU[1].product_terms[132][1] , 1'b0}),
     .in_45({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[133][0] , 
    1'b0}), .in_46({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[128][1] , 1'b0}), .in_47({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[129][0] }),
     .out_0({\level_6_sums[17][2] [9], UNCONNECTED83, UNCONNECTED82, 
    UNCONNECTED81,  \level_6_sums[17][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP752_group_359251 WALLACE_CSA_DUMMY_OP752_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[156][2] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[157][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[159][1] }), .in_3({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 1'b0}), .in_4({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}), .in_5({
    1'b0, \dot_product_and_ReLU[4].product_terms[166][0] , 1'b0}), .in_6({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[167][0] , 1'b0}), .in_7({
    1'b0, 1'b0, 1'b0, 1'b0, n_1403, n_1402, n_1401}), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, n_1212, n_1536}), .in_10({1'b0, 1'b0, 1'b0, n_1400, 
    n_1399, \dot_product_and_ReLU[1].product_terms[176][0] }), .in_11({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1398, n_1452}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[165][0] }), .in_14({
    1'b0, 1'b0, 1'b0,  \level_1_sums[2][73] [2:0] }), .in_15({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[144][0] , 1'b0, 1'b0}), .in_16({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[130][0] , 
    1'b0}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, n_1397, n_1396}), .in_18({1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[191][1] }), .in_20(
    \dot_product_and_ReLU[6].product_terms[188][1] ), .in_21({
    \dot_product_and_ReLU[0].product_terms[189][0] , 1'b0}), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[184][1] }), .in_23({
    1'b0, \dot_product_and_ReLU[5].product_terms[185][0] }), .in_24({
    \dot_product_and_ReLU[8].product_terms[182][0] , 1'b0}), .in_25(
    \dot_product_and_ReLU[18].product_terms[183][1] ), .in_26({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] , 1'b0}), .in_27({1'b0, 
    \dot_product_and_ReLU[3].product_terms[181][0] , 1'b0}), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[174][1] }),
     .in_29({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[175][0] }), .in_30({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[169][0] }), .in_31({1'b0, 1'b0, 
    1'b0, \level_1_sums[1][81][0] , 1'b0}), .in_32({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] }), .in_33({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}), .in_34({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] }),
     .in_35({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_36({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_37({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[152][0] }),
     .in_38({1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }), .in_39({
    1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }), .in_40({1'b0, 
    \dot_product_and_ReLU[1].product_terms[149][0] , 1'b0}), .in_41({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[142][0] , 1'b0}),
     .in_42({1'b0, \dot_product_and_ReLU[2].product_terms[143][0] }), .in_43({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0]}),
     .in_44({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[141][0] , 
    1'b0}), .out_0({\level_6_sums[5][2] [9], UNCONNECTED86, UNCONNECTED85, 
    UNCONNECTED84,  \level_6_sums[5][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP754_group_359252 WALLACE_CSA_DUMMY_OP754_groupi(.in_0({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[164][0] , 1'b0}),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[165][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, n_1403, n_1402, n_1401}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_5({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[185][0] , 1'b0}),
     .in_6({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] , 
    \dot_product_and_ReLU[3].product_terms[181][0] }), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[179][0] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] , 
    \dot_product_and_ReLU[10].product_terms[172][1] }), .in_9({1'b0, 1'b0, 
    1'b0, n_1386, n_1385, n_1384}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] , \level_1_sums[1][81][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, n_1393, n_1392}), .in_12({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_13({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] , 
    \dot_product_and_ReLU[9].product_terms[152][0] }), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, n_1383, n_1382}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] }), .in_16({1'b0, 
    \dot_product_and_ReLU[0].product_terms[189][0] , 1'b0}), .in_17({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[182][0] }),
     .in_18({1'b0, \dot_product_and_ReLU[18].product_terms[183][1] }), .in_19({
    \dot_product_and_ReLU[1].product_terms[176][0] , 1'b0}), .in_20({
    \dot_product_and_ReLU[0].product_terms[177][0] , 1'b0}), .in_21({
    \dot_product_and_ReLU[2].product_terms[174][1] , 1'b0}), .in_22({
    \dot_product_and_ReLU[2].product_terms[175][0] , 1'b0}), .in_23({
    \dot_product_and_ReLU[1].product_terms[170][0] , 1'b0, 1'b0}), .in_24(
    \dot_product_and_ReLU[1].product_terms[171][1] ), .in_25({1'b0, 
    \dot_product_and_ReLU[3].product_terms[168][0] }), .in_26(
    \dot_product_and_ReLU[0].product_terms[169][0] ), .in_27({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[5].product_terms[160][1] }), .in_28({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] }), .in_29({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[156][2] }),
     .in_30({1'b0, \dot_product_and_ReLU[0].product_terms[157][0] , 1'b0}),
     .in_31({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[150][0] , 
    1'b0}), .in_32({1'b0, \dot_product_and_ReLU[3].product_terms[151][0] , 
    1'b0}), .in_33({1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[146][0] }), .in_34({
    \dot_product_and_ReLU[1].product_terms[147][0] , 1'b0}), .in_35({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[145][1] }), .in_36({
    \dot_product_and_ReLU[0].product_terms[142][0] , 1'b0}), .in_37({
    \dot_product_and_ReLU[2].product_terms[143][0] , 1'b0}), .in_38({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 1'b0}), .in_39({
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[141][0] }), .in_40({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[138][0] }),
     .in_41({1'b0, \dot_product_and_ReLU[8].product_terms[139][0] }), .in_42({
    \dot_product_and_ReLU[4].product_terms[136][1] , 1'b0}), .in_43({
    \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}), .in_44({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[131][0] }), .in_45({
    1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }), .in_46({
    \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0, 1'b0}), .out_0({
    \level_6_sums[11][2] [9], UNCONNECTED88, UNCONNECTED87,  \level_6_sums[11][2] [6:0] }));
  WALLACE_CSA_DUMMY_OP758_group_359250 WALLACE_CSA_DUMMY_OP758_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[135][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }), .in_3({1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[129][0] }), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[141][0] }), .in_5({1'b0, 1'b0, 
    1'b0, 1'b0, n_1234, n_1233, n_1232}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[186][0] }), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[185][0] , 1'b0}), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[175][0] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0,  \level_1_sums[12][86] [1:0] }), .in_10({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[171][1] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1439, n_1448}), .in_13({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_14({
    1'b0, 1'b0, 1'b0, 1'b0, n_1383, n_1382}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, n_1409, n_1408}), .in_17({1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[191][1] }), .in_19({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] }),
     .in_20({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[189][0] }), .in_21({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[18].product_terms[183][1] , 1'b0}), .in_22({
    1'b0, \dot_product_and_ReLU[8].product_terms[180][0] }), .in_23({
    \dot_product_and_ReLU[3].product_terms[181][0] , 1'b0}), .in_24({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[166][0] }), .in_25({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[167][0] }),
     .in_26({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[165][0] }), .in_27({1'b0, 
    \level_1_sums[1][81][0] , 1'b0}), .in_28({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[163][0] , 1'b0}), .in_29(
    \dot_product_and_ReLU[1].product_terms[158][0] ), .in_30({
    \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0, 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[152][0] , 1'b0}),
     .in_32({1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[151][0] }), .in_34(
    \dot_product_and_ReLU[2].product_terms[144][0] ), .in_35(
    \dot_product_and_ReLU[0].product_terms[145][1] ), .in_36({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[19].product_terms[138][0] }), .in_37({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] }),
     .in_38({1'b0, \dot_product_and_ReLU[4].product_terms[136][1] }), .in_39({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[137][0] }),
     .in_40({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[132][1] }), .in_41({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[133][0] }), .in_42({
    1'b0, \dot_product_and_ReLU[0].product_terms[130][0] }), .in_43({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[131][0] }), .out_0({
    \level_6_sums[18][2] [9], UNCONNECTED91, UNCONNECTED90, UNCONNECTED89,  \level_6_sums[18][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP791_group_359281 WALLACE_CSA_DUMMY_OP791_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[186][0] }),
     .in_1({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 
    1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[137][0] }), .in_3({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[171][1] }), .in_5({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] , 1'b0}), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[191][1] , 
    1'b0}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[184][1] , 1'b0}), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[182][0] }), .in_9({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[179][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[176][0] , 1'b0}),
     .in_11({1'b0, 1'b0, 1'b0,  \level_1_sums[16][87] [2:1] , \dot_product_and_ReLU[2].product_terms[174][1] }),
     .in_12({1'b0, 1'b0, 1'b0, n_1386, n_1385, n_1384}), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[165][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[1][81][0] }), .in_15({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] , 
    \dot_product_and_ReLU[5].product_terms[160][1] }), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[150][0] , 1'b0}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[148][0] , 1'b0}), .in_18({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[144][0] }), .in_20({1'b0, 1'b0, 
    1'b0, n_1380, n_1379, \dot_product_and_ReLU[17].product_terms[140] [0]}),
     .in_21({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[128][1] , 1'b0}),
     .in_23(\dot_product_and_ReLU[8].product_terms[180][0] ), .in_24({
    \dot_product_and_ReLU[3].product_terms[181][0] , 1'b0}), .in_25({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[172][1] , 1'b0}), .in_26({
    1'b0, \dot_product_and_ReLU[8].product_terms[173][1] }), .in_27({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[168][0] }), .in_28({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[169][0] }),
     .in_29({1'b0, \dot_product_and_ReLU[1].product_terms[158][0] }), .in_30({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0}),
     .in_31(\dot_product_and_ReLU[17].product_terms[156][2] ), .in_32({
    \dot_product_and_ReLU[0].product_terms[157][0] , 1'b0}), .in_33({
    \dot_product_and_ReLU[9].product_terms[152][0] , 1'b0}), .in_34({
    \dot_product_and_ReLU[18].product_terms[153][0] , 1'b0}), .in_35({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[143][0] }),
     .in_36({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] , 
    1'b0}), .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[135][0] }), .in_38({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[130][0] , 1'b0}), .in_39({
    1'b0, \dot_product_and_ReLU[14].product_terms[131][0] , 1'b0}), .out_0({
    \level_6_sums[13][2] [9], UNCONNECTED94, UNCONNECTED93, UNCONNECTED92,  \level_6_sums[13][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP800_group_359276 WALLACE_CSA_DUMMY_OP800_groupi(.in_0({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] , 1'b0}),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[133][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[157][0] }), .in_3({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[143][0] }), .in_4({1'b0, 
    1'b0, 1'b0, \level_3_sums[19][22][4] , \level_3_sums[19][22][3] , 
    \level_3_sums[19][22][2] , \level_3_sums[19][22][1] , 
    \level_3_sums[19][22][0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] , 
    \dot_product_and_ReLU[0].product_terms[189][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[184][1] }),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[174][1] , 1'b0}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[170][0] }),
     .in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[168][0] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[165][0] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[1][81][0] }), .in_13({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[152][0] }), .in_14({1'b0, 
    \dot_product_and_ReLU[0].product_terms[150][0] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }), .in_16({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[136][1] , 
    1'b0}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] , 1'b0}), .in_18({1'b0, 
    1'b0, 1'b0, 1'b0, n_1441, n_1440}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[128][1] }), .in_20({
    \dot_product_and_ReLU[4].product_terms[190][1] , 1'b0}), .in_21({
    \dot_product_and_ReLU[0].product_terms[191][1] , 1'b0}), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] }), .in_23({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}),
     .in_24({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] , 
    1'b0}), .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[155][0] }), .in_27({
    1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }), .in_28({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[147][0] , 1'b0}), .in_29({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[145][1] }), .in_31({1'b0, 
    \dot_product_and_ReLU[17].product_terms[140] [0]}), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[141][0] }), .in_33({
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[138][0] }), .in_34({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] }),
     .out_0({\level_6_sums[19][2] [9], UNCONNECTED97, UNCONNECTED96, 
    UNCONNECTED95,  \level_6_sums[19][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP818_group_359286 WALLACE_CSA_DUMMY_OP818_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[135][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[137][0] }), .in_3({1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] , 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[167][0] , 1'b0}), .in_5({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, n_1441, n_1440}), .in_6({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] , 1'b0}), .in_7({1'b0, 
    \dot_product_and_ReLU[18].product_terms[183][1] , 1'b0}), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[174][1] }),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[173][1] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[164][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[1][81][0] }), .in_12({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[158][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, n_1439, n_1448}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[9].product_terms[152][0] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[143][0] }),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[138][0] }), .in_17({1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_18({
    \dot_product_and_ReLU[0].product_terms[191][1] , 1'b0}), .in_19({1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] , 1'b0}), .in_20({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }),
     .in_21({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[186][0] }), .in_22({1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[187][0] }), .in_23({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[184][1] }), .in_24({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[185][0] }),
     .in_25({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[178][0] }), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[179][0] }), .in_27({
    1'b0, \dot_product_and_ReLU[1].product_terms[176][0] }), .in_28({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[177][0] }), .in_29({
    1'b0, \dot_product_and_ReLU[1].product_terms[170][0] }), .in_30({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[171][1] , 1'b0}), .in_31({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[169][0] , 1'b0}),
     .in_32({1'b0, \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[161][0] }), .in_34({1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] , 1'b0}), .in_35({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}),
     .in_36({1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }),
     .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[148][0] }), .in_38({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[149][0] }), .in_39({
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }), .in_40({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[147][0] }),
     .in_41({1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 1'b0}),
     .in_42({1'b0, \dot_product_and_ReLU[0].product_terms[141][0] , 1'b0}),
     .in_43({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] , 
    1'b0}), .in_44({1'b0, \dot_product_and_ReLU[4].product_terms[133][0] }),
     .out_0({\level_6_sums[1][2] [9], UNCONNECTED100, UNCONNECTED99, 
    UNCONNECTED98,  \level_6_sums[1][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP850_group_359289 WALLACE_CSA_DUMMY_OP850_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[186][0] }),
     .in_1({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 
    1'b0}), .in_2({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] , 1'b0, 1'b0}), .in_3({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[184][1] , 1'b0}),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] }), .in_5({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[179][0] , 
    \dot_product_and_ReLU[3].product_terms[178][0] }), .in_6({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[175][0] }), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, n_1398, n_1452}), .in_8({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] , 1'b0, 1'b0}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, n_1388, n_1448}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] , 1'b0}), .in_11({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[152][0] , 1'b0}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[145][1] , 
    \dot_product_and_ReLU[2].product_terms[144][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[140] [0], 
    \dot_product_and_ReLU[0].product_terms[141][0] }), .in_14({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] }),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[132][1] , 1'b0}), .in_16({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] , 1'b0}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[191][1] }), .in_18({1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] }), .in_19({1'b0, 
    \dot_product_and_ReLU[3].product_terms[181][0] }), .in_20({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[176][0] }), .in_21({
    1'b0, \dot_product_and_ReLU[0].product_terms[177][0] , 1'b0, 1'b0}), .in_22({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[172][1] }),
     .in_23({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] , 
    1'b0}), .in_24(\dot_product_and_ReLU[3].product_terms[168][0] ), .in_25({
    \dot_product_and_ReLU[0].product_terms[169][0] , 1'b0}), .in_26({1'b0, 
    \dot_product_and_ReLU[3].product_terms[164][0] }), .in_27(
    \dot_product_and_ReLU[2].product_terms[165][0] ), .in_28({1'b0, 
    \level_1_sums[1][81][0] }), .in_29(
    \dot_product_and_ReLU[9].product_terms[163][0] ), .in_30({
    \dot_product_and_ReLU[5].product_terms[160][1] , 1'b0}), .in_31({
    \dot_product_and_ReLU[3].product_terms[161][0] , 1'b0, 1'b0}), .in_32({1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[158][0] , 1'b0, 1'b0}),
     .in_33({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[159][1] }), .in_34({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[150][0] , 1'b0}), .in_35({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[151][0] }),
     .in_36({1'b0, \dot_product_and_ReLU[1].product_terms[148][0] }), .in_37(
    \dot_product_and_ReLU[1].product_terms[149][0] ), .in_38(
    \dot_product_and_ReLU[4].product_terms[146][0] ), .in_39({
    \dot_product_and_ReLU[1].product_terms[147][0] , 1'b0}), .in_40({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[142][0] , 1'b0}), .in_41({
    1'b0, \dot_product_and_ReLU[2].product_terms[143][0] , 1'b0}), .in_42({1'b0, 
    \dot_product_and_ReLU[19].product_terms[138][0] }), .in_43({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[139][0] }), .in_44({
    1'b0, \dot_product_and_ReLU[4].product_terms[136][1] }), .in_45({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[137][0] }), .in_46(
    \dot_product_and_ReLU[0].product_terms[130][0] ), .in_47({1'b0, 
    \dot_product_and_ReLU[14].product_terms[131][0] }), .in_48({
    \dot_product_and_ReLU[9].product_terms[128][1] , 1'b0}), .in_49(
    \dot_product_and_ReLU[2].product_terms[129][0] ), .out_0({
    \level_6_sums[8][2] [9], UNCONNECTED102, UNCONNECTED101,  \level_6_sums[8][2] [6:0] }));
  WALLACE_CSA_DUMMY_OP875_group_359275 WALLACE_CSA_DUMMY_OP875_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[134][1] }),
     .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[135][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[142][0] }), .in_3({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[141][0] }),
     .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[159][1] }), .in_5({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0}), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[185][0] }), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[171][1] }),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[149][0] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] , 
    \dot_product_and_ReLU[0].product_terms[191][1] }), .in_11({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[180][0] , 
    \dot_product_and_ReLU[3].product_terms[181][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[178][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[173][1] }), .in_15({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[164][0] , 
    \dot_product_and_ReLU[2].product_terms[165][0] }), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[161][0] , 
    \dot_product_and_ReLU[5].product_terms[160][1] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[157][0] , 
    \dot_product_and_ReLU[17].product_terms[156][2] }), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[153][0] }),
     .in_19({1'b0, 1'b0, 1'b0, 1'b0, n_1391, n_1390}), .in_20({1'b0, 1'b0, 1'b0, 
    1'b0, \level_1_sums[2][73] [2], \level_1_sums[2][73] [0]}), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, n_1208, n_1404}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, n_1397, 
    n_1396}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] }), .in_24({1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[183][1] , 1'b0, 1'b0}), .in_25({
    1'b0, \dot_product_and_ReLU[0].product_terms[177][0] }), .in_26(
    \dot_product_and_ReLU[2].product_terms[174][1] ), .in_27(
    \dot_product_and_ReLU[2].product_terms[175][0] ), .in_28({1'b0, 
    \dot_product_and_ReLU[0].product_terms[169][0] }), .in_29({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[154][0] }), .in_30({
    1'b0, \dot_product_and_ReLU[0].product_terms[155][0] , 1'b0}), .in_31({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] }),
     .in_32({\dot_product_and_ReLU[19].product_terms[138][0] , 1'b0, 1'b0}),
     .in_33(\dot_product_and_ReLU[8].product_terms[139][0] ), .in_34({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[131][0] }),
     .out_0({\level_6_sums[14][2] [9], UNCONNECTED105, UNCONNECTED104, 
    UNCONNECTED103,  \level_6_sums[14][2] [5:0] }));
  WALLACE_CSA_DUMMY_OP1315_group_109833 WALLACE_CSA_DUMMY_OP1315_groupi(.in_0({
    B[247], 1'b0}), .in_1({1'b0, B[246]}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    B[221]}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, B[228]}), .in_4({1'b0, B[229], 
    1'b0}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, B[253]}), .in_6({1'b0, 1'b0, 1'b0, 
    B[237], 1'b0}), .in_7({1'b0, 1'b0, 1'b0, \level_6_sums[18][2] [9],  \level_6_sums[18][2] [5:0] }), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, n_1535, n_1534}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    B[250]}), .in_10({1'b0, B[251]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[242]}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_1517, n_1516}), .in_13({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[226]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[217]}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[212]}), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, n_1512, n_1511}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, B[203], 
    B[202]}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[201]}), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, n_1429, n_1428}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[194]}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[192]}), .in_22({1'b0, 
    1'b0, 1'b0, B[244], 1'b0}), .in_23({1'b0, 1'b0, 1'b0, 1'b0, B[245]}),
     .in_24(B[240]), .in_25({B[241], 1'b0}), .in_26({1'b0, 1'b0, 1'b0, B[235], 
    1'b0}), .in_27({1'b0, B[233], 1'b0}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, 
    B[230]}), .in_29({1'b0, 1'b0, B[231]}), .in_30({B[224], 1'b0}), .in_31({
    B[225], 1'b0}), .in_32({1'b0, 1'b0, 1'b0, B[223], 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, B[219], 1'b0}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[214]}),
     .in_35({1'b0, 1'b0, B[215]}), .in_36(B[210]), .in_37({B[211], 1'b0}),
     .in_38(B[208]), .in_39({1'b0, B[209]}), .in_40({B[204], 1'b0}), .in_41(
    B[205]), .in_42({1'b0, B[197]}), .out_0({\level_7_sums[18][1] [9], 
    UNCONNECTED107, UNCONNECTED106,  \level_7_sums[18][1] [6:0] }));
  WALLACE_CSA_DUMMY_OP1318_group_109815 WALLACE_CSA_DUMMY_OP1318_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0}), .in_1({1'b0, B[228], n_1245}), .in_2(n_1244),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, B[233]}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    B[253]}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_2631_danc, n_1495}), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[244]}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 
    B[243], 1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, B[238]}), .in_9({1'b0, 1'b0, 
    1'b0, 1'b0, B[239]}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, B[234], 1'b0}),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[222]}), .in_12({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[216]}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[212]}),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, n_1504, n_1529}), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[208]}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, B[203], B[202]}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[194]}), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, B[254]}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, B[255]}), .in_20({B[250], 
    1'b0}), .in_21({B[251], 1'b0}), .in_22({1'b0, B[248]}), .in_23({1'b0, 1'b0, 
    1'b0, B[249], 1'b0}), .in_24({1'b0, 1'b0, 1'b0, B[240], 1'b0}), .in_25({
    1'b0, B[241], 1'b0}), .in_26({1'b0, B[231], 1'b0, 1'b0}), .in_27({1'b0, 
    1'b0, 1'b0, B[226], 1'b0}), .in_28({1'b0, B[227], 1'b0}), .in_29({1'b0, 
    1'b0, 1'b0, B[224], 1'b0}), .in_30({1'b0, 1'b0, 1'b0, 1'b0, B[225]}),
     .in_31({1'b0, B[220]}), .in_32({1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_33({
    1'b0, 1'b0, 1'b0, 1'b0, B[218]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, B[219]}),
     .in_35({1'b0, 1'b0, 1'b0, 1'b0, B[214]}), .in_36({1'b0, 1'b0, 1'b0, B[215], 
    1'b0}), .in_37(B[206]), .in_38({B[207], 1'b0, 1'b0}), .in_39({1'b0, B[205]}),
     .in_40({1'b0, 1'b0, 1'b0, 1'b0, B[201]}), .in_41({1'b0, 1'b0, 1'b0, B[198], 
    1'b0}), .in_42({1'b0, B[199]}), .in_43({1'b0, 1'b0, B[196]}), .in_44({1'b0, 
    1'b0, 1'b0, 1'b0, B[197]}), .in_45({1'b0, B[192]}), .in_46({1'b0, 1'b0, 
    B[193]}), .out_0({\level_6_sums[7][3] [9], UNCONNECTED110, UNCONNECTED109, 
    UNCONNECTED108,  \level_6_sums[7][3] [5:0] }));
  WALLACE_CSA_DUMMY_OP_group_109839_6286_6339 WALLACE_CSA_DUMMY_OP_groupi(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, B[195]}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, B[218]}),
     .in_2({1'b0, B[219], 1'b0}), .in_3({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[187][0] , 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, \level_5_sums[9][4] [9],  \level_5_sums[9][4] [4:0] }), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 
    \level_4_sums[9][10] [8],  \level_4_sums[9][10] [3:0] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[248]}),
     .in_7({1'b0, 1'b0, 1'b0, 1'b0, B[242], 1'b0}), .in_8({1'b0, 1'b0, 1'b0, 
    n_1502, n_1501, n_1500}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[236]}),
     .in_10({1'b0, 1'b0, n_1552, n_1551, 1'b0, B[235]}), .in_11({1'b0, 1'b0, 
    1'b0, n_1550, n_1549, 1'b0}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, n_2667_danc, 
    n_1547}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[206]}), .in_14({1'b0, 
    1'b0, 1'b0, 1'b0,  B[202:203] }), .in_15({1'b0, 1'b0, 1'b0, n_1510, n_1509, B[201]}),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, n_1538, \level_1_sums[12][95] [0]}),
     .in_17({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[6].product_terms[188][1] }), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, n_1537, n_1536}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, B[254]}),
     .in_20({1'b0, B[255], 1'b0}), .in_21({1'b0, 1'b0, 1'b0, 1'b0, B[252]}),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, B[253]}), .in_23({1'b0, 1'b0, 1'b0, B[250], 
    1'b0}), .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[251]}), .in_25({1'b0, 1'b0, 1'b0, 
    1'b0, B[246]}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, B[247]}), .in_27({1'b0, 
    1'b0, 1'b0, B[244], 1'b0}), .in_28({1'b0, 1'b0, 1'b0, 1'b0, B[245]}),
     .in_29({1'b0, 1'b0, 1'b0, B[238], 1'b0}), .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    B[239]}), .in_31({1'b0, 1'b0, 1'b0, 1'b0, B[230]}), .in_32({1'b0, 1'b0, 
    1'b0, 1'b0, B[231]}), .in_33({1'b0, 1'b0, 1'b0, 1'b0, B[228]}), .in_34({
    1'b0, 1'b0, 1'b0, 1'b0, B[229]}), .in_35({1'b0, 1'b0, 1'b0, 1'b0, B[226]}),
     .in_36({1'b0, 1'b0, 1'b0, 1'b0, B[227]}), .in_37({1'b0, B[222]}), .in_38({
    1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_39({1'b0, 1'b0, 1'b0, 1'b0, B[220]}),
     .in_40({1'b0, 1'b0, 1'b0, 1'b0, B[221]}), .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    B[216]}), .in_42({1'b0, 1'b0, 1'b0, 1'b0, B[217]}), .in_43({1'b0, 1'b0, 
    1'b0, B[214], 1'b0}), .in_44({1'b0, 1'b0, 1'b0, B[215], 1'b0}), .in_45({
    1'b0, 1'b0, 1'b0, B[212], 1'b0}), .in_46({1'b0, 1'b0, 1'b0, B[213], 1'b0}),
     .in_47({1'b0, 1'b0, 1'b0, B[210], 1'b0}), .in_48({1'b0, 1'b0, 1'b0, B[211], 
    1'b0}), .in_49({1'b0, 1'b0, 1'b0, 1'b0, B[208]}), .in_50({1'b0, 1'b0, 
    B[209]}), .in_51({1'b0, 1'b0, 1'b0, 1'b0, B[204]}), .in_52({1'b0, B[205]}),
     .in_53({1'b0, 1'b0, 1'b0, 1'b0, B[198]}), .in_54({1'b0, 1'b0, 1'b0, B[199], 
    1'b0}), .in_55({1'b0, 1'b0, 1'b0, 1'b0, B[196]}), .in_56({1'b0, 1'b0, 
    B[197]}), .in_57({1'b0, 1'b0, 1'b0, B[192], 1'b0}), .in_58({1'b0, 1'b0, 
    1'b0, B[193], 1'b0}), .in_59({
    \dot_product_and_ReLU[3].product_terms[184][1] , 1'b0}), .in_60(
    \dot_product_and_ReLU[5].product_terms[185][0] ), .in_61({1'b0, 1'b0, 
    \dot_product_and_ReLU[8].product_terms[182][0] , 1'b0, 1'b0}), .in_62({
    1'b0, \dot_product_and_ReLU[18].product_terms[183][1] , 1'b0}), .in_63({
    1'b0, \dot_product_and_ReLU[8].product_terms[180][0] }), .in_64({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[181][0] , 1'b0}), .in_65({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[176][0] }),
     .in_66({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[177][0] , 
    1'b0}), .out_0({\level_7_sums[9][1] [9], UNCONNECTED111,  \level_7_sums[9][1] [7:0] }));
  WALLACE_CSA_DUMMY_OP_group_109839 WALLACE_CSA_DUMMY_OP_groupi4116(.in_0({
    \dot_product_and_ReLU[19].product_terms[46][2] , 1'b0}), .in_1({
    \dot_product_and_ReLU[3].product_terms[47][1] , 1'b0}), .in_2({1'b0, 1'b0, 
    1'b0, 1'b0, n_1241, n_1240, \dot_product_and_ReLU[0].product_terms[41][0] }),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[63][1] , 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, n_1494, n_2773_danc}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1493, 
    n_1492}), .in_6({1'b0, 1'b0, 1'b0, n_1491, n_1490, n_1489}), .in_7({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[39][0] }),
     .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[31][1] }), .in_9({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[26][2] , 1'b0}), .in_10({1'b0, 
    \dot_product_and_ReLU[0].product_terms[27][0] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[14][1] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] , 
    \dot_product_and_ReLU[0].product_terms[13][0] }), .in_14({
    \dot_product_and_ReLU[19].product_terms[60][2] , 1'b0}), .in_15({
    \dot_product_and_ReLU[15].product_terms[61][1] , 1'b0}), .in_16({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[37][1] }), .in_17({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[34][0] , 1'b0}), .in_18({
    1'b0, \dot_product_and_ReLU[2].product_terms[35][0] , 1'b0}), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }), .in_20({
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[33][0] }), .in_21({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[28][0] }), .in_22({
    1'b0, \dot_product_and_ReLU[0].product_terms[29][0] }), .in_23({1'b0, 
    \dot_product_and_ReLU[0].product_terms[22][0] }), .in_24({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_25({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }), .in_26({
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }), .in_27({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[16][0] }), .in_28({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[17][1] , 1'b0}),
     .in_29({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[11][1] , 
    1'b0}), .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[8][0] }), .in_31({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[6].product_terms[9][0] }), .in_32({1'b0, 
    \dot_product_and_ReLU[0].product_terms[6][2] , 1'b0, 1'b0}), .in_33({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[7][0] }), .in_34(
    \dot_product_and_ReLU[2].product_terms[4][0] ), .in_35(
    \dot_product_and_ReLU[0].product_terms[5][0] ), .in_36({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[3][0] , 1'b0}), .in_37(
    \dot_product_and_ReLU[0].product_terms[0][0] ), .in_38(
    \dot_product_and_ReLU[4].product_terms[1][0] ), .out_0({
    \level_6_sums[0][0] [9], UNCONNECTED114, UNCONNECTED113, UNCONNECTED112,  \level_6_sums[0][0] [5:0] }));
  WALLACE_CSA_DUMMY_OP_group_109839_6286 WALLACE_CSA_DUMMY_OP_groupi4212(.in_0({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[88][1] }), .in_1({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[113][1] }), .in_2({1'b0, 1'b0, 
    1'b0, \level_6_sums[7][0] [9],  \level_6_sums[7][0] [5:0] }), .in_3({1'b0, 1'b0, 1'b0, 
    \level_6_sums[7][3] [9],  \level_6_sums[7][3] [5:0] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_1389, 
    n_1408}), .in_5({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[17].product_terms[124][0] , 1'b0, 1'b0}), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, n_2925_danc, n_2926_danc}), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[117][0] }),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] }), .in_10({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}),
     .in_11({1'b0, 1'b0, 1'b0, \level_1_sums[3][46] [4], 
    \level_1_sums[3][46] [0], \dot_product_and_ReLU[8].product_terms[92][1] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[84][0] , 
    \dot_product_and_ReLU[1].product_terms[85][0] }), .in_13({1'b0, 1'b0, 1'b0, 
    n_2862_danc, n_1436, \dot_product_and_ReLU[10].product_terms[80][0] }),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[10].product_terms[78][1] , 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[6].product_terms[188][1] , 1'b0}),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[186][0] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0,  \level_1_sums[7][92] [1:0] }), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[183][1] }), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, n_1212, n_1536}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[174][1] }), .in_21({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[173][1] }),
     .in_22({1'b0, 1'b0, 1'b0, 1'b0, n_1453, n_1452}), .in_23({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[9].product_terms[163][0] , 
    \level_1_sums[1][81][0] }), .in_24({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[161][0] }), .in_25({1'b0, 1'b0, 
    1'b0, 1'b0, n_1393, n_1392}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, n_1388, 
    n_1448}), .in_27({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] , 1'b0}), .in_28({1'b0, 
    1'b0, 1'b0, 1'b0, n_1387, n_1390}), .in_29({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[146][0] }), .in_30({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 
    \dot_product_and_ReLU[2].product_terms[144][0] }), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[138][0] , 1'b0}),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[136][1] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[133][0] }),
     .in_34({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[130][0] }), .in_35({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_36({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[127][0] }),
     .in_37({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[111][0] }), .in_38({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[109][1] , 1'b0}), .in_39({
    1'b0, \dot_product_and_ReLU[16].product_terms[107][0] , 1'b0}), .in_40({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[16].product_terms[102][2] }),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[103][0] }), .in_42(
    \dot_product_and_ReLU[0].product_terms[100][0] ), .in_43(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .in_44({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[98][1] , 1'b0}), .in_45({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] }), .in_46({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[97][0] }),
     .in_47({1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[94][1] , 1'b0, 
    1'b0}), .in_48({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[95][0] }), .in_49({1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[86][0] }), .in_50(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .in_51({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[82][0] }), .in_52({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}), .in_53({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[76][0] , 1'b0}), .in_54({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[77][0] }),
     .in_55({1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] }), .in_56({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[75][0] }), .in_57({
    1'b0, \dot_product_and_ReLU[5].product_terms[72][0] }), .in_58({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[73][0] }), .in_59({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[70][0] , 1'b0}), .in_60({
    1'b0, \dot_product_and_ReLU[16].product_terms[71][0] }), .in_61({1'b0, 
    \dot_product_and_ReLU[4].product_terms[68][0] }), .in_62({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[1].product_terms[69][1] }), .in_63({1'b0, 
    \dot_product_and_ReLU[0].product_terms[66][0] }), .in_64({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[67][0] }), .in_65({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[64][1] , 1'b0}), .in_66({1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] , 1'b0}), .in_67({1'b0, 
    \dot_product_and_ReLU[4].product_terms[190][1] }), .in_68(
    \dot_product_and_ReLU[0].product_terms[191][1] ), .in_69({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[8].product_terms[180][0] }), .in_70({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[181][0] }),
     .in_71(\dot_product_and_ReLU[1].product_terms[176][0] ), .in_72({1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[177][0] }), .in_73({
    \dot_product_and_ReLU[3].product_terms[168][0] , 1'b0}), .in_74({
    \dot_product_and_ReLU[0].product_terms[169][0] , 1'b0}), .in_75({1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] , 1'b0}), .in_76({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[167][0] }),
     .in_77({1'b0, \dot_product_and_ReLU[2].product_terms[165][0] , 1'b0}),
     .in_78(\dot_product_and_ReLU[9].product_terms[152][0] ), .in_79(
    \dot_product_and_ReLU[18].product_terms[153][0] ), .in_80({1'b0, 
    \dot_product_and_ReLU[1].product_terms[149][0] }), .in_81(
    \dot_product_and_ReLU[2].product_terms[134][1] ), .in_82({1'b0, 
    \dot_product_and_ReLU[1].product_terms[135][0] }), .in_83({1'b0, 
    \dot_product_and_ReLU[9].product_terms[128][1] , 1'b0}), .in_84({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[129][0] , 1'b0}),
     .out_0({\level_8_sums[7] [8], UNCONNECTED115,  \level_8_sums[7] [7:0] }));
  csa_tree_dot_product_and_ReLU_0__product_terms_gen_255__final_adder_adder_inst_add_47_23_group_359257 
    csa_tree_dot_product_and_ReLU_0__product_terms_gen_255__final_adder_adder_inst_add_47_23_groupi(
    .in_0({1'b0, 1'b0, 1'b0, \level_6_sums[0][0] [9],  \level_6_sums[0][0] [5:0] }), .in_1({1'b0, 1'b0, 1'b0, 
    \level_6_sums[0][3] [9],  \level_6_sums[0][3] [5:0] }), .in_2({1'b0, 1'b0, 1'b0, n_1238, n_1237, n_1236, 
    n_1235}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[183][1] }), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, n_1234, n_1233, n_1232}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \level_1_sums[1][81][0] , 1'b0}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    n_1460, n_1459}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[126][1] }), .in_8({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] }), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, n_2925_danc, n_2926_danc}), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[112][2] }), .in_11({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[108][0] , 
    1'b0}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] }), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[98][1] }), .in_14({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[90][0] }), .in_15({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[86][0] }), .in_16({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[72][0] }),
     .in_17({1'b0, 1'b0, 1'b0, n_1458, n_1457, 1'b0}), .in_18({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[68][0] }), .in_19({1'b0, 
    1'b0, 1'b0, 1'b0, n_1456, n_1455}), .in_20({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[65][0] }), .in_21({1'b0, 1'b0, 1'b0, 
    1'b0, n_1454, \level_1_sums[16][87] [1]}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[172][1] }), .in_23({1'b0, 
    1'b0, 1'b0, 1'b0, n_1453, n_1452}), .in_24({1'b0, 1'b0, 1'b0, n_1451, 
    n_1450, \dot_product_and_ReLU[2].product_terms[165][0] }), .in_25({1'b0, 
    1'b0, 1'b0, 1'b0, n_1449, n_1448}), .in_26({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[18].product_terms[153][0] }), .in_27({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[146][0] }),
     .in_28({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[134][1] }), .in_29({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[132][1] }),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[130][0] }), .in_31({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[9].product_terms[128][1] }),
     .in_32({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[122][0] }), .in_33({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[123][1] }), .in_34({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] , 1'b0}),
     .in_35({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[119][0] }), .in_36({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[117][0] , 1'b0}), .in_37({
    1'b0, \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}), .in_38({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] , 1'b0}),
     .in_39({1'b0, \dot_product_and_ReLU[7].product_terms[111][0] }), .in_40({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}),
     .in_41({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[105][0] }), .in_42({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[96][0] }), .in_43({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[97][0] }), .in_44({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[94][1] , 1'b0}),
     .in_45({1'b0, \dot_product_and_ReLU[2].product_terms[95][0] , 1'b0}),
     .in_46(\dot_product_and_ReLU[8].product_terms[92][1] ), .in_47(
    \dot_product_and_ReLU[0].product_terms[93][0] ), .in_48({1'b0, 
    \dot_product_and_ReLU[0].product_terms[88][1] , 1'b0}), .in_49({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[13].product_terms[89][0] , 1'b0}), .in_50({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}),
     .in_51({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[85][0] }), .in_52(
    \dot_product_and_ReLU[4].product_terms[82][0] ), .in_53({
    \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0}), .in_54({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[10].product_terms[80][0] }), .in_55({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[81][0] }),
     .in_56({1'b0, \dot_product_and_ReLU[0].product_terms[76][0] }), .in_57({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[77][0] , 1'b0}),
     .in_58({1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] }), .in_59({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[75][0] }), .in_60({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[190][1] }),
     .in_61({1'b0, \dot_product_and_ReLU[0].product_terms[191][1] , 1'b0}),
     .in_62({1'b0, \dot_product_and_ReLU[0].product_terms[189][0] }), .in_63({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[18].product_terms[186][0] , 1'b0}),
     .in_64({1'b0, \dot_product_and_ReLU[0].product_terms[187][0] }), .in_65({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[184][1] }),
     .in_66({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[5].product_terms[185][0] , 
    1'b0}), .in_67({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[169][0] }), .in_68({1'b0, 
    \dot_product_and_ReLU[4].product_terms[166][0] }), .in_69({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[167][0] }), .in_70({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[158][0] }),
     .in_71({1'b0, \dot_product_and_ReLU[0].product_terms[159][1] , 1'b0}),
     .in_72({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[14].product_terms[154][0] }), .in_73({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[155][0] }), .in_74({
    1'b0, \dot_product_and_ReLU[0].product_terms[150][0] }), .in_75({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[3].product_terms[151][0] , 1'b0}), .in_76({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[149][0] , 1'b0}),
     .in_77({1'b0, \dot_product_and_ReLU[2].product_terms[144][0] }), .in_78({
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[145][1] , 1'b0}),
     .in_79({\dot_product_and_ReLU[19].product_terms[138][0] , 1'b0}), .in_80(
    \dot_product_and_ReLU[8].product_terms[139][0] ), .in_81({1'b0, 
    \dot_product_and_ReLU[4].product_terms[136][1] }), .in_82({1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[137][0] , 1'b0, 1'b0}), .out_0({
    \level_8_sums[0] [8], UNCONNECTED116,  \level_8_sums[0] [7:0] }));
  csa_tree_dot_product_and_ReLU_1__product_terms_gen_127__adder_32s_adder_inst_add_38_20_group_100063 
    csa_tree_dot_product_and_ReLU_1__product_terms_gen_127__adder_32s_adder_inst_add_38_20_groupi(
    .in_0({1'b0, \dot_product_and_ReLU[0].product_terms[122][0] }), .in_1({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[123][1] , 1'b0}), .in_2(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .in_3(
    \dot_product_and_ReLU[0].product_terms[119][0] ), .in_4({1'b0, 1'b0, 1'b0, 
    1'b0, n_1447, n_1446}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1445, n_1444}),
     .in_6({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[100][0] , 1'b0}), .in_7({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[14].product_terms[99][0] }), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[5].product_terms[96][0] }), .in_9({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }),
     .in_11({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[110][0] }), .in_12({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[7].product_terms[111][0] }), .in_13({
    1'b0, \dot_product_and_ReLU[0].product_terms[106][0] }), .in_14({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[16].product_terms[107][0] , 1'b0}), .in_15({
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[104] [1]}), .in_16({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[105][0] , 1'b0}),
     .in_17({\dot_product_and_ReLU[16].product_terms[102][2] , 1'b0}), .in_18({
    \dot_product_and_ReLU[7].product_terms[103][0] , 1'b0}), .out_0({
    \level_5_sums[1][3] [9], UNCONNECTED120, UNCONNECTED119, UNCONNECTED118, 
    UNCONNECTED117,  \level_5_sums[1][3] [4:0] }));
  csa_tree_dot_product_and_ReLU_1__product_terms_gen_255__adder_64s_adder_inst_add_47_23_group_109831 
    csa_tree_dot_product_and_ReLU_1__product_terms_gen_255__adder_64s_adder_inst_add_47_23_groupi(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, n_1503, n_1525}), .in_1({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, B[248]}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, n_1533, n_1532}),
     .in_3({1'b0, 1'b0, n_1554, n_1553,  B[242:243] }), .in_4({1'b0, 1'b0, 1'b0, n_1502, 
    n_1501, n_1500}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, n_1499, n_1498}), .in_6({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[234]}), .in_7({1'b0, 1'b0, 1'b0, B[228], 
    1'b0, 1'b0}), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B[227]}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[223]}), .in_10({1'b0, 1'b0, 1'b0, 1'b0, n_1497, 
    n_1513}), .in_11({1'b0, 1'b0, 1'b0, n_1544, n_1543, B[216]}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, B[214], 1'b0}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[212]}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, n_1504, n_1529}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, B[207]}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    B[204]}), .in_17({1'b0, 1'b0, 1'b0, 1'b0, B[202]}), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, B[200]}), .in_19({1'b0, 1'b0, 1'b0, n_1508, n_1507, n_1527}),
     .in_20({1'b0, 1'b0, 1'b0, 1'b0, B[254]}), .in_21({1'b0, 1'b0, 1'b0, B[255], 
    1'b0}), .in_22({1'b0, 1'b0, 1'b0, 1'b0, B[252]}), .in_23({1'b0, B[253]}),
     .in_24({1'b0, 1'b0, 1'b0, 1'b0, B[247]}), .in_25({1'b0, 1'b0, B[238]}),
     .in_26({1'b0, 1'b0, 1'b0, B[239], 1'b0}), .in_27({B[232], 1'b0}), .in_28({
    B[233], 1'b0}), .in_29({1'b0, B[230]}), .in_30({1'b0, 1'b0, 1'b0, B[231], 
    1'b0}), .in_31({1'b0, 1'b0, 1'b0, 1'b0, B[224]}), .in_32({1'b0, 1'b0, 1'b0, 
    B[225], 1'b0}), .in_33({1'b0, B[218]}), .in_34({1'b0, 1'b0, 1'b0, 1'b0, 
    B[219]}), .in_35({1'b0, 1'b0, 1'b0, 1'b0, B[208]}), .in_36({1'b0, 1'b0, 
    1'b0, 1'b0, B[209]}), .in_37({1'b0, B[198]}), .in_38({1'b0, 1'b0, 1'b0, 
    1'b0, B[199]}), .in_39({1'b0, 1'b0, B[196]}), .in_40({1'b0, 1'b0, 1'b0, 
    1'b0, B[197]}), .in_41({1'b0, 1'b0, B[192]}), .in_42({1'b0, 1'b0, 1'b0, 
    1'b0, B[193]}), .out_0({\level_6_sums[1][3] [9], UNCONNECTED123, 
    UNCONNECTED122, UNCONNECTED121,  \level_6_sums[1][3] [5:0] }));
  csa_tree_dot_product_and_ReLU_2__product_terms_gen_127__adder_64s_adder_inst_add_47_23_group_100071 
    csa_tree_dot_product_and_ReLU_2__product_terms_gen_127__adder_64s_adder_inst_add_47_23_groupi(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, \level_3_sums[2][12][3] , 
    \level_3_sums[2][12][2] , \level_3_sums[2][12][1] , 
    \level_3_sums[2][12][0] }), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[122][0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[110][0] }), .in_3({1'b0, 
    1'b0, 1'b0, 1'b0, n_1445, n_1444}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[0].product_terms[106][0] }), .in_5({1'b0, 1'b0, 1'b0, 
    n_1438, n_1437, \dot_product_and_ReLU[0].product_terms[105][0] }), .in_6({
    1'b0, 1'b0, 1'b0, n_1435, n_2928_danc, 
    \dot_product_and_ReLU[2].product_terms[95][0] }), .in_7({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[88][1] }), .in_8({1'b0, 
    1'b0, 1'b0, n_2862_danc, n_1436, 
    \dot_product_and_ReLU[10].product_terms[80][0] }), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[10].product_terms[78][1] }), .in_10({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[79][0] }), .in_11({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \level_1_sums[4][37][1] }), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[69][1] }),
     .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[64][1] }), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[4].product_terms[127][0] }), .in_15(
    \dot_product_and_ReLU[17].product_terms[124][0] ), .in_16(
    \dot_product_and_ReLU[4].product_terms[125][1] ), .in_17({1'b0, 
    \dot_product_and_ReLU[2].product_terms[121][1] , 1'b0}), .in_18({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] , 1'b0}),
     .in_19({1'b0, \dot_product_and_ReLU[0].product_terms[119][0] , 1'b0}),
     .in_20(\dot_product_and_ReLU[2].product_terms[116][0] ), .in_21(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .in_22({1'b0, 
    \dot_product_and_ReLU[0].product_terms[114][1] , 1'b0}), .in_23({1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }),
     .in_24({1'b0, 1'b0, \dot_product_and_ReLU[17].product_terms[112][2] }),
     .in_25({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[113][1] , 
    1'b0}), .in_26({1'b0, \dot_product_and_ReLU[0].product_terms[93][0] }),
     .in_27({1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[90][0] }),
     .in_28({1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[91][1] , 
    1'b0}), .in_29({1'b0, \dot_product_and_ReLU[3].product_terms[84][0] , 1'b0}),
     .in_30({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[85][0] }), .in_31({1'b0, 
    \dot_product_and_ReLU[4].product_terms[82][0] }), .in_32({1'b0, 1'b0, 
    \dot_product_and_ReLU[3].product_terms[83][0] , 1'b0, 1'b0}), .in_33(
    \dot_product_and_ReLU[5].product_terms[72][0] ), .in_34(
    \dot_product_and_ReLU[1].product_terms[73][0] ), .in_35({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[2].product_terms[70][0] }), .in_36({1'b0, 
    \dot_product_and_ReLU[16].product_terms[71][0] , 1'b0}), .in_37({
    \dot_product_and_ReLU[0].product_terms[66][0] , 1'b0}), .in_38(
    \dot_product_and_ReLU[2].product_terms[67][0] ), .out_0({
    \level_6_sums[2][1] [9], UNCONNECTED126, UNCONNECTED125, UNCONNECTED124,  \level_6_sums[2][1] [5:0] }));
  csa_tree_dot_product_and_ReLU_14__product_terms_gen_127__adder_128s_adder_inst_add_47_23_group_106211 
    csa_tree_dot_product_and_ReLU_14__product_terms_gen_127__adder_128s_adder_inst_add_47_23_groupi(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, \level_5_sums[14][2] [9],  \level_5_sums[14][2] [4:0] }), .in_1({1'b0, 
    1'b0, 1'b0, 1'b0, \level_4_sums[14][6] [8],  \level_4_sums[14][6] [3:0] }), .in_2({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[3].product_terms[123][1] }), .in_3({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[30][1] , 1'b0}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[126][1] , 1'b0}), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[125][1] , 
    \dot_product_and_ReLU[17].product_terms[124][0] }), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[118][0] }), .in_7({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[63][1] , 
    \dot_product_and_ReLU[1].product_terms[62][0] }), .in_8({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[1].product_terms[55][0] , n_1433, n_1432}), .in_9({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[52][0] }), .in_10({1'b0, 1'b0, 
    n_1485, n_2818_danc, \dot_product_and_ReLU[2].product_terms[44][1] , 
    \dot_product_and_ReLU[3].product_terms[45][1] }), .in_11({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[42][1] , 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[40][0] }),
     .in_13({1'b0, 1'b0, 1'b0, n_2950_danc, n_1414, 
    \dot_product_and_ReLU[8].product_terms[36][0] }), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[27][0] , 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[24][0] }),
     .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[16].product_terms[12][0] }), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, n_2980_danc, n_2981_danc}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[0].product_terms[8][0] }), .in_19({1'b0, 1'b0, 
    1'b0, n_1470, n_1469, \dot_product_and_ReLU[2].product_terms[4][0] }),
     .in_20({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[2].product_terms[116][0] }), .in_21({1'b0, 
    \dot_product_and_ReLU[2].product_terms[117][0] }), .in_22({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[114][1] }), .in_23({
    1'b0, \dot_product_and_ReLU[1].product_terms[115][0] }), .in_24({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[17].product_terms[112][2] , 1'b0}), .in_25({
    1'b0, \dot_product_and_ReLU[2].product_terms[113][1] }), .in_26({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[19].product_terms[60][2] }), .in_27({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[15].product_terms[61][1] }),
     .in_28({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[59][1] }), .in_29({1'b0, 
    \dot_product_and_ReLU[1].product_terms[56][1] }), .in_30({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[7].product_terms[57][2] , 1'b0}), .in_31({1'b0, 1'b0, 
    \dot_product_and_ReLU[11].product_terms[50][0] }), .in_32({1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[5].product_terms[51][1] , 1'b0}), .in_33(
    \dot_product_and_ReLU[19].product_terms[48][1] ), .in_34({1'b0, 
    \dot_product_and_ReLU[0].product_terms[49][0] }), .in_35({1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[19].product_terms[46][2] , 1'b0}), .in_36({1'b0, 
    \dot_product_and_ReLU[3].product_terms[47][1] }), .in_37({1'b0, 1'b0, 1'b0, 
    1'b0, \dot_product_and_ReLU[7].product_terms[38][1] }), .in_38({1'b0, 
    \dot_product_and_ReLU[0].product_terms[39][0] , 1'b0}), .in_39({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[34][0] }), .in_40({1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[35][0] , 1'b0}), .in_41({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[8].product_terms[32][1] }),
     .in_42({1'b0, \dot_product_and_ReLU[2].product_terms[33][0] , 1'b0, 1'b0}),
     .in_43({1'b0, \dot_product_and_ReLU[0].product_terms[23][0] }), .in_44({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[2].product_terms[21][1] }),
     .in_45({1'b0, \dot_product_and_ReLU[14].product_terms[18][0] }), .in_46({
    1'b0, 1'b0, 1'b0, 1'b0, \dot_product_and_ReLU[1].product_terms[19][1] }),
     .in_47({1'b0, 1'b0, \dot_product_and_ReLU[0].product_terms[17][1] }),
     .in_48({1'b0, 1'b0, 1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[15][0] }), .in_49(
    \dot_product_and_ReLU[0].product_terms[6][2] ), .in_50({
    \dot_product_and_ReLU[7].product_terms[7][0] , 1'b0}), .in_51({1'b0, 1'b0, 
    1'b0, 1'b0, \dot_product_and_ReLU[4].product_terms[3][0] }), .in_52({1'b0, 
    \dot_product_and_ReLU[0].product_terms[0][0] }), .in_53({1'b0, 1'b0, 
    \dot_product_and_ReLU[4].product_terms[1][0] , 1'b0, 1'b0}), .out_0({
    \level_7_sums[14][0] [9], UNCONNECTED128, UNCONNECTED127,  \level_7_sums[14][0] [6:0] }));
  INVX1 g16309(.Y(n_1212), .A(n_1243));
  INVX1 g16310(.Y(n_1453), .A(n_1225));
  INVX1 g16313(.Y(n_1214), .A(n_1246));
  INVX1 g16308(.Y(n_1406), .A(n_1222));
  INVX1 g16311(.Y(n_1216), .A(n_1239));
  INVX1 g16314(.Y(n_1215), .A(n_1221));
  INVX1 g16315(.Y(n_1465), .A(n_1226));
  INVX1 g16312(.Y(n_1213), .A(n_1220));
  INVX1 g16317(.Y(n_1209), .A(n_1242));
  INVX1 g16316(.Y(n_1208), .A(n_1228));
  INVX1 g16323(.Y(n_1207), .A(\dot_product_and_ReLU[1].product_terms[176][0] ));
  INVX1 g16336(.Y(n_1206), .A(\dot_product_and_ReLU[0].product_terms[94][1] ));
  INVX1 g16328(.Y(n_1205), .A(\dot_product_and_ReLU[0].product_terms[150][0] ));
  INVX1 g16320(.Y(n_1204), .A(\dot_product_and_ReLU[7].product_terms[111][0] ));
  INVX1 g16319(.Y(n_1203), .A(\dot_product_and_ReLU[4].product_terms[133][0] ));
  INVX1 g16324(.Y(n_1202), .A(\dot_product_and_ReLU[0].product_terms[76][0] ));
  INVX1 g16329(.Y(n_1201), .A(\dot_product_and_ReLU[3].product_terms[45][1] ));
  INVX1 g16334(.Y(n_1200), .A(\dot_product_and_ReLU[2].product_terms[44][1] ));
  INVX1 g16331(.Y(n_1199), .A(\dot_product_and_ReLU[0].product_terms[41][0] ));
  INVX1 g16322(.Y(n_1198), .A(\dot_product_and_ReLU[1].product_terms[132][1] ));
  INVX1 g16325(.Y(n_1197), .A(\dot_product_and_ReLU[7].product_terms[7][0] ));
  INVX1 g16326(.Y(n_1196), .A(\dot_product_and_ReLU[0].product_terms[6][2] ));
  INVX1 g16318(.Y(n_1195), .A(\dot_product_and_ReLU[19].product_terms[26][2] ));
  INVX1 g16327(.Y(n_1194), .A(\dot_product_and_ReLU[2].product_terms[40][0] ));
  INVX1 g16332(.Y(n_1193), .A(\dot_product_and_ReLU[0].product_terms[177][0] ));
  INVX1 g16321(.Y(n_1192), .A(\dot_product_and_ReLU[7].product_terms[16][0] ));
  INVX1 g16337(.Y(n_1191), .A(\dot_product_and_ReLU[3].product_terms[151][0] ));
  INVX1 g16335(.Y(n_1190), .A(\dot_product_and_ReLU[2].product_terms[95][0] ));
  INVX1 g16333(.Y(n_1211), .A(B[242]));
  INVX1 g16330(.Y(n_1210), .A(B[243]));
  DFFRHQX1 \out_reg_reg[2][5] (.Q(out[23]), .D(n_1182), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][7] (.Q(out[25]), .D(n_1181), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][8] (.Q(out[26]), .D(n_1189), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][1] (.Q(out[19]), .D(n_1183), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][6] (.Q(out[24]), .D(n_1188), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][4] (.Q(out[22]), .D(n_1187), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][0] (.Q(out[18]), .D(n_1186), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][3] (.Q(out[21]), .D(n_1185), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[2][2] (.Q(out[20]), .D(n_1184), .RN(rst_n), .CK(clk));
  NOR2BX1 g16338(.Y(n_1189), .AN(\final_sums[2] [8]), .B(\final_sums[2] [9]));
  NOR2BX1 g16339(.Y(n_1188), .AN(\final_sums[2] [6]), .B(\final_sums[2] [9]));
  NOR2BX1 g16340(.Y(n_1187), .AN(\final_sums[2] [4]), .B(\final_sums[2] [9]));
  NOR2BX1 g16341(.Y(n_1186), .AN(\final_sums[2] [0]), .B(\final_sums[2] [9]));
  NOR2BX1 g16342(.Y(n_1185), .AN(\final_sums[2] [3]), .B(\final_sums[2] [9]));
  NOR2BX1 g16343(.Y(n_1184), .AN(\final_sums[2] [2]), .B(\final_sums[2] [9]));
  NOR2BX1 g16344(.Y(n_1183), .AN(\final_sums[2] [1]), .B(\final_sums[2] [9]));
  NOR2BX1 g16345(.Y(n_1182), .AN(\final_sums[2] [5]), .B(\final_sums[2] [9]));
  NOR2BX1 g16346(.Y(n_1181), .AN(\final_sums[2] [7]), .B(\final_sums[2] [9]));
  DFFRHQX1 \out_reg_reg[4][4] (.Q(out[40]), .D(n_1178), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][6] (.Q(out[42]), .D(n_1179), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][7] (.Q(out[43]), .D(n_1173), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][0] (.Q(out[36]), .D(n_1180), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][2] (.Q(out[38]), .D(n_1176), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][5] (.Q(out[41]), .D(n_1175), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][3] (.Q(out[39]), .D(n_1174), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[4][1] (.Q(out[37]), .D(n_1177), .RN(rst_n), .CK(clk));
  NOR2BX1 g16347(.Y(n_1180), .AN(\final_sums[4] [0]), .B(\final_sums[4] [9]));
  NOR2BX1 g16348(.Y(n_1179), .AN(\final_sums[4] [6]), .B(\final_sums[4] [9]));
  NOR2BX1 g16349(.Y(n_1178), .AN(\final_sums[4] [4]), .B(\final_sums[4] [9]));
  NOR2BX1 g16350(.Y(n_1177), .AN(\final_sums[4] [1]), .B(\final_sums[4] [9]));
  NOR2BX1 g16351(.Y(n_1176), .AN(\final_sums[4] [2]), .B(\final_sums[4] [9]));
  NOR2BX1 g16352(.Y(n_1175), .AN(\final_sums[4] [5]), .B(\final_sums[4] [9]));
  NOR2BX1 g16353(.Y(n_1174), .AN(\final_sums[4] [3]), .B(\final_sums[4] [9]));
  NOR2BX1 g16354(.Y(n_1173), .AN(\final_sums[4] [7]), .B(\final_sums[4] [9]));
  DFFRHQX1 \out_reg_reg[5][4] (.Q(out[49]), .D(n_1170), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][6] (.Q(out[51]), .D(n_1171), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][7] (.Q(out[52]), .D(n_1165), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][0] (.Q(out[45]), .D(n_1172), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][2] (.Q(out[47]), .D(n_1168), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][5] (.Q(out[50]), .D(n_1167), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][3] (.Q(out[48]), .D(n_1166), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[5][1] (.Q(out[46]), .D(n_1169), .RN(rst_n), .CK(clk));
  NOR2BX1 g16355(.Y(n_1172), .AN(\final_sums[5] [0]), .B(\final_sums[5] [9]));
  NOR2BX1 g16356(.Y(n_1171), .AN(\final_sums[5] [6]), .B(\final_sums[5] [9]));
  NOR2BX1 g16357(.Y(n_1170), .AN(\final_sums[5] [4]), .B(\final_sums[5] [9]));
  NOR2BX1 g16358(.Y(n_1169), .AN(\final_sums[5] [1]), .B(\final_sums[5] [9]));
  NOR2BX1 g16359(.Y(n_1168), .AN(\final_sums[5] [2]), .B(\final_sums[5] [9]));
  NOR2BX1 g16360(.Y(n_1167), .AN(\final_sums[5] [5]), .B(\final_sums[5] [9]));
  NOR2BX1 g16361(.Y(n_1166), .AN(\final_sums[5] [3]), .B(\final_sums[5] [9]));
  NOR2BX1 g16362(.Y(n_1165), .AN(\final_sums[5] [7]), .B(\final_sums[5] [9]));
  AO21XL g17798(.Y(\level_5_sums[14][2] [4]), .A0(n_1153), .A1(n_1164), .B0(
    \level_5_sums[14][2] [9]));
  NOR2X1 g17799(.Y(\level_5_sums[14][2] [9]), .A(n_1153), .B(n_1164));
  ADDFX1 g17800(.CO(n_1164), .S(\level_5_sums[14][2] [3]), .A(n_1152), .B(n_1157),
     .CI(n_1162));
  INVX1 g17801(.Y(\level_4_sums[14][6] [8]), .A(n_1163));
  ADDFX1 g17802(.CO(n_1163), .S(\level_4_sums[14][6] [3]), .A(n_1102), .B(n_1143),
     .CI(n_1161));
  ADDFX1 g17803(.CO(n_1162), .S(\level_5_sums[14][2] [2]), .A(n_1155), .B(n_1158),
     .CI(n_1160));
  ADDFX1 g17804(.CO(n_1161), .S(\level_4_sums[14][6] [2]), .A(n_1150), .B(n_1144),
     .CI(n_1159));
  ADDFX1 g17805(.CO(n_1160), .S(\level_5_sums[14][2] [1]), .A(n_1149), .B(n_1154),
     .CI(n_1156));
  ADDFX1 g17806(.CO(n_1159), .S(\level_4_sums[14][6] [1]), .A(n_1122), .B(n_1147),
     .CI(n_1151));
  ADDFX1 g17807(.CO(n_1157), .S(n_1158), .A(n_1139), .B(n_1148), .CI(n_1146));
  ADDFX1 g17808(.CO(n_1155), .S(n_1156), .A(n_1132), .B(n_1140), .CI(n_1141));
  ADDFX1 g17809(.CO(n_1154), .S(\level_5_sums[14][2] [0]), .A(n_1128), .B(n_1124),
     .CI(n_1142));
  ADDHX1 g17810(.CO(n_1153), .S(n_1152), .A(n_1125), .B(n_1145));
  ADDFX1 g17811(.CO(n_1150), .S(n_1151), .A(n_1129), .B(n_1137), .CI(n_1135));
  ADDFX1 g17812(.CO(n_1148), .S(n_1149), .A(n_1127), .B(n_1123), .CI(n_1133));
  ADDFX1 g17813(.CO(n_1147), .S(\level_4_sums[14][6] [0]), .A(n_1130), .B(n_1138),
     .CI(n_1136));
  ADDFX1 g17814(.CO(n_1145), .S(n_1146), .A(n_1088), .B(n_1131), .CI(n_1126));
  ADDFX1 g17815(.CO(n_1143), .S(n_1144), .A(n_1111), .B(n_1087), .CI(n_1121));
  ADDFX1 g17816(.CO(n_1141), .S(n_1142), .A(n_1089), .B(n_2871_danc), .CI(n_1134));
  ADDFX1 g17817(.CO(n_1139), .S(n_1140), .A(
    \dot_product_and_ReLU[5].product_terms[75][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[77][0] ), .CI(n_2870_danc));
  ADDFX1 g17818(.CO(n_1137), .S(n_1138), .A(
    \dot_product_and_ReLU[3].product_terms[110][0] ), .B(n_1091), .CI(n_1097));
  ADDFX1 g17819(.CO(n_1135), .S(n_1136), .A(n_1094), .B(
    \dot_product_and_ReLU[7].product_terms[103][0] ), .CI(n_1119));
  ADDFX1 g17820(.CO(n_1133), .S(n_1134), .A(
    \dot_product_and_ReLU[0].product_terms[94][1] ), .B(n_1099), .CI(n_1095));
  ADDFX1 g17821(.CO(n_1131), .S(n_1132), .A(
    \dot_product_and_ReLU[0].product_terms[65][0] ), .B(n_1090), .CI(n_1100));
  ADDFX1 g17822(.CO(n_1129), .S(n_1130), .A(
    \dot_product_and_ReLU[14].product_terms[99][0] ), .B(n_1098), .CI(
    \dot_product_and_ReLU[4].product_terms[98][1] ));
  ADDFX1 g17823(.CO(n_1127), .S(n_1128), .A(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .B(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .CI(
    \dot_product_and_ReLU[0].product_terms[66][0] ));
  ADDFX1 g17824(.CO(n_1125), .S(n_1126), .A(
    \dot_product_and_ReLU[3].product_terms[86][0] ), .B(n_1093), .CI(
    \dot_product_and_ReLU[4].product_terms[82][0] ));
  ADDFX1 g17825(.CO(n_1123), .S(n_1124), .A(
    \dot_product_and_ReLU[0].product_terms[88][1] ), .B(n_1096), .CI(
    \dot_product_and_ReLU[1].product_terms[73][0] ));
  OAI2BB1X1 g17826(.Y(n_1122), .A0N(n_1120), .A1N(n_1118), .B0(n_1121));
  OR2X1 g17827(.Y(n_1121), .A(n_1120), .B(n_1118));
  ADDHX1 g17828(.CO(n_2870_danc), .S(n_2871_danc), .A(
    \dot_product_and_ReLU[4].product_terms[68][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[69][1] ));
  ADDHX1 g17829(.CO(n_1120), .S(n_1119), .A(
    \dot_product_and_ReLU[7].product_terms[109][1] ), .B(
    \dot_product_and_ReLU[16].product_terms[107][0] ));
  OR2X1 g17830(.Y(n_1527), .A(n_1508), .B(n_1116));
  NAND2X2 g17831(.Y(n_2981_danc), .A(n_1224), .B(n_1117));
  OAI21X1 g17832(.Y(n_1513), .A0(B[220]), .A1(n_1113), .B0(n_1227));
  OR2X1 g17833(.Y(n_1469), .A(n_1108), .B(n_1470));
  AND2X1 g17834(.Y(n_1534), .A(n_1518), .B(n_1242));
  NAND2BX1 g17835(.Y(n_1117), .AN(\dot_product_and_ReLU[1].product_terms[11][1] ),
     .B(n_2980_danc));
  OR2X1 g17836(.Y(n_1549), .A(n_1103), .B(n_1515));
  AOI21X1 g17837(.Y(n_1509), .A0(B[201]), .A1(B[200]), .B0(n_1112));
  NOR2BX1 g17838(.Y(n_1116), .AN(n_1507), .B(B[194]));
  OAI2BB1X1 g17839(.Y(n_1404), .A0N(
    \dot_product_and_ReLU[1].product_terms[132][1] ), .A1N(n_1101), .B0(n_1228));
  OR2X1 g17840(.Y(n_1414), .A(n_1109), .B(n_2950_danc));
  AOI21XL g17841(.Y(n_1118), .A0(\dot_product_and_ReLU[7].product_terms[111][0] ),
     .A1(n_1092), .B0(n_1111));
  AOI21X1 g17842(.Y(n_2818_danc), .A0(
    \dot_product_and_ReLU[3].product_terms[45][1] ), .A1(
    \dot_product_and_ReLU[2].product_terms[44][1] ), .B0(n_1104));
  AOI2BB1X1 g17843(.Y(n_1432), .A0N(
    \dot_product_and_ReLU[3].product_terms[54][0] ), .A1N(
    \dot_product_and_ReLU[1].product_terms[55][0] ), .B0(n_1433));
  AOI21X1 g17844(.Y(\level_1_sums[2][73] [0]), .A0(
    \dot_product_and_ReLU[1].product_terms[147][0] ), .A1(
    \dot_product_and_ReLU[4].product_terms[146][0] ), .B0(n_1115));
  AOI21X1 g17845(.Y(n_1523), .A0(B[231]), .A1(B[230]), .B0(n_1105));
  AOI2BB1X1 g17846(.Y(n_1541), .A0N(B[205]), .A1N(B[204]), .B0(n_1542));
  OR2X1 g17847(.Y(n_1396), .A(n_1110), .B(n_1397));
  AOI21X1 g17848(.Y(n_1390), .A0(\dot_product_and_ReLU[0].product_terms[150][0] ),
     .A1(\dot_product_and_ReLU[3].product_terms[151][0] ), .B0(n_1106));
  AOI21X1 g17849(.Y(n_1511), .A0(B[207]), .A1(B[206]), .B0(n_1114));
  AOI21X1 g17850(.Y(n_1516), .A0(B[238]), .A1(B[239]), .B0(n_1107));
  INVX1 g17852(.Y(n_1115), .A(\level_1_sums[2][73] [2]));
  INVX1 g17853(.Y(n_1512), .A(n_1114));
  INVX1 g17854(.Y(n_1514), .A(n_1113));
  INVX1 g17855(.Y(n_1510), .A(n_1112));
  NOR2BX1 g17856(.Y(n_1110), .AN(\dot_product_and_ReLU[9].product_terms[128][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[129][0] ));
  NOR2BX1 g17857(.Y(n_1109), .AN(\dot_product_and_ReLU[2].product_terms[37][1] ),
     .B(\dot_product_and_ReLU[8].product_terms[36][0] ));
  NOR2BX1 g17858(.Y(n_1108), .AN(\dot_product_and_ReLU[0].product_terms[5][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[4][0] ));
  NAND2BX1 g17859(.Y(n_1227), .AN(B[221]), .B(B[220]));
  NAND2X1 g17860(.Y(n_1242), .A(B[255]), .B(B[254]));
  OR2X1 g17861(.Y(\level_1_sums[2][73] [2]), .A(
    \dot_product_and_ReLU[1].product_terms[147][0] ), .B(
    \dot_product_and_ReLU[4].product_terms[146][0] ));
  OR2X1 g17862(.Y(n_2980_danc), .A(
    \dot_product_and_ReLU[7].product_terms[10][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[11][1] ));
  NAND2BX1 g17863(.Y(n_1228), .AN(
    \dot_product_and_ReLU[1].product_terms[132][1] ), .B(
    \dot_product_and_ReLU[4].product_terms[133][0] ));
  NOR2X1 g17864(.Y(n_1114), .A(B[207]), .B(B[206]));
  AND2X1 g17865(.Y(n_1542), .A(B[205]), .B(B[204]));
  NOR2BX1 g17866(.Y(n_1508), .AN(B[194]), .B(B[195]));
  NOR2X1 g17867(.Y(n_1113), .A(B[221]), .B(B[220]));
  NOR2X1 g17868(.Y(n_1112), .A(B[201]), .B(B[200]));
  NOR2X1 g17869(.Y(n_1111), .A(\dot_product_and_ReLU[7].product_terms[111][0] ),
     .B(n_1092));
  INVX1 g17870(.Y(n_1517), .A(n_1107));
  INVX1 g17871(.Y(n_1391), .A(n_1106));
  INVX1 g17872(.Y(n_1524), .A(n_1105));
  INVX1 g17873(.Y(n_1485), .A(n_1104));
  NOR2BX1 g17874(.Y(n_1103), .AN(B[233]), .B(B[232]));
  NAND2BX1 g17875(.Y(n_1224), .AN(\dot_product_and_ReLU[7].product_terms[10][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[11][1] ));
  NOR2X1 g17876(.Y(n_1107), .A(B[238]), .B(B[239]));
  NOR2BX1 g17877(.Y(n_1515), .AN(B[232]), .B(B[233]));
  OR2X1 g17878(.Y(n_1518), .A(B[255]), .B(B[254]));
  OR2X1 g17879(.Y(n_1507), .A(B[195]), .B(B[194]));
  NOR2X1 g17880(.Y(n_1106), .A(\dot_product_and_ReLU[3].product_terms[151][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[150][0] ));
  AND2X1 g17881(.Y(n_1433), .A(\dot_product_and_ReLU[1].product_terms[55][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[54][0] ));
  NOR2X1 g17882(.Y(n_1105), .A(B[231]), .B(B[230]));
  NOR2X1 g17883(.Y(n_1104), .A(\dot_product_and_ReLU[3].product_terms[45][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[44][1] ));
  NOR2BX1 g17884(.Y(n_1397), .AN(\dot_product_and_ReLU[2].product_terms[129][0] ),
     .B(\dot_product_and_ReLU[9].product_terms[128][1] ));
  NOR2BX1 g17885(.Y(n_2950_danc), .AN(
    \dot_product_and_ReLU[8].product_terms[36][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[37][1] ));
  NOR2X1 g17886(.Y(n_1102), .A(\dot_product_and_ReLU[14].product_terms[99][0] ),
     .B(\dot_product_and_ReLU[7].product_terms[103][0] ));
  NOR2BX1 g17887(.Y(n_1470), .AN(\dot_product_and_ReLU[2].product_terms[4][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[5][0] ));
  INVXL g17888(.Y(n_1101), .A(\dot_product_and_ReLU[4].product_terms[133][0] ));
  INVX1 g17889(.Y(n_1100), .A(\level_1_sums[4][37][1] ));
  INVX1 g17890(.Y(n_1099), .A(\dot_product_and_ReLU[4].product_terms[79][0] ));
  INVX1 g17891(.Y(n_1098), .A(\dot_product_and_ReLU[0].product_terms[106][0] ));
  INVX1 g17892(.Y(n_1097), .A(\dot_product_and_ReLU[5].product_terms[96][0] ));
  INVX1 g17893(.Y(n_1096), .A(\dot_product_and_ReLU[2].product_terms[95][0] ));
  INVX1 g17894(.Y(n_1095), .A(\dot_product_and_ReLU[0].product_terms[76][0] ));
  INVX1 g17895(.Y(n_1094), .A(\dot_product_and_ReLU[0].product_terms[105][0] ));
  INVX1 g17897(.Y(n_1093), .A(\dot_product_and_ReLU[12].product_terms[87][0] ));
  INVX1 g17898(.Y(n_1092), .A(\dot_product_and_ReLU[16].product_terms[102][2] ));
  INVX1 g17899(.Y(n_1091), .A(\dot_product_and_ReLU[4].product_terms[101][1] ));
  INVX1 g17900(.Y(n_1090), .A(\dot_product_and_ReLU[10].product_terms[80][0] ));
  INVX1 g17901(.Y(n_1089), .A(\dot_product_and_ReLU[5].product_terms[72][0] ));
  INVX1 g17903(.Y(n_1088), .A(\dot_product_and_ReLU[1].product_terms[77][0] ));
  CLKXOR2X1 g2(.Y(n_1087), .A(\dot_product_and_ReLU[14].product_terms[99][0] ),
     .B(\dot_product_and_ReLU[7].product_terms[103][0] ));
  OAI2BB1X1 g16637(.Y(n_1241), .A0N(
    \dot_product_and_ReLU[6].product_terms[43][0] ), .A1N(n_1083), .B0(n_1086));
  NAND2BX1 g16638(.Y(\level_2_sums[17][25][2] ), .AN(\level_2_sums[17][25][0] ),
     .B(n_1084));
  OAI2BB1X1 g16639(.Y(n_1240), .A0N(
    \dot_product_and_ReLU[0].product_terms[42][1] ), .A1N(n_1083), .B0(n_1086));
  CLKXOR2X1 g16640(.Y(\level_2_sums[17][29][1] ), .A(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .B(n_1411));
  OR2X1 g16641(.Y(n_1489), .A(n_1490), .B(n_1085));
  OR2X1 g16642(.Y(n_1086), .A(\dot_product_and_ReLU[0].product_terms[42][1] ),
     .B(n_1083));
  OAI21X1 g16643(.Y(n_2867_danc), .A0(
    \dot_product_and_ReLU[1].product_terms[77][0] ), .A1(n_1078), .B0(n_1221));
  OAI2BB1X1 g16644(.Y(\level_2_sums[17][29][2] ), .A0N(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .A1N(n_1081), .B0(n_1080));
  XNOR2X1 g16645(.Y(\level_2_sums[17][25][1] ), .A(
    \dot_product_and_ReLU[0].product_terms[100][0] ), .B(n_1223));
  NOR2BX1 g16646(.Y(n_1085), .AN(n_1491), .B(
    \dot_product_and_ReLU[19].product_terms[48][1] ));
  NAND2BX1 g16647(.Y(\level_1_sums[16][87] [1]), .AN(n_1454), .B(n_1218));
  NAND2BXL g16648(.Y(n_1084), .AN(n_1223), .B(
    \dot_product_and_ReLU[0].product_terms[100][0] ));
  OR2X1 g16649(.Y(n_2773_danc), .A(n_1494), .B(n_1082));
  AND2X1 g16650(.Y(\level_2_sums[17][25][0] ), .A(\level_2_sums[17][25][4] ), .B(
    n_1223));
  AOI21X1 g16651(.Y(n_1436), .A0(\dot_product_and_ReLU[3].product_terms[81][0] ),
     .A1(\dot_product_and_ReLU[10].product_terms[80][0] ), .B0(n_1079));
  OR2X1 g16652(.Y(n_1437), .A(n_1077), .B(n_1438));
  OAI2BB1X1 g16653(.Y(n_1479), .A0N(
    \dot_product_and_ReLU[19].product_terms[60][2] ), .A1N(n_1076), .B0(n_1220));
  AOI2BB1X1 g16654(.Y(n_1440), .A0N(
    \dot_product_and_ReLU[0].product_terms[130][0] ), .A1N(
    \dot_product_and_ReLU[14].product_terms[131][0] ), .B0(n_1441));
  NAND2X1 g16655(.Y(n_1411), .A(n_1081), .B(n_1080));
  XNOR2X1 g16656(.Y(n_1083), .A(\dot_product_and_ReLU[0].product_terms[41][0] ),
     .B(\dot_product_and_ReLU[6].product_terms[43][0] ));
  INVX1 g16657(.Y(n_1226), .A(n_1082));
  NOR2BX1 g16658(.Y(n_1082), .AN(\dot_product_and_ReLU[19].product_terms[59][1] ),
     .B(\dot_product_and_ReLU[7].product_terms[58][0] ));
  OR2X1 g16659(.Y(\level_2_sums[17][25][4] ), .A(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .B(
    \dot_product_and_ReLU[16].product_terms[102][2] ));
  NOR2BX1 g16660(.Y(n_1438), .AN(\dot_product_and_ReLU[0].product_terms[105][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[104] [1]));
  NAND2BX1 g16661(.Y(n_1081), .AN(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[119][0] ));
  NOR2BX1 g16662(.Y(n_1454), .AN(\dot_product_and_ReLU[2].product_terms[175][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[174][1] ));
  NOR2BX1 g16663(.Y(n_1490), .AN(\dot_product_and_ReLU[19].product_terms[48][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[49][0] ));
  OR2X1 g16664(.Y(n_1220), .A(\dot_product_and_ReLU[19].product_terms[60][2] ),
     .B(n_1076));
  OR2X1 g16665(.Y(n_1491), .A(\dot_product_and_ReLU[0].product_terms[49][0] ),
     .B(\dot_product_and_ReLU[19].product_terms[48][1] ));
  NAND2X1 g16666(.Y(n_1223), .A(\dot_product_and_ReLU[4].product_terms[101][1] ),
     .B(\dot_product_and_ReLU[16].product_terms[102][2] ));
  INVX1 g16667(.Y(n_2862_danc), .A(n_1079));
  INVX1 g16668(.Y(n_1078), .A(n_2866_danc));
  NOR2BX1 g16669(.Y(n_1077), .AN(\dot_product_and_ReLU[2].product_terms[104] [1]),
     .B(\dot_product_and_ReLU[0].product_terms[105][0] ));
  OR2X1 g16670(.Y(n_1405), .A(\dot_product_and_ReLU[8].product_terms[36][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[37][1] ));
  AND2XL g16671(.Y(n_1506), .A(B[255]), .B(n_1242));
  NOR2BX1 g16672(.Y(n_1494), .AN(\dot_product_and_ReLU[7].product_terms[58][0] ),
     .B(\dot_product_and_ReLU[19].product_terms[59][1] ));
  NAND2BX1 g16673(.Y(n_1080), .AN(
    \dot_product_and_ReLU[0].product_terms[119][0] ), .B(
    \dot_product_and_ReLU[4].product_terms[118][0] ));
  AND2X1 g16674(.Y(n_1441), .A(\dot_product_and_ReLU[14].product_terms[131][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[130][0] ));
  NOR2X1 g16675(.Y(n_1079), .A(\dot_product_and_ReLU[10].product_terms[80][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[81][0] ));
  NAND2BX1 g16676(.Y(n_1218), .AN(
    \dot_product_and_ReLU[2].product_terms[175][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[174][1] ));
  OR2X1 g16677(.Y(n_2866_danc), .A(
    \dot_product_and_ReLU[0].product_terms[76][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[77][0] ));
  NAND2BX1 g16678(.Y(n_1221), .AN(\dot_product_and_ReLU[0].product_terms[76][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[77][0] ));
  INVX1 g16679(.Y(n_1076), .A(\dot_product_and_ReLU[15].product_terms[61][1] ));
  INVX1 g17114(.Y(\level_4_sums[18][4] [8]), .A(n_1075));
  ADDFX1 g17115(.CO(n_1075), .S(\level_4_sums[18][4] [3]), .A(n_1053), .B(n_1071),
     .CI(n_1074));
  ADDFX1 g17116(.CO(n_1074), .S(\level_4_sums[18][4] [2]), .A(n_1069), .B(n_1072),
     .CI(n_1073));
  ADDFX1 g17117(.CO(n_1073), .S(\level_4_sums[18][4] [1]), .A(n_1065), .B(n_1070),
     .CI(n_1068));
  ADDFX1 g17118(.CO(n_1071), .S(n_1072), .A(n_1044), .B(n_1054), .CI(n_1064));
  ADDFX1 g17119(.CO(n_1069), .S(n_1070), .A(n_1051), .B(n_1060), .CI(n_1055));
  ADDFX1 g17120(.CO(n_1068), .S(\level_4_sums[18][4] [0]), .A(n_1046), .B(n_1061),
     .CI(n_1056));
  NAND2BX1 g17121(.Y(\level_3_sums[18][10] [1]), .AN(\level_3_sums[18][10] [2]),
     .B(n_1067));
  NOR2BX1 g17122(.Y(\level_3_sums[18][10] [2]), .AN(n_1062), .B(n_1066));
  NAND2BX1 g17123(.Y(n_1067), .AN(n_1062), .B(n_1066));
  ADDFX1 g17124(.CO(n_1066), .S(\level_3_sums[18][10] [0]), .A(
    \dot_product_and_ReLU[3].product_terms[86][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[81][0] ), .CI(n_1063));
  XNOR2X1 g17125(.Y(n_1234), .A(n_1399), .B(n_1052));
  ADDFX1 g17126(.CO(n_1064), .S(n_1065), .A(n_2870_danc), .B(n_1221), .CI(n_1047));
  INVX1 g17127(.Y(n_1063), .A(n_1059));
  INVX1 g17128(.Y(n_1061), .A(n_1058));
  INVX1 g17129(.Y(n_1060), .A(n_1057));
  ADDFX1 g17130(.CO(n_1062), .S(n_1059), .A(
    \dot_product_and_ReLU[3].product_terms[83][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[84][0] ), .CI(n_1038));
  ADDFX1 g17131(.CO(n_1057), .S(n_1058), .A(
    \dot_product_and_ReLU[4].product_terms[79][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[65][0] ), .CI(
    \dot_product_and_ReLU[16].product_terms[71][0] ));
  ADDFX1 g17132(.CO(n_1055), .S(n_1056), .A(
    \dot_product_and_ReLU[5].product_terms[72][0] ), .B(n_1037), .CI(
    n_2871_danc));
  OA21X1 g17133(.Y(n_1233), .A0(\dot_product_and_ReLU[1].product_terms[176][0] ),
     .A1(n_1050), .B0(n_1052));
  XNOR2X1 g17134(.Y(n_1054), .A(\dot_product_and_ReLU[0].product_terms[66][0] ),
     .B(n_1039));
  NOR2BX1 g17135(.Y(n_1053), .AN(n_1039), .B(
    \dot_product_and_ReLU[0].product_terms[66][0] ));
  CLKXOR2X1 g17136(.Y(n_1232), .A(
    \dot_product_and_ReLU[0].product_terms[179][0] ), .B(n_1399));
  NAND2X1 g17137(.Y(n_1052), .A(\dot_product_and_ReLU[1].product_terms[176][0] ),
     .B(n_1050));
  INVX1 g17138(.Y(n_1051), .A(n_1222));
  INVX1 g17139(.Y(n_1407), .A(n_1044));
  OAI2BB1X1 g17140(.Y(n_1050), .A0N(
    \dot_product_and_ReLU[0].product_terms[179][0] ), .A1N(
    \dot_product_and_ReLU[1].product_terms[176][0] ), .B0(n_1048));
  NAND2BX1 g17141(.Y(n_1448), .AN(n_1439), .B(n_1049));
  AOI21X1 g17142(.Y(n_2780_danc), .A0(
    \dot_product_and_ReLU[2].product_terms[40][0] ), .A1(
    \dot_product_and_ReLU[0].product_terms[41][0] ), .B0(n_1040));
  AOI21X1 g17143(.Y(\level_1_sums[12][86] [0]), .A0(
    \dot_product_and_ReLU[10].product_terms[172][1] ), .A1(
    \dot_product_and_ReLU[8].product_terms[173][1] ), .B0(n_1041));
  NAND2BXL g17144(.Y(n_1049), .AN(n_1388), .B(
    \dot_product_and_ReLU[0].product_terms[157][0] ));
  OA21X1 g17145(.Y(n_1492), .A0(\dot_product_and_ReLU[7].product_terms[57][2] ),
     .A1(\dot_product_and_ReLU[1].product_terms[56][1] ), .B0(n_1239));
  AOI21X1 g17146(.Y(n_1474), .A0(\dot_product_and_ReLU[2].product_terms[35][0] ),
     .A1(\dot_product_and_ReLU[2].product_terms[34][0] ), .B0(n_1045));
  OR2X1 g17147(.Y(n_1394), .A(n_1042), .B(n_1395));
  AO21X1 g17148(.Y(n_1222), .A0(\dot_product_and_ReLU[5].product_terms[72][0] ),
     .A1(\dot_product_and_ReLU[1].product_terms[73][0] ), .B0(n_1044));
  AOI2BB1X1 g17149(.Y(n_1428), .A0N(B[199]), .A1N(B[198]), .B0(n_1429));
  OR2X1 g17150(.Y(n_1382), .A(n_1043), .B(n_1383));
  OAI21XL g17151(.Y(n_1048), .A0(\dot_product_and_ReLU[0].product_terms[179][0] ),
     .A1(\dot_product_and_ReLU[1].product_terms[176][0] ), .B0(
    \dot_product_and_ReLU[0].product_terms[177][0] ));
  AOI2BB1X1 g17152(.Y(n_1408), .A0N(
    \dot_product_and_ReLU[0].product_terms[142][0] ), .A1N(
    \dot_product_and_ReLU[2].product_terms[143][0] ), .B0(n_1409));
  XNOR2X1 g17153(.Y(n_1047), .A(\dot_product_and_ReLU[7].product_terms[64][1] ),
     .B(\dot_product_and_ReLU[10].product_terms[78][1] ));
  OAI21X1 g17154(.Y(n_1046), .A0(\dot_product_and_ReLU[1].product_terms[77][0] ),
     .A1(n_1202), .B0(n_1221));
  CLKXOR2X1 g17155(.Y(n_1399), .A(
    \dot_product_and_ReLU[1].product_terms[176][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[177][0] ));
  INVX1 g17156(.Y(n_1475), .A(n_1045));
  NOR2BX1 g17157(.Y(n_1043), .AN(\dot_product_and_ReLU[1].product_terms[148][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[149][0] ));
  NOR2BX1 g17158(.Y(n_1042), .AN(\dot_product_and_ReLU[4].product_terms[97][0] ),
     .B(\dot_product_and_ReLU[5].product_terms[96][0] ));
  NOR2BX1 g17159(.Y(n_1395), .AN(\dot_product_and_ReLU[5].product_terms[96][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[97][0] ));
  NAND2X1 g17160(.Y(n_1239), .A(\dot_product_and_ReLU[7].product_terms[57][2] ),
     .B(\dot_product_and_ReLU[1].product_terms[56][1] ));
  NOR2X1 g17161(.Y(n_1045), .A(\dot_product_and_ReLU[2].product_terms[35][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[34][0] ));
  AND2X1 g17162(.Y(n_1388), .A(\dot_product_and_ReLU[17].product_terms[156][2] ),
     .B(\dot_product_and_ReLU[0].product_terms[157][0] ));
  AND2X1 g17163(.Y(n_1429), .A(B[198]), .B(B[199]));
  NOR2X1 g17164(.Y(n_1044), .A(\dot_product_and_ReLU[5].product_terms[72][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[73][0] ));
  INVX1 g17165(.Y(\level_1_sums[12][86] [1]), .A(n_1041));
  INVX1 g17166(.Y(n_2779_danc), .A(n_1040));
  NOR2X1 g17167(.Y(n_2817_danc), .A(n_1201), .B(n_1200));
  AND2XL g17168(.Y(n_1535), .A(B[254]), .B(n_1242));
  NOR2X1 g17169(.Y(n_1041), .A(\dot_product_and_ReLU[10].product_terms[172][1] ),
     .B(\dot_product_and_ReLU[8].product_terms[173][1] ));
  NOR2X1 g17170(.Y(n_1040), .A(\dot_product_and_ReLU[2].product_terms[40][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[41][0] ));
  NOR2BX1 g17171(.Y(n_1383), .AN(\dot_product_and_ReLU[1].product_terms[149][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[148][0] ));
  AND2X1 g17172(.Y(n_1409), .A(\dot_product_and_ReLU[0].product_terms[142][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[143][0] ));
  NOR2BX1 g17173(.Y(n_1439), .AN(
    \dot_product_and_ReLU[17].product_terms[156][2] ), .B(
    \dot_product_and_ReLU[0].product_terms[157][0] ));
  NOR2BX1 g17174(.Y(n_1039), .AN(\dot_product_and_ReLU[10].product_terms[78][1] ),
     .B(\dot_product_and_ReLU[7].product_terms[64][1] ));
  INVX1 g17175(.Y(n_1038), .A(\dot_product_and_ReLU[10].product_terms[80][0] ));
  INVX1 g17176(.Y(n_1037), .A(\dot_product_and_ReLU[5].product_terms[75][0] ));
  AOI21X1 g17904(.Y(n_2976_danc), .A0(
    \dot_product_and_ReLU[0].product_terms[27][0] ), .A1(
    \dot_product_and_ReLU[19].product_terms[26][2] ), .B0(n_1036));
  AND2X1 g17905(.Y(n_2788_danc), .A(n_1482), .B(n_1034));
  AOI21X1 g17906(.Y(n_2823_danc), .A0(
    \dot_product_and_ReLU[0].product_terms[42][1] ), .A1(
    \dot_product_and_ReLU[6].product_terms[43][0] ), .B0(n_1033));
  OR2X1 g17907(.Y(n_1392), .A(n_1035), .B(n_1393));
  INVX1 g17908(.Y(n_2996_danc), .A(n_1036));
  NOR2BX1 g17909(.Y(n_1035), .AN(\dot_product_and_ReLU[0].product_terms[159][1] ),
     .B(\dot_product_and_ReLU[1].product_terms[158][0] ));
  NAND2XL g17910(.Y(n_1034), .A(\dot_product_and_ReLU[0].product_terms[17][1] ),
     .B(\dot_product_and_ReLU[7].product_terms[16][0] ));
  OR2X1 g17911(.Y(n_1381), .A(\dot_product_and_ReLU[0].product_terms[130][0] ),
     .B(\dot_product_and_ReLU[14].product_terms[131][0] ));
  NOR2BX1 g17912(.Y(n_1393), .AN(\dot_product_and_ReLU[1].product_terms[158][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[159][1] ));
  NOR2X1 g16363(.Y(n_1036), .A(\dot_product_and_ReLU[0].product_terms[27][0] ),
     .B(\dot_product_and_ReLU[19].product_terms[26][2] ));
  INVX1 g16364(.Y(n_2822_danc), .A(n_1033));
  NAND2X1 g16365(.Y(n_1378), .A(n_1203), .B(n_1198));
  NAND2X1 g16366(.Y(n_1400), .A(n_1193), .B(n_1207));
  NOR2X1 g16367(.Y(n_2929_danc), .A(n_1194), .B(n_1199));
  NOR2X1 g16368(.Y(n_1033), .A(\dot_product_and_ReLU[0].product_terms[42][1] ),
     .B(\dot_product_and_ReLU[6].product_terms[43][0] ));
  OR2X1 g16369(.Y(n_1482), .A(\dot_product_and_ReLU[0].product_terms[17][1] ),
     .B(\dot_product_and_ReLU[7].product_terms[16][0] ));
  INVX1 g16370(.Y(\level_1_sums[16][87] [2]), .A(n_1218));
  OA21X1 g17106(.Y(\level_4_sums[11][5] [4]), .A0(n_1030), .A1(n_1032), .B0(
    \level_4_sums[11][5] [8]));
  NAND2X1 g17107(.Y(\level_4_sums[11][5] [8]), .A(n_1030), .B(n_1032));
  ADDFX1 g17108(.CO(n_1032), .S(\level_4_sums[11][5] [3]), .A(n_1008), .B(n_1029),
     .CI(n_1031));
  ADDFX1 g17109(.CO(n_1031), .S(\level_4_sums[11][5] [2]), .A(n_1009), .B(n_1028),
     .CI(n_1027));
  ADDFX1 g17110(.CO(n_1030), .S(n_1029), .A(n_1003), .B(n_1019), .CI(n_1026));
  ADDFX1 g17111(.CO(n_1028), .S(\level_4_sums[11][5] [1]), .A(n_1017), .B(n_1023),
     .CI(n_1025));
  ADDFX1 g17112(.CO(n_1026), .S(n_1027), .A(n_1021), .B(n_1020), .CI(n_1024));
  ADDFX1 g17113(.CO(n_1024), .S(n_1025), .A(
    \dot_product_and_ReLU[0].product_terms[88][1] ), .B(n_1004), .CI(n_1022));
  ADDFX1 g17913(.CO(n_1023), .S(\level_4_sums[11][5] [0]), .A(
    \dot_product_and_ReLU[0].product_terms[88][1] ), .B(n_1016), .CI(n_1018));
  ADDFX1 g17914(.CO(n_1021), .S(n_1022), .A(
    \dot_product_and_ReLU[3].product_terms[81][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[85][0] ), .CI(n_1015));
  ADDFX1 g17915(.CO(n_1019), .S(n_1020), .A(n_999), .B(n_996), .CI(n_1010));
  ADDFX1 g17916(.CO(n_1017), .S(n_1018), .A(n_997), .B(
    \dot_product_and_ReLU[0].product_terms[94][1] ), .CI(n_1011));
  ADDFX1 g17917(.CO(n_1015), .S(n_1016), .A(
    \dot_product_and_ReLU[2].product_terms[91][1] ), .B(n_1000), .CI(n_998));
  AO21X1 g17918(.Y(n_1402), .A0(n_1228), .A1(n_1014), .B0(n_1403));
  NOR2X1 g17919(.Y(n_1403), .A(n_1228), .B(n_1014));
  ADDHX1 g17920(.CO(n_1014), .S(n_1401), .A(
    \dot_product_and_ReLU[2].product_terms[134][1] ), .B(n_1404));
  OR2X1 g17921(.Y(n_2603_danc), .A(n_2602_danc), .B(n_1013));
  OR2X1 g17922(.Y(n_1384), .A(n_1386), .B(n_1012));
  OR2X1 g17923(.Y(n_1553), .A(n_1007), .B(n_1531));
  NOR2BX1 g17924(.Y(n_1013), .AN(n_1487), .B(B[223]));
  NOR2BX1 g17925(.Y(n_1012), .AN(n_1385), .B(
    \dot_product_and_ReLU[4].product_terms[166][0] ));
  OR2X1 g17926(.Y(n_1495), .A(n_1006), .B(n_1496));
  OR2X1 g17927(.Y(n_1426), .A(n_1002), .B(n_1427));
  OR2X1 g17928(.Y(n_2926_danc), .A(n_1001), .B(n_2925_danc));
  OR2X1 g17929(.Y(n_1529), .A(n_1005), .B(n_1530));
  OA21X1 g17930(.Y(n_1547), .A0(B[225]), .A1(B[224]), .B0(n_1246));
  OAI2BB1X1 g17931(.Y(n_1011), .A0N(
    \dot_product_and_ReLU[10].product_terms[80][0] ), .A1N(
    \dot_product_and_ReLU[3].product_terms[84][0] ), .B0(n_1004));
  OAI21X1 g17932(.Y(n_1010), .A0(\dot_product_and_ReLU[8].product_terms[92][1] ),
     .A1(\dot_product_and_ReLU[2].product_terms[91][1] ), .B0(n_1003));
  AOI21X1 g17933(.Y(n_1009), .A0(\dot_product_and_ReLU[13].product_terms[89][0] ),
     .A1(\dot_product_and_ReLU[0].product_terms[88][1] ), .B0(n_1008));
  AND2X1 g17934(.Y(n_1528), .A(B[195]), .B(B[194]));
  NOR2BX1 g17935(.Y(n_1007), .AN(B[242]), .B(B[243]));
  OR2XL g17936(.Y(n_1471), .A(\dot_product_and_ReLU[0].product_terms[5][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[4][0] ));
  NOR2BX1 g17937(.Y(n_1006), .AN(B[247]), .B(B[246]));
  NOR2BX1 g17938(.Y(n_1005), .AN(B[211]), .B(B[210]));
  NOR2BX1 g17939(.Y(n_1386), .AN(\dot_product_and_ReLU[4].product_terms[166][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[167][0] ));
  NOR2BX1 g17940(.Y(n_1531), .AN(B[243]), .B(B[242]));
  NOR2BX1 g17941(.Y(n_1530), .AN(B[210]), .B(B[211]));
  NAND2X1 g17942(.Y(n_1246), .A(B[225]), .B(B[224]));
  NOR2X1 g17943(.Y(n_1008), .A(\dot_product_and_ReLU[13].product_terms[89][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[88][1] ));
  NOR2BX1 g17944(.Y(n_1002), .AN(\dot_product_and_ReLU[1].product_terms[108][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[110][0] ));
  NOR2BX1 g17945(.Y(n_1001), .AN(\dot_product_and_ReLU[3].product_terms[120][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[121][1] ));
  OR2X1 g17946(.Y(n_1487), .A(B[222]), .B(B[223]));
  NOR2BX1 g17947(.Y(n_1496), .AN(B[246]), .B(B[247]));
  NOR2BX1 g17948(.Y(n_1427), .AN(\dot_product_and_ReLU[3].product_terms[110][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[108][0] ));
  NOR2BX1 g17949(.Y(n_2602_danc), .AN(B[223]), .B(B[222]));
  OR2X1 g17950(.Y(n_1385), .A(\dot_product_and_ReLU[0].product_terms[167][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[166][0] ));
  NOR2BX1 g17951(.Y(n_2925_danc), .AN(
    \dot_product_and_ReLU[2].product_terms[121][1] ), .B(
    \dot_product_and_ReLU[3].product_terms[120][1] ));
  OR2X1 g17952(.Y(n_1004), .A(\dot_product_and_ReLU[10].product_terms[80][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[84][0] ));
  NAND2X1 g17953(.Y(n_1003), .A(\dot_product_and_ReLU[2].product_terms[91][1] ),
     .B(\dot_product_and_ReLU[8].product_terms[92][1] ));
  INVX1 g17954(.Y(n_1497), .A(n_1227));
  INVX1 g17955(.Y(n_1000), .A(\dot_product_and_ReLU[3].product_terms[83][0] ));
  INVX1 g17956(.Y(n_999), .A(\dot_product_and_ReLU[0].product_terms[94][1] ));
  INVX1 g17957(.Y(n_998), .A(\dot_product_and_ReLU[0].product_terms[90][0] ));
  INVX1 g17958(.Y(n_997), .A(\dot_product_and_ReLU[3].product_terms[86][0] ));
  INVX1 g17959(.Y(n_996), .A(\dot_product_and_ReLU[1].product_terms[85][0] ));
  OR2X1 g16443(.Y(\level_1_sums[8][55] [0]), .A(\level_1_sums[8][55] [1]), .B(
    n_995));
  OAI21X1 g16444(.Y(n_1452), .A0(\dot_product_and_ReLU[1].product_terms[170][0] ),
     .A1(n_992), .B0(n_1225));
  NOR2BX1 g16445(.Y(n_995), .AN(\level_1_sums[8][55] [4]), .B(
    \dot_product_and_ReLU[3].product_terms[110][0] ));
  OR2X1 g16446(.Y(n_1498), .A(n_993), .B(n_1499));
  AOI2BB1X1 g16447(.Y(n_1539), .A0N(B[197]), .A1N(B[196]), .B0(n_1540));
  AOI2BB1X1 g16448(.Y(n_1430), .A0N(
    \dot_product_and_ReLU[6].product_terms[9][0] ), .A1N(
    \dot_product_and_ReLU[0].product_terms[8][0] ), .B0(n_1431));
  OR2X1 g16449(.Y(n_1463), .A(n_994), .B(n_1464));
  NOR2BX1 g16450(.Y(n_994), .AN(\dot_product_and_ReLU[4].product_terms[24][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[25][0] ));
  NOR2BX1 g16451(.Y(n_993), .AN(B[236]), .B(B[237]));
  NOR2BX1 g16452(.Y(n_1499), .AN(B[237]), .B(B[236]));
  AND2X1 g16453(.Y(n_1540), .A(B[197]), .B(B[196]));
  NOR2BX1 g16454(.Y(\level_1_sums[8][55] [1]), .AN(
    \dot_product_and_ReLU[3].product_terms[110][0] ), .B(
    \dot_product_and_ReLU[7].product_terms[111][0] ));
  OR2X1 g16455(.Y(\level_1_sums[8][55] [4]), .A(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[110][0] ));
  INVX1 g16456(.Y(n_1398), .A(n_992));
  AND2X1 g16457(.Y(n_2667_danc), .A(n_1246), .B(B[225]));
  OR2X1 g16458(.Y(n_2772_danc), .A(
    \dot_product_and_ReLU[19].product_terms[59][1] ), .B(
    \dot_product_and_ReLU[7].product_terms[58][0] ));
  NAND2BX1 g16459(.Y(n_1225), .AN(
    \dot_product_and_ReLU[1].product_terms[171][1] ), .B(
    \dot_product_and_ReLU[1].product_terms[170][0] ));
  AND2X1 g16460(.Y(n_1431), .A(\dot_product_and_ReLU[0].product_terms[8][0] ),
     .B(\dot_product_and_ReLU[6].product_terms[9][0] ));
  NOR2BX1 g16461(.Y(n_1464), .AN(\dot_product_and_ReLU[3].product_terms[25][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[24][0] ));
  NOR2X1 g16462(.Y(n_992), .A(\dot_product_and_ReLU[1].product_terms[171][1] ),
     .B(\dot_product_and_ReLU[1].product_terms[170][0] ));
  AOI2BB1X1 g16388(.Y(\level_1_sums[7][92] [0]), .A0N(
    \dot_product_and_ReLU[3].product_terms[184][1] ), .A1N(
    \dot_product_and_ReLU[5].product_terms[185][0] ), .B0(
    \level_1_sums[7][92] [1]));
  AOI21X1 g16389(.Y(n_2757_danc), .A0(
    \dot_product_and_ReLU[4].product_terms[1][0] ), .A1(
    \dot_product_and_ReLU[0].product_terms[0][0] ), .B0(n_990));
  OR2X1 g16390(.Y(n_1443), .A(n_991), .B(n_2826_danc));
  AOI21X1 g16391(.Y(\level_1_sums[3][46] [0]), .A0(
    \dot_product_and_ReLU[0].product_terms[93][0] ), .A1(
    \dot_product_and_ReLU[8].product_terms[92][1] ), .B0(n_989));
  OA21X1 g16392(.Y(n_1536), .A0(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .A1(\dot_product_and_ReLU[0].product_terms[179][0] ), .B0(n_1243));
  OR2XL g16393(.Y(n_1389), .A(\dot_product_and_ReLU[0].product_terms[142][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[143][0] ));
  AND2X1 g16394(.Y(n_2631_danc), .A(B[246]), .B(B[247]));
  NOR2BX1 g16395(.Y(n_991), .AN(\dot_product_and_ReLU[0].product_terms[23][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[22][0] ));
  OR2X1 g16396(.Y(n_1245), .A(B[228]), .B(B[229]));
  NOR2BX1 g16397(.Y(n_2826_danc), .AN(
    \dot_product_and_ReLU[0].product_terms[22][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[23][0] ));
  AND2X1 g16398(.Y(\level_1_sums[7][92] [1]), .A(
    \dot_product_and_ReLU[5].product_terms[185][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[184][1] ));
  INVX1 g16399(.Y(n_1461), .A(n_990));
  INVX1 g16400(.Y(\level_1_sums[3][46] [4]), .A(n_989));
  AND2XL g16401(.Y(n_1244), .A(B[228]), .B(B[229]));
  OR2X1 g16402(.Y(n_1504), .A(B[211]), .B(B[210]));
  NOR2X1 g16403(.Y(n_1387), .A(n_1205), .B(n_1191));
  NAND2XL g16404(.Y(n_1243), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[179][0] ));
  NOR2X1 g16405(.Y(n_990), .A(\dot_product_and_ReLU[4].product_terms[1][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[0][0] ));
  NOR2X1 g16406(.Y(n_989), .A(\dot_product_and_ReLU[0].product_terms[93][0] ),
     .B(\dot_product_and_ReLU[8].product_terms[92][1] ));
  INVX1 g16407(.Y(n_1442), .A(n_1224));
  OR2X1 g17960(.Y(n_1500), .A(n_1501), .B(n_988));
  AOI21X1 g16463(.Y(n_1483), .A0(\dot_product_and_ReLU[0].product_terms[29][0] ),
     .A1(\dot_product_and_ReLU[0].product_terms[28][0] ), .B0(n_984));
  OR2X1 g16464(.Y(n_1480), .A(n_985), .B(n_1481));
  NOR2BX1 g16465(.Y(n_988), .AN(n_1502), .B(B[240]));
  AOI21X1 g16466(.Y(n_1543), .A0(B[217]), .A1(B[216]), .B0(n_987));
  AOI21X1 g16467(.Y(n_1525), .A0(B[250]), .A1(B[251]), .B0(n_986));
  OR2X1 g16468(.Y(n_1532), .A(n_982), .B(n_1533));
  OR2X1 g16469(.Y(n_1444), .A(n_981), .B(n_1445));
  AOI21X1 g16470(.Y(n_1446), .A0(\dot_product_and_ReLU[2].product_terms[113][1] ),
     .A1(\dot_product_and_ReLU[17].product_terms[112][2] ), .B0(n_983));
  INVX1 g16471(.Y(n_1544), .A(n_987));
  INVX1 g16472(.Y(n_1503), .A(n_986));
  NOR2BX1 g16473(.Y(n_985), .AN(\dot_product_and_ReLU[0].product_terms[6][2] ),
     .B(\dot_product_and_ReLU[7].product_terms[7][0] ));
  OR2X1 g16474(.Y(n_1502), .A(B[241]), .B(B[240]));
  NOR2X1 g16475(.Y(n_987), .A(B[217]), .B(B[216]));
  NOR2BX1 g16476(.Y(n_1533), .AN(B[244]), .B(B[245]));
  NOR2BX1 g16477(.Y(n_1445), .AN(\dot_product_and_ReLU[7].product_terms[109][1] ),
     .B(\dot_product_and_ReLU[1].product_terms[108][0] ));
  NOR2XL g16478(.Y(n_986), .A(B[250]), .B(B[251]));
  INVX1 g16479(.Y(n_1484), .A(n_984));
  INVX1 g16480(.Y(n_1447), .A(n_983));
  NAND2X1 g16481(.Y(n_1554), .A(n_1210), .B(n_1211));
  NOR2BX1 g16482(.Y(n_982), .AN(B[245]), .B(B[244]));
  NOR2BX1 g16483(.Y(n_981), .AN(\dot_product_and_ReLU[1].product_terms[108][0] ),
     .B(\dot_product_and_ReLU[7].product_terms[109][1] ));
  NOR2X1 g16484(.Y(n_984), .A(\dot_product_and_ReLU[0].product_terms[29][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[28][0] ));
  NOR2BX1 g16485(.Y(n_1481), .AN(\dot_product_and_ReLU[7].product_terms[7][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[6][2] ));
  NOR2X1 g16486(.Y(n_983), .A(\dot_product_and_ReLU[2].product_terms[113][1] ),
     .B(\dot_product_and_ReLU[17].product_terms[112][2] ));
  NOR2BX1 g16487(.Y(n_1501), .AN(B[240]), .B(B[241]));
  DFFRHQX1 \out_reg_reg[19][4] (.Q(out[175]), .D(n_976), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][6] (.Q(out[177]), .D(n_973), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][7] (.Q(out[178]), .D(n_979), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][0] (.Q(out[171]), .D(n_978), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][2] (.Q(out[173]), .D(n_975), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][5] (.Q(out[176]), .D(n_980), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][3] (.Q(out[174]), .D(n_977), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[19][1] (.Q(out[172]), .D(n_974), .RN(rst_n), .CK(clk));
  NOR2X1 g16521(.Y(n_980), .A(n_967), .B(n_972));
  NOR2X1 g16522(.Y(n_979), .A(n_970), .B(n_972));
  NOR2X1 g16523(.Y(n_978), .A(\level_8_sums[19] [0]), .B(n_972));
  NOR2X1 g16524(.Y(n_977), .A(n_962), .B(n_972));
  NOR2X1 g16525(.Y(n_976), .A(n_964), .B(n_972));
  NOR2X1 g16526(.Y(n_975), .A(n_959), .B(n_972));
  NOR2X1 g16527(.Y(n_974), .A(n_957), .B(n_972));
  NOR2X1 g16528(.Y(n_973), .A(n_969), .B(n_972));
  XNOR2X1 g16529(.Y(n_972), .A(\level_8_sums[19] [9]), .B(n_971));
  NAND3BXL g16530(.Y(n_971), .AN(n_968), .B(\level_8_sums[19] [7]), .C(
    \level_8_sums[19] [8]));
  XOR2XL g16531(.Y(n_970), .A(n_968), .B(\level_8_sums[19] [7]));
  XNOR2X1 g16532(.Y(n_969), .A(\level_8_sums[19] [6]), .B(n_966));
  NAND2X1 g16533(.Y(n_968), .A(\level_8_sums[19] [6]), .B(n_966));
  AOI21X1 g16534(.Y(n_967), .A0(n_963), .A1(\level_8_sums[19] [5]), .B0(n_965));
  INVX1 g16535(.Y(n_966), .A(n_965));
  NOR2X1 g16536(.Y(n_965), .A(n_963), .B(\level_8_sums[19] [5]));
  XNOR2X1 g16537(.Y(n_964), .A(\level_8_sums[19] [4]), .B(n_961));
  AND2XL g16538(.Y(n_963), .A(\level_8_sums[19] [4]), .B(n_961));
  AOI21X1 g16539(.Y(n_962), .A0(n_958), .A1(\level_8_sums[19] [3]), .B0(n_960));
  INVX1 g16540(.Y(n_961), .A(n_960));
  NOR2XL g16541(.Y(n_960), .A(n_958), .B(\level_8_sums[19] [3]));
  XNOR2X1 g16542(.Y(n_959), .A(n_956), .B(\level_8_sums[19] [2]));
  AND2XL g16543(.Y(n_958), .A(n_956), .B(\level_8_sums[19] [2]));
  XNOR2X1 g16544(.Y(n_957), .A(\level_8_sums[19] [0]), .B(\level_8_sums[19] [1]));
  AND2XL g16545(.Y(n_956), .A(\level_8_sums[19] [0]), .B(\level_8_sums[19] [1]));
  AO21XL g17961(.Y(\level_4_sums[16][10][3] ), .A0(n_946), .A1(n_955), .B0(
    \level_4_sums[16][10][7] ));
  NOR2X1 g17962(.Y(\level_4_sums[16][10][7] ), .A(n_946), .B(n_955));
  XNOR2X1 g17963(.Y(\level_3_sums[16][15] [3]), .A(n_951), .B(n_954));
  ADDFX1 g17964(.CO(n_955), .S(\level_4_sums[16][10][2] ), .A(n_947), .B(n_944),
     .CI(n_953));
  ADDFX1 g17965(.CO(n_954), .S(\level_3_sums[16][15] [2]), .A(n_941), .B(n_950),
     .CI(n_952));
  ADDFX1 g17966(.CO(n_953), .S(\level_4_sums[16][10][1] ), .A(n_923), .B(n_927),
     .CI(n_945));
  ADDFX1 g17177(.CO(n_952), .S(\level_3_sums[16][15] [1]), .A(n_932), .B(n_942),
     .CI(n_948));
  XNOR2X1 g17178(.Y(n_951), .A(n_949), .B(n_943));
  ADDFX1 g17179(.CO(n_949), .S(n_950), .A(
    \dot_product_and_ReLU[3].product_terms[123][1] ), .B(n_931), .CI(n_936));
  ADDFX1 g17180(.CO(n_948), .S(\level_3_sums[16][15] [0]), .A(
    \dot_product_and_ReLU[3].product_terms[123][1] ), .B(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .CI(n_929));
  XNOR2X1 g17181(.Y(n_947), .A(n_937), .B(n_940));
  AOI221X1 g17182(.Y(n_946), .A0(n_935), .A1(n_918), .B0(n_937), .B1(n_938), .C0(
    n_933));
  ADDFX1 g17183(.CO(n_944), .S(n_945), .A(
    \dot_product_and_ReLU[0].product_terms[167][0] ), .B(n_922), .CI(n_911));
  XNOR2X1 g17184(.Y(n_943), .A(n_939), .B(n_936));
  ADDFX1 g17185(.CO(n_941), .S(n_942), .A(
    \dot_product_and_ReLU[4].product_terms[126][1] ), .B(
    \dot_product_and_ReLU[3].product_terms[123][1] ), .CI(n_928));
  OR2X1 g17186(.Y(n_1478), .A(n_919), .B(n_926));
  MXI2XL g17187(.Y(n_940), .A(n_934), .B(n_935), .S0(n_918));
  XNOR2X1 g17188(.Y(n_939), .A(\dot_product_and_ReLU[3].product_terms[123][1] ),
     .B(n_930));
  OR2XL g17189(.Y(n_938), .A(n_935), .B(n_918));
  AO21X1 g17190(.Y(n_1477), .A0(n_921), .A1(n_925), .B0(n_926));
  AOI21X1 g17191(.Y(n_937), .A0(n_1218), .A1(n_924), .B0(n_933));
  INVX1 g17192(.Y(n_935), .A(n_934));
  ADDFX1 g17193(.CO(n_931), .S(n_932), .A(
    \dot_product_and_ReLU[17].product_terms[124][0] ), .B(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .CI(n_917));
  ADDFX1 g17194(.CO(n_930), .S(n_936), .A(
    \dot_product_and_ReLU[4].product_terms[126][1] ), .B(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .CI(n_917));
  ADDFX1 g17195(.CO(n_928), .S(n_929), .A(
    \dot_product_and_ReLU[17].product_terms[124][0] ), .B(
    \dot_product_and_ReLU[4].product_terms[125][1] ), .CI(n_2926_danc));
  ADDFX1 g17196(.CO(n_934), .S(n_927), .A(
    \dot_product_and_ReLU[1].product_terms[170][0] ), .B(
    \dot_product_and_ReLU[5].product_terms[160][1] ), .CI(
    \level_1_sums[1][81][0] ));
  NOR2X1 g17197(.Y(n_933), .A(n_1218), .B(n_924));
  NOR2XL g17198(.Y(n_926), .A(n_921), .B(n_925));
  ADDFX1 g17199(.CO(n_923), .S(\level_4_sums[16][10][0] ), .A(
    \dot_product_and_ReLU[2].product_terms[174][1] ), .B(n_913), .CI(n_916));
  ADDFX1 g17200(.CO(n_925), .S(n_1476), .A(
    \dot_product_and_ReLU[0].product_terms[63][1] ), .B(
    \dot_product_and_ReLU[1].product_terms[62][0] ), .CI(n_1479));
  ADDFX1 g17201(.CO(n_924), .S(n_922), .A(
    \dot_product_and_ReLU[3].product_terms[164][0] ), .B(n_912), .CI(n_914));
  AOI21X1 g17202(.Y(n_1379), .A0(\dot_product_and_ReLU[0].product_terms[141][0] ),
     .A1(\dot_product_and_ReLU[17].product_terms[140] [0]), .B0(n_920));
  AO21XL g17203(.Y(n_921), .A0(n_915), .A1(n_1220), .B0(n_919));
  INVX1 g17205(.Y(n_1380), .A(n_920));
  OR2XL g17206(.Y(n_1415), .A(\dot_product_and_ReLU[3].product_terms[184][1] ),
     .B(\dot_product_and_ReLU[5].product_terms[185][0] ));
  NOR2X1 g17207(.Y(n_920), .A(\dot_product_and_ReLU[17].product_terms[140] [0]),
     .B(\dot_product_and_ReLU[0].product_terms[141][0] ));
  NOR2X1 g17208(.Y(n_919), .A(n_915), .B(n_1220));
  INVX1 g17210(.Y(n_1219), .A(n_917));
  NAND2X1 g17211(.Y(n_1462), .A(n_1196), .B(n_1197));
  NOR2X1 g17212(.Y(n_2975_danc), .A(
    \dot_product_and_ReLU[0].product_terms[27][0] ), .B(n_1195));
  NOR2X1 g17213(.Y(n_918), .A(\dot_product_and_ReLU[3].product_terms[168][0] ),
     .B(\level_1_sums[16][87] [1]));
  NOR2BX1 g17214(.Y(n_917), .AN(\dot_product_and_ReLU[3].product_terms[120][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[121][1] ));
  INVX1 g17215(.Y(n_916), .A(\dot_product_and_ReLU[2].product_terms[165][0] ));
  INVX1 g17216(.Y(n_915), .A(\dot_product_and_ReLU[1].product_terms[62][0] ));
  INVX1 g17217(.Y(n_914), .A(\dot_product_and_ReLU[4].product_terms[166][0] ));
  INVX1 g17218(.Y(n_913), .A(\dot_product_and_ReLU[1].product_terms[171][1] ));
  INVX1 g17219(.Y(n_912), .A(\dot_product_and_ReLU[8].product_terms[173][1] ));
  AO21XL g17967(.Y(n_911), .A0(\dot_product_and_ReLU[3].product_terms[168][0] ),
     .A1(\level_1_sums[16][87] [1]), .B0(n_918));
  AOI2BB1X1 g17968(.Y(n_2928_danc), .A0N(
    \dot_product_and_ReLU[2].product_terms[95][0] ), .A1N(
    \dot_product_and_ReLU[0].product_terms[94][1] ), .B0(n_2927_danc));
  AOI2BB1X1 g17969(.Y(n_1466), .A0N(
    \dot_product_and_ReLU[4].product_terms[15][0] ), .A1N(
    \dot_product_and_ReLU[6].product_terms[14][1] ), .B0(n_1467));
  OR2X1 g17970(.Y(n_1434), .A(n_910), .B(n_2864_danc));
  NOR2BX1 g17971(.Y(n_2864_danc), .AN(B[203]), .B(B[202]));
  AND2X1 g17972(.Y(n_1467), .A(\dot_product_and_ReLU[4].product_terms[15][0] ),
     .B(\dot_product_and_ReLU[6].product_terms[14][1] ));
  AND2X1 g17973(.Y(n_2927_danc), .A(
    \dot_product_and_ReLU[2].product_terms[95][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[94][1] ));
  AND2X1 g16371(.Y(n_1413), .A(\dot_product_and_ReLU[0].product_terms[42][1] ),
     .B(\dot_product_and_ReLU[6].product_terms[43][0] ));
  NOR2BX1 g16372(.Y(n_910), .AN(B[202]), .B(B[203]));
  AND2X1 g16373(.Y(n_1526), .A(B[251]), .B(B[250]));
  INVX1 g16374(.Y(n_3001_danc), .A(n_1219));
  AOI21X1 g17974(.Y(\level_4_sums[12][8] [8]), .A0(n_825), .A1(n_879), .B0(n_909));
  ADDFX1 g17975(.CO(n_909), .S(\level_4_sums[12][8] [3]), .A(n_887), .B(n_898),
     .CI(n_907));
  INVX1 g17976(.Y(\level_4_sums[12][11][6] ), .A(n_908));
  ADDFX1 g17977(.CO(n_908), .S(\level_4_sums[12][11][3] ), .A(n_855), .B(n_900),
     .CI(n_906));
  AO21XL g17978(.Y(\level_4_sums[12][6] [3]), .A0(n_884), .A1(n_905), .B0(
    \level_4_sums[12][6] [8]));
  ADDFX1 g17979(.CO(n_907), .S(\level_4_sums[12][8] [2]), .A(n_889), .B(n_899),
     .CI(n_903));
  ADDFX1 g17980(.CO(n_906), .S(\level_4_sums[12][11][2] ), .A(n_896), .B(n_901),
     .CI(n_904));
  NOR2X1 g17981(.Y(\level_4_sums[12][6] [8]), .A(n_884), .B(n_905));
  ADDFX1 g17982(.CO(n_905), .S(\level_4_sums[12][6] [2]), .A(n_893), .B(n_881),
     .CI(n_902));
  ADDFX1 g17983(.CO(n_904), .S(\level_4_sums[12][11][1] ), .A(n_886), .B(n_895),
     .CI(n_897));
  ADDFX1 g17984(.CO(n_903), .S(\level_4_sums[12][8] [1]), .A(n_850), .B(n_880),
     .CI(n_890));
  ADDFX1 g17985(.CO(n_902), .S(\level_4_sums[12][6] [1]), .A(n_870), .B(n_894),
     .CI(n_888));
  ADDFX1 g17986(.CO(n_900), .S(n_901), .A(n_875), .B(n_856), .CI(n_885));
  ADDFX1 g17987(.CO(n_898), .S(n_899), .A(n_847), .B(n_865), .CI(n_877));
  ADDFX1 g17851(.CO(n_896), .S(n_897), .A(n_832), .B(n_867), .CI(n_876));
  INVX1 g17988(.Y(\level_4_sums[12][11][0] ), .A(n_892));
  INVX1 g17989(.Y(n_895), .A(n_891));
  ADDFX1 g17990(.CO(n_893), .S(n_894), .A(n_829), .B(n_861), .CI(n_852));
  ADDFX1 g17991(.CO(n_891), .S(n_892), .A(
    \dot_product_and_ReLU[0].product_terms[177][0] ), .B(n_860), .CI(n_858));
  ADDFX1 g17992(.CO(n_889), .S(n_890), .A(n_871), .B(n_866), .CI(n_864));
  ADDFX1 g17993(.CO(n_888), .S(\level_4_sums[12][6] [0]), .A(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .B(n_853), .CI(n_862));
  MX2XL g17994(.Y(n_887), .A(n_825), .B(
    \dot_product_and_ReLU[9].product_terms[128][1] ), .S0(n_879));
  AOI221X1 g17995(.Y(\level_3_sums[12][19] [3]), .A0(n_842), .A1(n_846), .B0(
    n_873), .B1(n_878), .C0(n_868));
  XNOR2X1 g17996(.Y(\level_3_sums[12][19] [2]), .A(n_878), .B(n_874));
  INVX1 g17997(.Y(n_886), .A(n_883));
  INVX1 g17998(.Y(n_885), .A(n_882));
  ADDFX1 g17999(.CO(n_882), .S(n_883), .A(
    \dot_product_and_ReLU[1].product_terms[176][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[187][0] ), .CI(n_854));
  ADDHX1 g18000(.CO(n_884), .S(n_881), .A(n_839), .B(n_869));
  ADDFX1 g18001(.CO(n_880), .S(\level_4_sums[12][8] [0]), .A(n_1379), .B(n_1440),
     .CI(n_872));
  ADDFX1 g18002(.CO(n_879), .S(n_877), .A(
    \dot_product_and_ReLU[9].product_terms[128][1] ), .B(
    \dot_product_and_ReLU[17].product_terms[140] [0]), .CI(n_863));
  ADDFX1 g18003(.CO(n_875), .S(n_876), .A(
    \dot_product_and_ReLU[5].product_terms[185][0] ), .B(n_827), .CI(n_840));
  ADDFX1 g18004(.CO(n_878), .S(\level_3_sums[12][19] [1]), .A(n_843), .B(n_844),
     .CI(n_851));
  NAND2BX1 g18005(.Y(n_874), .AN(n_868), .B(n_873));
  ADDFX1 g18006(.CO(n_871), .S(n_872), .A(
    \dot_product_and_ReLU[0].product_terms[142][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[134][1] ), .CI(
    \dot_product_and_ReLU[9].product_terms[128][1] ));
  ADDFX1 g18007(.CO(n_869), .S(n_870), .A(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[105][0] ), .CI(n_1420));
  NAND2X1 g18008(.Y(n_873), .A(n_837), .B(n_857));
  NOR2X1 g18009(.Y(n_868), .A(n_837), .B(n_857));
  INVX1 g18010(.Y(n_867), .A(n_859));
  ADDFX1 g18011(.CO(n_865), .S(n_866), .A(
    \dot_product_and_ReLU[2].product_terms[143][0] ), .B(
    \dot_product_and_ReLU[1].product_terms[135][0] ), .CI(n_831));
  ADDFX1 g18012(.CO(n_863), .S(n_864), .A(
    \dot_product_and_ReLU[2].product_terms[134][1] ), .B(
    \dot_product_and_ReLU[0].product_terms[141][0] ), .CI(n_830));
  ADDFX1 g18013(.CO(n_861), .S(n_862), .A(
    \dot_product_and_ReLU[2].product_terms[104] [1]), .B(
    \dot_product_and_ReLU[3].product_terms[110][0] ), .CI(
    \dot_product_and_ReLU[1].product_terms[108][0] ));
  ADDFX1 g18014(.CO(n_859), .S(n_860), .A(
    \dot_product_and_ReLU[8].product_terms[180][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .CI(
    \dot_product_and_ReLU[0].product_terms[189][0] ));
  XNOR2X1 g18015(.Y(n_858), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\level_1_sums[12][95] [0]));
  XNOR2X1 g18016(.Y(n_857), .A(n_841), .B(n_846));
  ADDHX1 g18017(.CO(n_855), .S(n_856), .A(
    \dot_product_and_ReLU[6].product_terms[188][1] ), .B(n_833));
  NAND2X1 g18018(.Y(n_854), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\level_1_sums[12][95] [0]));
  XNOR2X1 g18019(.Y(\level_3_sums[12][19] [0]), .A(
    \dot_product_and_ReLU[0].product_terms[155][0] ), .B(n_845));
  XOR2XL g18020(.Y(n_853), .A(\dot_product_and_ReLU[16].product_terms[102][2] ),
     .B(n_1231));
  INVX1 g18021(.Y(n_1421), .A(n_839));
  OR2X1 g18022(.Y(n_1423), .A(n_1424), .B(n_849));
  OAI22X1 g18023(.Y(n_852), .A0(\dot_product_and_ReLU[4].product_terms[98][1] ),
     .A1(n_835), .B0(\dot_product_and_ReLU[5].product_terms[96][0] ), .B1(n_828));
  OAI2BB1X1 g18024(.Y(n_851), .A0N(
    \dot_product_and_ReLU[9].product_terms[152][0] ), .A1N(
    \dot_product_and_ReLU[0].product_terms[155][0] ), .B0(n_848));
  XNOR2X1 g18025(.Y(n_850), .A(\dot_product_and_ReLU[1].product_terms[132][1] ),
     .B(n_836));
  NOR2BX1 g18026(.Y(n_849), .AN(n_1425), .B(
    \dot_product_and_ReLU[3].product_terms[123][1] ));
  NAND2BXL g18027(.Y(n_848), .AN(n_842), .B(
    \dot_product_and_ReLU[17].product_terms[156][2] ));
  OR2X1 g18028(.Y(n_1521), .A(n_834), .B(n_1505));
  OR2X1 g18029(.Y(\level_1_sums[12][95] [0]), .A(n_838), .B(n_840));
  NOR2BX1 g18030(.Y(n_847), .AN(n_836), .B(
    \dot_product_and_ReLU[1].product_terms[132][1] ));
  XNOR2X1 g18031(.Y(n_845), .A(\dot_product_and_ReLU[17].product_terms[156][2] ),
     .B(\dot_product_and_ReLU[9].product_terms[152][0] ));
  CLKXOR2X1 g17896(.Y(n_1231), .A(\dot_product_and_ReLU[5].product_terms[96][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[98][1] ));
  XNOR2X1 g18032(.Y(n_846), .A(\dot_product_and_ReLU[1].product_terms[158][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[155][0] ));
  OAI2BB1X1 g18033(.Y(n_844), .A0N(
    \dot_product_and_ReLU[1].product_terms[158][0] ), .A1N(n_826), .B0(n_841));
  XOR2XL g18034(.Y(n_843), .A(\dot_product_and_ReLU[18].product_terms[153][0] ),
     .B(\dot_product_and_ReLU[14].product_terms[154][0] ));
  NOR2BX1 g18035(.Y(n_838), .AN(\dot_product_and_ReLU[4].product_terms[190][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[191][1] ));
  NOR2BX1 g17902(.Y(n_1424), .AN(\dot_product_and_ReLU[3].product_terms[123][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[122][0] ));
  NOR2XL g18036(.Y(n_842), .A(\dot_product_and_ReLU[0].product_terms[155][0] ),
     .B(\dot_product_and_ReLU[9].product_terms[152][0] ));
  NOR2BX1 g18037(.Y(n_1505), .AN(B[226]), .B(B[227]));
  OR2XL g18038(.Y(n_841), .A(\dot_product_and_ReLU[1].product_terms[158][0] ),
     .B(n_826));
  NOR2BX1 g18039(.Y(n_840), .AN(\dot_product_and_ReLU[0].product_terms[191][1] ),
     .B(\dot_product_and_ReLU[4].product_terms[190][1] ));
  NOR2X1 g18040(.Y(n_839), .A(\dot_product_and_ReLU[0].product_terms[100][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[101][1] ));
  NOR2BX1 g18041(.Y(n_835), .AN(\dot_product_and_ReLU[5].product_terms[96][0] ),
     .B(\dot_product_and_ReLU[16].product_terms[102][2] ));
  AND2X1 g18042(.Y(n_2861_danc), .A(B[233]), .B(B[232]));
  NOR2BX1 g18043(.Y(n_834), .AN(B[227]), .B(B[226]));
  NAND2X1 g18044(.Y(n_837), .A(\dot_product_and_ReLU[14].product_terms[154][0] ),
     .B(\dot_product_and_ReLU[18].product_terms[153][0] ));
  OR2X1 g18045(.Y(n_1425), .A(\dot_product_and_ReLU[0].product_terms[122][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[123][1] ));
  NOR2XL g18046(.Y(n_833), .A(\dot_product_and_ReLU[4].product_terms[190][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[191][1] ));
  NAND2BX1 g18047(.Y(n_836), .AN(\dot_product_and_ReLU[0].product_terms[141][0] ),
     .B(\dot_product_and_ReLU[17].product_terms[140] [0]));
  INVX1 g18048(.Y(n_832), .A(\dot_product_and_ReLU[6].product_terms[188][1] ));
  INVX1 g18049(.Y(n_831), .A(n_1381));
  INVX1 g18050(.Y(n_830), .A(\dot_product_and_ReLU[2].product_terms[129][0] ));
  INVX1 g18051(.Y(n_829), .A(\dot_product_and_ReLU[0].product_terms[106][0] ));
  INVX1 g18052(.Y(n_828), .A(\dot_product_and_ReLU[16].product_terms[102][2] ));
  INVX1 g18053(.Y(n_827), .A(\dot_product_and_ReLU[0].product_terms[179][0] ));
  INVX1 g18054(.Y(n_826), .A(\dot_product_and_ReLU[9].product_terms[152][0] ));
  INVX1 g18055(.Y(n_825), .A(\dot_product_and_ReLU[9].product_terms[128][1] ));
  CLKXOR2X1 g18056(.Y(n_1420), .A(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .B(
    \dot_product_and_ReLU[0].product_terms[100][0] ));
  DFFRHQX1 \out_reg_reg[10][3] (.Q(out[93]), .D(n_818), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][4] (.Q(out[94]), .D(n_823), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][7] (.Q(out[97]), .D(n_817), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][2] (.Q(out[92]), .D(n_819), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][5] (.Q(out[95]), .D(n_821), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][0] (.Q(out[90]), .D(n_822), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][6] (.Q(out[96]), .D(n_820), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[10][1] (.Q(out[91]), .D(n_824), .RN(rst_n), .CK(clk));
  NOR2X1 g16494(.Y(n_824), .A(n_802), .B(n_816));
  AND2XL g16495(.Y(n_823), .A(n_808), .B(n_815));
  NOR2X1 g16496(.Y(n_822), .A(\level_8_sums[10] [0]), .B(n_816));
  NOR2X1 g16497(.Y(n_821), .A(n_811), .B(n_816));
  NOR2X1 g16498(.Y(n_820), .A(n_813), .B(n_816));
  AOI21X1 g16499(.Y(n_819), .A0(n_804), .A1(n_803), .B0(n_816));
  NOR2X1 g16500(.Y(n_818), .A(n_806), .B(n_816));
  NOR3BX1 g16501(.Y(n_817), .AN(\level_8_sums[10] [7]), .B(n_812), .C(n_816));
  INVX1 g16502(.Y(n_816), .A(n_815));
  NOR2X1 g16503(.Y(n_815), .A(\level_8_sums[10] [8]), .B(n_814));
  NOR2BX1 g16504(.Y(n_814), .AN(n_812), .B(\level_8_sums[10] [7]));
  AOI21X1 g16505(.Y(n_813), .A0(\level_8_sums[10] [6]), .A1(n_810), .B0(n_812));
  NOR2X1 g16506(.Y(n_812), .A(\level_8_sums[10] [6]), .B(n_810));
  AOI21X1 g16507(.Y(n_811), .A0(\level_8_sums[10] [5]), .A1(n_807), .B0(n_809));
  INVX1 g16508(.Y(n_810), .A(n_809));
  NOR2X1 g16509(.Y(n_809), .A(\level_8_sums[10] [5]), .B(n_807));
  XNOR2X1 g16510(.Y(n_808), .A(n_805), .B(\level_8_sums[10] [4]));
  NOR2BX1 g16511(.Y(n_807), .AN(\level_8_sums[10] [4]), .B(n_805));
  XNOR2X1 g16512(.Y(n_806), .A(n_803), .B(\level_8_sums[10] [3]));
  NAND2X1 g16513(.Y(n_805), .A(n_803), .B(\level_8_sums[10] [3]));
  NAND2BX1 g16514(.Y(n_804), .AN(n_801), .B(\level_8_sums[10] [2]));
  NAND2BX1 g16515(.Y(n_803), .AN(\level_8_sums[10] [2]), .B(n_801));
  AOI21X1 g16516(.Y(n_802), .A0(\level_8_sums[10] [0]), .A1(
    \level_8_sums[10] [1]), .B0(n_801));
  NOR2X1 g16517(.Y(n_801), .A(\level_8_sums[10] [0]), .B(\level_8_sums[10] [1]));
  AO21XL g18057(.Y(\level_4_sums[9][10] [3]), .A0(n_773), .A1(n_800), .B0(
    \level_4_sums[9][10] [8]));
  NOR2X1 g18058(.Y(\level_4_sums[9][10] [8]), .A(n_773), .B(n_800));
  ADDFX1 g18059(.CO(n_800), .S(\level_4_sums[9][10] [2]), .A(n_779), .B(n_787),
     .CI(n_799));
  ADDFX1 g18060(.CO(n_799), .S(\level_4_sums[9][10] [1]), .A(n_767), .B(n_788),
     .CI(n_789));
  XNOR2X1 g18061(.Y(\level_3_sums[9][8] [7]), .A(n_793), .B(n_798));
  XNOR2X1 g18062(.Y(\level_3_sums[9][8] [3]), .A(n_797), .B(n_795));
  OAI21X1 g18063(.Y(n_798), .A0(n_796), .A1(n_786), .B0(n_791));
  XNOR2X1 g17204(.Y(\level_3_sums[9][8] [2]), .A(n_792), .B(n_794));
  NAND2X1 g18064(.Y(n_797), .A(n_785), .B(n_796));
  NAND2BX1 g18065(.Y(n_796), .AN(n_790), .B(n_792));
  NAND2BX1 g18066(.Y(n_795), .AN(n_786), .B(n_791));
  NAND2BX1 g18067(.Y(n_794), .AN(n_790), .B(n_785));
  XNOR2X1 g17209(.Y(n_793), .A(n_781), .B(n_780));
  ADDFX1 g18068(.CO(n_789), .S(\level_4_sums[9][10] [0]), .A(
    \dot_product_and_ReLU[9].product_terms[163][0] ), .B(n_771), .CI(n_776));
  ADDFX1 g18069(.CO(n_792), .S(\level_3_sums[9][8] [1]), .A(n_769), .B(n_765),
     .CI(n_774));
  ADDFX1 g18070(.CO(n_787), .S(n_788), .A(
    \dot_product_and_ReLU[3].product_terms[168][0] ), .B(n_770), .CI(n_775));
  NAND2X1 g18071(.Y(n_791), .A(n_782), .B(n_784));
  NOR2X1 g18072(.Y(n_790), .A(n_777), .B(n_783));
  NOR2XL g18073(.Y(n_786), .A(n_782), .B(n_784));
  NAND2X1 g18074(.Y(n_785), .A(n_777), .B(n_783));
  ADDFX1 g18075(.CO(n_781), .S(n_784), .A(n_764), .B(n_762), .CI(n_761));
  ADDFX1 g18076(.CO(n_782), .S(n_783), .A(n_746), .B(n_768), .CI(n_747));
  XNOR2X1 g18077(.Y(n_780), .A(n_763), .B(n_778));
  XNOR2X1 g17220(.Y(n_779), .A(\dot_product_and_ReLU[9].product_terms[163][0] ),
     .B(n_772));
  XOR2XL g17221(.Y(n_778), .A(n_766), .B(n_761));
  ADDFX1 g17222(.CO(n_775), .S(n_776), .A(
    \dot_product_and_ReLU[2].product_terms[174][1] ), .B(
    \dot_product_and_ReLU[10].product_terms[172][1] ), .CI(
    \dot_product_and_ReLU[1].product_terms[170][0] ));
  ADDFX1 g17223(.CO(n_777), .S(n_774), .A(
    \dot_product_and_ReLU[4].product_terms[68][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[70][0] ), .CI(n_754));
  NOR2BX1 g17224(.Y(n_773), .AN(n_772), .B(
    \dot_product_and_ReLU[9].product_terms[163][0] ));
  ADDFX1 g17225(.CO(n_770), .S(n_771), .A(
    \dot_product_and_ReLU[4].product_terms[166][0] ), .B(n_753), .CI(n_752));
  ADDFX1 g17226(.CO(n_768), .S(n_769), .A(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .B(
    \dot_product_and_ReLU[0].product_terms[66][0] ), .CI(
    \dot_product_and_ReLU[16].product_terms[71][0] ));
  ADDFX1 g17227(.CO(n_772), .S(n_767), .A(
    \dot_product_and_ReLU[2].product_terms[175][0] ), .B(n_751), .CI(
    \dot_product_and_ReLU[8].product_terms[173][1] ));
  OAI21XL g17228(.Y(n_766), .A0(n_1230), .A1(n_756), .B0(n_755));
  OAI21X1 g17229(.Y(n_765), .A0(n_756), .A1(n_759), .B0(n_755));
  OAI21X1 g17230(.Y(n_764), .A0(n_749), .A1(n_756), .B0(n_755));
  XNOR2X1 g17231(.Y(n_763), .A(n_745), .B(n_760));
  XNOR2X1 g17232(.Y(n_762), .A(n_1230), .B(n_745));
  MXI2XL g17234(.Y(\level_3_sums[9][8] [0]), .A(n_748), .B(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .S0(n_1229));
  XNOR2X1 g17235(.Y(n_761), .A(n_749), .B(n_746));
  OAI21X1 g17237(.Y(n_760), .A0(n_749), .A1(n_757), .B0(n_1230));
  AOI21X1 g17238(.Y(n_1551), .A0(B[234]), .A1(B[235]), .B0(n_758));
  XNOR2X1 g17240(.Y(n_759), .A(\dot_product_and_ReLU[1].product_terms[69][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[65][0] ));
  MX2XL g17241(.Y(n_1229), .A(\dot_product_and_ReLU[0].product_terms[65][0] ),
     .B(n_750), .S0(n_2871_danc));
  INVX1 g17243(.Y(n_1552), .A(n_758));
  OR2X1 g17244(.Y(n_1550), .A(B[232]), .B(B[233]));
  NOR2X1 g17245(.Y(n_758), .A(B[235]), .B(B[234]));
  NOR2X1 g17246(.Y(n_757), .A(\dot_product_and_ReLU[0].product_terms[66][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[65][0] ));
  NOR2X1 g17247(.Y(n_756), .A(\dot_product_and_ReLU[4].product_terms[68][0] ),
     .B(\dot_product_and_ReLU[7].product_terms[64][1] ));
  OR2XL g17249(.Y(n_1537), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[179][0] ));
  NOR2BX1 g17250(.Y(n_1538), .AN(\dot_product_and_ReLU[4].product_terms[190][1] ),
     .B(\dot_product_and_ReLU[0].product_terms[191][1] ));
  NAND2X1 g17251(.Y(n_755), .A(\dot_product_and_ReLU[4].product_terms[68][0] ),
     .B(\dot_product_and_ReLU[7].product_terms[64][1] ));
  NOR2BX1 g17252(.Y(n_754), .AN(\dot_product_and_ReLU[1].product_terms[69][1] ),
     .B(n_750));
  NAND2X1 g17253(.Y(n_1230), .A(\dot_product_and_ReLU[0].product_terms[66][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[65][0] ));
  INVX1 g17254(.Y(n_753), .A(\dot_product_and_ReLU[3].product_terms[164][0] ));
  INVX1 g17255(.Y(n_752), .A(\dot_product_and_ReLU[3].product_terms[161][0] ));
  INVX1 g17256(.Y(n_751), .A(\dot_product_and_ReLU[0].product_terms[169][0] ));
  INVX1 g17257(.Y(n_750), .A(\dot_product_and_ReLU[0].product_terms[65][0] ));
  INVX1 g17259(.Y(n_749), .A(\dot_product_and_ReLU[2].product_terms[70][0] ));
  INVX1 g17260(.Y(n_748), .A(\dot_product_and_ReLU[7].product_terms[64][1] ));
  XOR2XL g18078(.Y(n_747), .A(\dot_product_and_ReLU[2].product_terms[70][0] ),
     .B(n_745));
  NOR2BX1 g17261(.Y(n_746), .AN(n_1230), .B(n_757));
  MXI2XL g17262(.Y(n_745), .A(n_748), .B(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .S0(
    \dot_product_and_ReLU[4].product_terms[68][0] ));
  OR2XL g18079(.Y(n_1522), .A(B[227]), .B(B[226]));
  OR2X1 g18080(.Y(n_1486), .A(B[197]), .B(B[196]));
  NOR2X1 g18081(.Y(n_2787_danc), .A(
    \dot_product_and_ReLU[0].product_terms[17][1] ), .B(n_1192));
  AND2XL g18082(.Y(n_1493), .A(\dot_product_and_ReLU[7].product_terms[57][2] ),
     .B(n_1239));
  NOR2X1 g18083(.Y(n_1488), .A(n_1210), .B(n_1211));
  OR2XL g18084(.Y(n_1416), .A(n_744), .B(n_1417));
  AOI2BB1X1 g18085(.Y(n_1418), .A0N(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .A1N(
    \dot_product_and_ReLU[3].product_terms[86][0] ), .B0(n_1419));
  OR2X1 g18086(.Y(n_1449), .A(\dot_product_and_ReLU[17].product_terms[156][2] ),
     .B(\dot_product_and_ReLU[0].product_terms[157][0] ));
  AND2X1 g18087(.Y(n_1468), .A(n_1239), .B(
    \dot_product_and_ReLU[1].product_terms[56][1] ));
  NOR2BX1 g18088(.Y(n_1417), .AN(\dot_product_and_ReLU[3].product_terms[84][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[85][0] ));
  NOR2BX1 g18089(.Y(n_744), .AN(\dot_product_and_ReLU[1].product_terms[85][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[84][0] ));
  NOR2X1 g18090(.Y(n_1422), .A(\dot_product_and_ReLU[3].product_terms[110][0] ),
     .B(n_1204));
  AND2X1 g18091(.Y(n_1419), .A(\dot_product_and_ReLU[3].product_terms[86][0] ),
     .B(\dot_product_and_ReLU[12].product_terms[87][0] ));
  AO21X1 g18092(.Y(n_1237), .A0(n_735), .A1(n_743), .B0(n_1238));
  NOR2X1 g18093(.Y(n_1238), .A(n_735), .B(n_743));
  ADDFX1 g18094(.CO(n_743), .S(n_1236), .A(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .B(
    \dot_product_and_ReLU[7].product_terms[103][0] ), .CI(n_742));
  NAND2X1 g18095(.Y(n_742), .A(n_741), .B(n_1223));
  AOI21X1 g18096(.Y(n_1450), .A0(\dot_product_and_ReLU[3].product_terms[164][0] ),
     .A1(\dot_product_and_ReLU[2].product_terms[165][0] ), .B0(n_740));
  AOI21X1 g18097(.Y(n_1519), .A0(B[209]), .A1(B[208]), .B0(n_739));
  AOI21X1 g18098(.Y(n_1459), .A0(\dot_product_and_ReLU[0].product_terms[141][0] ),
     .A1(\dot_product_and_ReLU[0].product_terms[142][0] ), .B0(n_737));
  OAI21XL g18099(.Y(n_741), .A0(\dot_product_and_ReLU[4].product_terms[101][1] ),
     .A1(\dot_product_and_ReLU[16].product_terms[102][2] ), .B0(
    \dot_product_and_ReLU[0].product_terms[100][0] ));
  OR2XL g18100(.Y(n_1457), .A(n_736), .B(n_1458));
  AOI21X1 g18101(.Y(n_1455), .A0(\dot_product_and_ReLU[2].product_terms[67][0] ),
     .A1(\dot_product_and_ReLU[0].product_terms[66][0] ), .B0(n_738));
  CLKXOR2X1 g18102(.Y(n_1235), .A(
    \dot_product_and_ReLU[16].product_terms[102][2] ), .B(n_1420));
  INVX1 g18103(.Y(n_1451), .A(n_740));
  INVX1 g16488(.Y(n_1520), .A(n_739));
  NOR2X1 g16489(.Y(n_740), .A(\dot_product_and_ReLU[2].product_terms[165][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[164][0] ));
  NOR2BX1 g16490(.Y(n_1458), .AN(\dot_product_and_ReLU[2].product_terms[70][0] ),
     .B(\dot_product_and_ReLU[16].product_terms[71][0] ));
  NOR2X1 g16491(.Y(n_739), .A(B[209]), .B(B[208]));
  INVX1 g16492(.Y(n_1456), .A(n_738));
  INVX1 g16493(.Y(n_1460), .A(n_737));
  NOR2BX1 g18104(.Y(n_736), .AN(\dot_product_and_ReLU[16].product_terms[71][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[70][0] ));
  NOR2X1 g18105(.Y(n_738), .A(\dot_product_and_ReLU[2].product_terms[67][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[66][0] ));
  NOR2X1 g18106(.Y(n_737), .A(\dot_product_and_ReLU[0].product_terms[141][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[142][0] ));
  INVX1 g18107(.Y(n_735), .A(\dot_product_and_ReLU[4].product_terms[101][1] ));
  DFFRHQX1 \out_reg_reg[0][0] (.Q(out[0]), .D(n_675), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][1] (.Q(out[1]), .D(n_680), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][2] (.Q(out[2]), .D(n_673), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][3] (.Q(out[3]), .D(n_667), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][4] (.Q(out[4]), .D(n_663), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][5] (.Q(out[5]), .D(n_671), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][6] (.Q(out[6]), .D(n_662), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[0][7] (.Q(out[7]), .D(n_659), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][0] (.Q(out[9]), .D(n_672), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][1] (.Q(out[10]), .D(n_666), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][2] (.Q(out[11]), .D(n_665), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][3] (.Q(out[12]), .D(n_661), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][4] (.Q(out[13]), .D(n_670), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][5] (.Q(out[14]), .D(n_660), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][6] (.Q(out[15]), .D(n_669), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[1][7] (.Q(out[16]), .D(n_658), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][0] (.Q(out[27]), .D(n_559), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][1] (.Q(out[28]), .D(n_560), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][2] (.Q(out[29]), .D(n_561), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][3] (.Q(out[30]), .D(n_558), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][4] (.Q(out[31]), .D(n_557), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][5] (.Q(out[32]), .D(n_554), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][6] (.Q(out[33]), .D(n_555), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[3][7] (.Q(out[34]), .D(n_552), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][0] (.Q(out[54]), .D(n_730), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][1] (.Q(out[55]), .D(n_729), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][2] (.Q(out[56]), .D(n_728), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][3] (.Q(out[57]), .D(n_718), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][4] (.Q(out[58]), .D(n_734), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][5] (.Q(out[59]), .D(n_725), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][6] (.Q(out[60]), .D(n_717), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][7] (.Q(out[61]), .D(n_719), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[6][8] (.Q(out[62]), .D(n_724), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][0] (.Q(out[63]), .D(n_694), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][1] (.Q(out[64]), .D(n_692), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][2] (.Q(out[65]), .D(n_690), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][3] (.Q(out[66]), .D(n_688), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][4] (.Q(out[67]), .D(n_689), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][5] (.Q(out[68]), .D(n_695), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][6] (.Q(out[69]), .D(n_693), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[7][7] (.Q(out[70]), .D(n_696), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][0] (.Q(out[72]), .D(n_726), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][1] (.Q(out[73]), .D(n_723), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][2] (.Q(out[74]), .D(n_733), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][3] (.Q(out[75]), .D(n_722), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][4] (.Q(out[76]), .D(n_732), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][5] (.Q(out[77]), .D(n_731), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][6] (.Q(out[78]), .D(n_721), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][7] (.Q(out[79]), .D(n_727), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[8][8] (.Q(out[80]), .D(n_720), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][0] (.Q(out[81]), .D(n_706), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][1] (.Q(out[82]), .D(n_697), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][2] (.Q(out[83]), .D(n_700), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][3] (.Q(out[84]), .D(n_703), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][4] (.Q(out[85]), .D(n_702), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][5] (.Q(out[86]), .D(n_701), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][6] (.Q(out[87]), .D(n_699), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][7] (.Q(out[88]), .D(n_704), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[9][8] (.Q(out[89]), .D(n_698), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][0] (.Q(out[99]), .D(n_713), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][1] (.Q(out[100]), .D(n_708), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][2] (.Q(out[101]), .D(n_712), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][3] (.Q(out[102]), .D(n_711), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][4] (.Q(out[103]), .D(n_707), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][5] (.Q(out[104]), .D(n_710), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][6] (.Q(out[105]), .D(n_714), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[11][7] (.Q(out[106]), .D(n_709), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][0] (.Q(out[108]), .D(n_599), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][1] (.Q(out[109]), .D(n_600), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][2] (.Q(out[110]), .D(n_601), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][3] (.Q(out[111]), .D(n_598), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][4] (.Q(out[112]), .D(n_597), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][5] (.Q(out[113]), .D(n_596), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][6] (.Q(out[114]), .D(n_595), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[12][7] (.Q(out[115]), .D(n_594), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][0] (.Q(out[117]), .D(n_446), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][1] (.Q(out[118]), .D(n_448), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][2] (.Q(out[119]), .D(n_453), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][3] (.Q(out[120]), .D(n_452), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][4] (.Q(out[121]), .D(n_451), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][5] (.Q(out[122]), .D(n_454), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][6] (.Q(out[123]), .D(n_450), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[13][7] (.Q(out[124]), .D(n_447), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][0] (.Q(out[126]), .D(n_313), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][1] (.Q(out[127]), .D(n_317), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][2] (.Q(out[128]), .D(n_285), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][3] (.Q(out[129]), .D(n_307), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][4] (.Q(out[130]), .D(n_280), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][5] (.Q(out[131]), .D(n_306), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][6] (.Q(out[132]), .D(n_279), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[14][7] (.Q(out[133]), .D(n_318), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][0] (.Q(out[135]), .D(n_674), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][1] (.Q(out[136]), .D(n_668), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][2] (.Q(out[137]), .D(n_679), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][3] (.Q(out[138]), .D(n_664), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][4] (.Q(out[139]), .D(n_678), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][5] (.Q(out[140]), .D(n_677), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][6] (.Q(out[141]), .D(n_676), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[15][7] (.Q(out[142]), .D(n_657), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][0] (.Q(out[144]), .D(n_636), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][1] (.Q(out[145]), .D(n_639), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][2] (.Q(out[146]), .D(n_638), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][3] (.Q(out[147]), .D(n_631), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][4] (.Q(out[148]), .D(n_625), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][5] (.Q(out[149]), .D(n_630), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][6] (.Q(out[150]), .D(n_633), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[16][7] (.Q(out[151]), .D(n_626), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][0] (.Q(out[153]), .D(n_282), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][1] (.Q(out[154]), .D(n_283), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][2] (.Q(out[155]), .D(n_315), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][3] (.Q(out[156]), .D(n_314), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][4] (.Q(out[157]), .D(n_287), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][5] (.Q(out[158]), .D(n_309), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][6] (.Q(out[159]), .D(n_316), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][7] (.Q(out[160]), .D(n_286), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[17][8] (.Q(out[161]), .D(n_310), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][0] (.Q(out[162]), .D(n_637), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][1] (.Q(out[163]), .D(n_640), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][2] (.Q(out[164]), .D(n_632), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][3] (.Q(out[165]), .D(n_635), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][4] (.Q(out[166]), .D(n_629), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][5] (.Q(out[167]), .D(n_634), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][6] (.Q(out[168]), .D(n_628), .RN(rst_n), .CK(clk));
  DFFRHQX1 \out_reg_reg[18][7] (.Q(out[169]), .D(n_627), .RN(rst_n), .CK(clk));
  NOR2X1 g21585(.Y(n_734), .A(n_540), .B(n_716));
  NOR2XL g21586(.Y(n_733), .A(n_430), .B(n_715));
  NOR2XL g21587(.Y(n_732), .A(n_545), .B(n_715));
  NOR2BX1 g21588(.Y(n_731), .AN(n_587), .B(n_715));
  NOR2X1 g21589(.Y(n_730), .A(\level_8_sums[6] [0]), .B(n_716));
  NOR2X1 g21590(.Y(n_729), .A(n_360), .B(n_716));
  NOR2BX1 g21591(.Y(n_728), .AN(n_413), .B(n_716));
  NOR2XL g21592(.Y(n_727), .A(n_651), .B(n_715));
  NOR2XL g21593(.Y(n_726), .A(\level_8_sums[8] [0]), .B(n_715));
  NOR2X1 g21594(.Y(n_725), .A(n_581), .B(n_716));
  NOR2X1 g21595(.Y(n_724), .A(n_686), .B(n_716));
  NOR2XL g21596(.Y(n_723), .A(n_338), .B(n_715));
  AOI21X1 g21597(.Y(n_722), .A0(n_474), .A1(n_482), .B0(n_715));
  NOR2XL g21598(.Y(n_721), .A(n_614), .B(n_715));
  NOR2XL g21599(.Y(n_720), .A(n_687), .B(n_715));
  NOR2X1 g21600(.Y(n_719), .A(n_650), .B(n_716));
  NOR2X1 g21601(.Y(n_718), .A(n_490), .B(n_716));
  NOR2X1 g21602(.Y(n_717), .A(n_616), .B(n_716));
  XNOR2X1 g21611(.Y(n_716), .A(\level_8_sums[6] [9]), .B(n_683));
  XNOR2X1 g21612(.Y(n_715), .A(\level_8_sums[8] [9]), .B(n_681));
  NOR2X1 g21621(.Y(n_714), .A(n_613), .B(n_705));
  NOR2X1 g21622(.Y(n_713), .A(\level_8_sums[11] [0]), .B(n_705));
  NOR2X1 g21623(.Y(n_712), .A(n_431), .B(n_705));
  NOR2BX1 g21624(.Y(n_711), .AN(n_491), .B(n_705));
  NOR2X1 g21625(.Y(n_710), .A(n_583), .B(n_705));
  NOR2X1 g21626(.Y(n_709), .A(n_648), .B(n_705));
  NOR2X1 g21627(.Y(n_708), .A(n_339), .B(n_705));
  NOR2X1 g21628(.Y(n_707), .A(n_539), .B(n_705));
  NOR2BX1 g21630(.Y(n_706), .AN(\final_sums[9][0] ), .B(n_691));
  NOR2XL g21639(.Y(n_704), .A(n_617), .B(n_691));
  NOR2BX1 g21640(.Y(n_703), .AN(n_411), .B(n_691));
  NOR2XL g21641(.Y(n_702), .A(n_499), .B(n_691));
  NOR2BX1 g21642(.Y(n_701), .AN(n_541), .B(n_691));
  NOR2XL g21643(.Y(n_700), .A(n_359), .B(n_691));
  NOR2XL g21644(.Y(n_699), .A(n_582), .B(n_691));
  NOR2XL g21645(.Y(n_698), .A(n_647), .B(n_691));
  NOR2XL g21646(.Y(n_697), .A(\level_8_sums[9][1] ), .B(n_691));
  XNOR2X1 g21647(.Y(n_705), .A(\level_8_sums[11] [9]), .B(n_682));
  AND2XL g21648(.Y(n_696), .A(n_649), .B(n_685));
  AND2XL g21649(.Y(n_695), .A(n_584), .B(n_685));
  NOR2XL g21650(.Y(n_694), .A(\level_8_sums[7] [0]), .B(n_684));
  NOR2XL g21651(.Y(n_693), .A(n_615), .B(n_684));
  NOR2XL g21652(.Y(n_692), .A(n_342), .B(n_684));
  NOR2XL g21653(.Y(n_690), .A(n_410), .B(n_684));
  NOR2XL g21654(.Y(n_689), .A(n_538), .B(n_684));
  NOR2XL g21655(.Y(n_688), .A(n_497), .B(n_684));
  XNOR2X1 g21656(.Y(n_687), .A(n_645), .B(\level_8_sums[8] [8]));
  XNOR2X1 g21657(.Y(n_686), .A(n_644), .B(\level_8_sums[6] [8]));
  XNOR2X1 g21658(.Y(n_691), .A(\level_8_sums[9][9] ), .B(n_641));
  INVX1 g21673(.Y(n_684), .A(n_685));
  NAND2X1 g21684(.Y(n_683), .A(n_644), .B(\level_8_sums[6] [8]));
  NAND3BXL g21685(.Y(n_682), .AN(n_606), .B(\level_8_sums[11] [7]), .C(
    \level_8_sums[11] [8]));
  NAND2X1 g21686(.Y(n_681), .A(n_645), .B(\level_8_sums[8] [8]));
  OAI2BB1X1 g21687(.Y(n_685), .A0N(n_608), .A1N(\level_8_sums[7] [7]), .B0(
    \level_8_sums[7] [8]));
  NOR2X1 g21688(.Y(n_680), .A(n_361), .B(n_656));
  NOR2X1 g21689(.Y(n_679), .A(n_428), .B(n_654));
  NOR2X1 g21690(.Y(n_678), .A(n_546), .B(n_654));
  AND2XL g21691(.Y(n_677), .A(n_585), .B(n_653));
  NOR2X1 g21692(.Y(n_676), .A(n_620), .B(n_654));
  NOR2X1 g21693(.Y(n_675), .A(\level_8_sums[0] [0]), .B(n_656));
  NOR2X1 g21694(.Y(n_674), .A(\level_8_sums[15] [0]), .B(n_654));
  AND2XL g21695(.Y(n_673), .A(n_429), .B(n_655));
  NOR2X1 g21696(.Y(n_672), .A(\level_8_sums[1] [0]), .B(n_652));
  NOR2X1 g21697(.Y(n_671), .A(n_589), .B(n_656));
  NOR2X1 g21698(.Y(n_670), .A(n_544), .B(n_652));
  NOR2X1 g21699(.Y(n_669), .A(n_619), .B(n_652));
  NOR2X1 g21700(.Y(n_668), .A(n_347), .B(n_654));
  NOR2X1 g21701(.Y(n_667), .A(n_488), .B(n_656));
  NOR2X1 g21702(.Y(n_666), .A(n_341), .B(n_652));
  NOR2X1 g21703(.Y(n_665), .A(n_414), .B(n_652));
  AOI21X1 g21704(.Y(n_664), .A0(n_473), .A1(n_484), .B0(n_654));
  NOR2X1 g21705(.Y(n_663), .A(n_542), .B(n_656));
  NOR2X1 g21706(.Y(n_662), .A(n_618), .B(n_656));
  NOR2X1 g21707(.Y(n_661), .A(n_500), .B(n_652));
  NOR2X1 g21708(.Y(n_660), .A(n_586), .B(n_652));
  NOR3BX1 g21709(.Y(n_659), .AN(\level_8_sums[0] [7]), .B(n_607), .C(n_656));
  NOR3BX1 g21710(.Y(n_658), .AN(\level_8_sums[1] [7]), .B(n_610), .C(n_652));
  NOR3BX1 g21711(.Y(n_657), .AN(\level_8_sums[15] [7]), .B(n_604), .C(n_654));
  XNOR2X1 g21712(.Y(\level_3_sums[10][22][3] ), .A(n_603), .B(n_646));
  INVX1 g21713(.Y(n_656), .A(n_655));
  INVX1 g21714(.Y(n_654), .A(n_653));
  XNOR2X1 g21715(.Y(n_651), .A(n_611), .B(\level_8_sums[8] [7]));
  NOR2X1 g21716(.Y(n_655), .A(\level_8_sums[0] [8]), .B(n_642));
  AOI21X1 g21717(.Y(n_653), .A0(n_604), .A1(n_275), .B0(\level_8_sums[15] [8]));
  OR2X1 g21718(.Y(n_652), .A(\level_8_sums[1] [8]), .B(n_643));
  XNOR2X1 g21719(.Y(n_650), .A(n_609), .B(\level_8_sums[6] [7]));
  XOR2XL g21720(.Y(n_649), .A(n_608), .B(\level_8_sums[7] [7]));
  XOR2XL g21721(.Y(n_648), .A(n_606), .B(\level_8_sums[11] [7]));
  XNOR2X1 g21722(.Y(n_647), .A(n_605), .B(\level_8_sums[9][8] ));
  ADDFX1 g21723(.CO(n_646), .S(\level_3_sums[10][22][2] ), .A(n_495), .B(n_591),
     .CI(n_576));
  NOR2BX1 g21740(.Y(n_643), .AN(n_610), .B(\level_8_sums[1] [7]));
  NOR2BX1 g21741(.Y(n_642), .AN(n_607), .B(\level_8_sums[0] [7]));
  NAND2X1 g21742(.Y(n_641), .A(n_605), .B(\level_8_sums[9][8] ));
  AND2XL g21743(.Y(n_645), .A(n_611), .B(\level_8_sums[8] [7]));
  AND2XL g21744(.Y(n_644), .A(n_609), .B(\level_8_sums[6] [7]));
  NOR2X1 g21745(.Y(n_640), .A(\level_8_sums[18][1] ), .B(n_622));
  NOR2X1 g21746(.Y(n_639), .A(\level_8_sums[16][1] ), .B(n_624));
  NOR2X1 g21747(.Y(n_638), .A(n_363), .B(n_624));
  AND2XL g21748(.Y(n_637), .A(\final_sums[18][0] ), .B(n_621));
  AND2XL g21749(.Y(n_636), .A(\level_8_sums[16][0] ), .B(n_623));
  NOR2X1 g21750(.Y(n_635), .A(n_427), .B(n_622));
  NOR2X1 g21751(.Y(n_634), .A(n_547), .B(n_622));
  NOR2X1 g21752(.Y(n_633), .A(n_588), .B(n_624));
  AO21XL g21753(.Y(\level_3_sums[10][12] [3]), .A0(n_471), .A1(n_612), .B0(
    \level_3_sums[10][12] [7]));
  NOR2X1 g21754(.Y(n_632), .A(n_340), .B(n_622));
  AOI21X1 g21755(.Y(n_631), .A0(n_389), .A1(n_393), .B0(n_624));
  NOR2X1 g21756(.Y(n_630), .A(n_543), .B(n_624));
  AOI21X1 g21757(.Y(n_629), .A0(n_462), .A1(n_485), .B0(n_622));
  AOI21X1 g21758(.Y(n_628), .A0(n_564), .A1(n_565), .B0(n_622));
  NOR3BX1 g21759(.Y(n_627), .AN(\level_8_sums[18][7] ), .B(n_602), .C(n_622));
  NOR3BX1 g21760(.Y(n_626), .AN(\level_8_sums[16][7] ), .B(n_566), .C(n_624));
  NOR2X1 g21761(.Y(n_625), .A(n_489), .B(n_624));
  INVX1 g21762(.Y(n_624), .A(n_623));
  INVX1 g21763(.Y(n_622), .A(n_621));
  AOI21X1 g21764(.Y(n_620), .A0(n_573), .A1(\level_8_sums[15] [6]), .B0(n_604));
  AOI21X1 g21765(.Y(n_619), .A0(\level_8_sums[1] [6]), .A1(n_568), .B0(n_610));
  NOR2X1 g21766(.Y(\level_3_sums[10][12] [7]), .A(n_471), .B(n_612));
  AOI21X1 g21767(.Y(n_623), .A0(n_566), .A1(n_269), .B0(\level_8_sums[16][8] ));
  AOI2BB1X1 g21768(.Y(n_621), .A0N(n_565), .A1N(\level_8_sums[18][7] ), .B0(
    \level_8_sums[18][8] ));
  AOI21X1 g21769(.Y(n_618), .A0(\level_8_sums[0] [6]), .A1(n_570), .B0(n_607));
  XNOR2X1 g21770(.Y(n_617), .A(n_572), .B(\level_8_sums[9][7] ));
  XNOR2X1 g21771(.Y(n_616), .A(\level_8_sums[6] [6]), .B(n_571));
  XNOR2X1 g21772(.Y(n_615), .A(\level_8_sums[7] [6]), .B(n_578));
  XNOR2X1 g21773(.Y(n_614), .A(n_580), .B(\level_8_sums[8] [6]));
  XNOR2X1 g21774(.Y(n_613), .A(n_579), .B(\level_8_sums[11] [6]));
  ADDFX1 g21775(.CO(n_612), .S(\level_3_sums[10][12] [2]), .A(n_504), .B(n_408),
     .CI(n_575));
  XNOR2X1 g21784(.Y(n_603), .A(n_590), .B(n_509));
  AND2XL g21785(.Y(n_611), .A(n_580), .B(\level_8_sums[8] [6]));
  NOR2X1 g21786(.Y(n_610), .A(\level_8_sums[1] [6]), .B(n_568));
  AND2XL g21787(.Y(n_609), .A(n_571), .B(\level_8_sums[6] [6]));
  AND2XL g21788(.Y(n_608), .A(\level_8_sums[7] [6]), .B(n_578));
  NOR2X1 g21789(.Y(n_607), .A(\level_8_sums[0] [6]), .B(n_570));
  NAND2X1 g21790(.Y(n_606), .A(n_579), .B(\level_8_sums[11] [6]));
  AND2XL g21791(.Y(n_605), .A(n_572), .B(\level_8_sums[9][7] ));
  NOR2X1 g21792(.Y(n_604), .A(n_573), .B(\level_8_sums[15] [6]));
  INVX1 g21793(.Y(n_602), .A(n_565));
  NOR2X1 g21794(.Y(n_601), .A(\level_8_sums[12][2] ), .B(n_592));
  AND2XL g21795(.Y(n_600), .A(\final_sums[12][1] ), .B(n_593));
  AND2XL g21796(.Y(n_599), .A(\final_sums[12][0] ), .B(n_593));
  NOR2X1 g21797(.Y(n_598), .A(n_362), .B(n_592));
  AND2XL g21798(.Y(n_597), .A(n_412), .B(n_593));
  NOR2X1 g21799(.Y(n_596), .A(n_498), .B(n_592));
  AOI21X1 g21800(.Y(n_595), .A0(n_522), .A1(n_536), .B0(n_592));
  NOR3BX1 g21801(.Y(n_594), .AN(\level_8_sums[12][7] ), .B(n_562), .C(n_592));
  OAI211X1 g21802(.Y(\level_3_sums[19][22][3] ), .A0(n_436), .A1(n_556), .B0(
    n_519), .C0(n_563));
  XNOR2X1 g21803(.Y(\level_3_sums[2][17] [3]), .A(n_510), .B(n_574));
  XNOR2X1 g21804(.Y(\level_3_sums[2][12][3] ), .A(n_511), .B(n_577));
  INVX1 g21805(.Y(n_592), .A(n_593));
  ADDFX1 g21806(.CO(n_590), .S(n_591), .A(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .B(n_502), .CI(n_464));
  AOI21X1 g21807(.Y(n_589), .A0(n_531), .A1(\level_8_sums[0] [5]), .B0(n_569));
  AOI21X1 g21808(.Y(n_588), .A0(\level_8_sums[16][6] ), .A1(n_534), .B0(n_566));
  XNOR2X1 g21809(.Y(n_587), .A(n_525), .B(\level_8_sums[8] [5]));
  AOI21X1 g21810(.Y(n_586), .A0(\level_8_sums[1] [5]), .A1(n_529), .B0(n_567));
  AOI2BB1X1 g21811(.Y(n_593), .A0N(n_536), .A1N(\level_8_sums[12][7] ), .B0(
    \level_8_sums[12][9] ));
  XNOR2X1 g21812(.Y(n_585), .A(n_526), .B(\level_8_sums[15] [5]));
  XNOR2X1 g21813(.Y(n_584), .A(\level_8_sums[7] [5]), .B(n_521));
  XNOR2X1 g21814(.Y(n_583), .A(n_520), .B(\level_8_sums[11] [5]));
  XNOR2X1 g21815(.Y(\level_3_sums[19][22][2] ), .A(n_512), .B(n_556));
  XNOR2X1 g21816(.Y(n_582), .A(\level_8_sums[9][6] ), .B(n_532));
  XNOR2X1 g21817(.Y(n_581), .A(n_527), .B(\level_8_sums[6] [5]));
  ADDFX1 g21818(.CO(n_577), .S(\level_3_sums[2][12][2] ), .A(n_407), .B(n_476),
     .CI(n_524));
  ADDFX1 g21819(.CO(n_576), .S(\level_3_sums[10][22][1] ), .A(n_503), .B(n_487),
     .CI(n_494));
  ADDFX1 g21820(.CO(n_575), .S(\level_3_sums[10][12] [1]), .A(n_416), .B(n_505),
     .CI(n_457));
  ADDFX1 g21821(.CO(n_574), .S(\level_3_sums[2][17] [2]), .A(n_422), .B(n_442),
     .CI(n_523));
  NOR2BX1 g21830(.Y(n_580), .AN(\level_8_sums[8] [5]), .B(n_525));
  AND2XL g21831(.Y(n_579), .A(n_520), .B(\level_8_sums[11] [5]));
  NOR2BX1 g21832(.Y(n_578), .AN(\level_8_sums[7] [5]), .B(n_521));
  INVX1 g21833(.Y(n_570), .A(n_569));
  INVX1 g21834(.Y(n_568), .A(n_567));
  NAND2BX1 g21835(.Y(n_564), .AN(n_535), .B(\level_8_sums[18][6] ));
  XNOR2X1 g21836(.Y(\level_3_sums[2][21] [2]), .A(n_517), .B(n_551));
  NAND2X1 g21837(.Y(n_563), .A(n_456), .B(n_556));
  NAND2BX1 g21838(.Y(\level_3_sums[2][21] [3]), .AN(\level_3_sums[2][21] [7]),
     .B(n_553));
  XNOR2X1 g21839(.Y(\level_3_sums[19][8] [2]), .A(n_537), .B(n_548));
  NOR2BX1 g21840(.Y(n_573), .AN(\level_8_sums[15] [5]), .B(n_526));
  AND2XL g21841(.Y(n_572), .A(n_532), .B(\level_8_sums[9][6] ));
  AND2XL g21842(.Y(n_571), .A(n_527), .B(\level_8_sums[6] [5]));
  NOR2X1 g21843(.Y(n_569), .A(n_531), .B(\level_8_sums[0] [5]));
  NOR2X1 g21844(.Y(n_567), .A(\level_8_sums[1] [5]), .B(n_529));
  NOR2X1 g21845(.Y(n_566), .A(n_534), .B(\level_8_sums[16][6] ));
  NAND2BX1 g21846(.Y(n_565), .AN(\level_8_sums[18][6] ), .B(n_535));
  INVX1 g21847(.Y(n_562), .A(n_536));
  AND2XL g21848(.Y(n_561), .A(\level_8_sums[3][2] ), .B(n_550));
  AND2XL g21849(.Y(n_560), .A(\level_8_sums[3][1] ), .B(n_550));
  AND2XL g21850(.Y(n_559), .A(\level_8_sums[3][0] ), .B(n_550));
  NOR2X1 g21851(.Y(n_558), .A(\level_8_sums[3][3] ), .B(n_549));
  NOR2X1 g21852(.Y(n_557), .A(n_346), .B(n_549));
  NOR2X1 g21853(.Y(n_555), .A(n_496), .B(n_549));
  AOI21X1 g21854(.Y(n_554), .A0(n_378), .A1(n_386), .B0(n_549));
  NAND3BXL g21855(.Y(n_553), .AN(n_514), .B(n_515), .C(n_551));
  NOR3BX1 g21856(.Y(n_552), .AN(\level_8_sums[3][7] ), .B(n_465), .C(n_549));
  NOR3BX1 g21857(.Y(\level_3_sums[2][21] [7]), .AN(n_514), .B(n_516), .C(n_551));
  XNOR2X1 g21858(.Y(n_556), .A(n_258), .B(n_518));
  INVX1 g21859(.Y(n_549), .A(n_550));
  ADDFX1 g21860(.CO(n_551), .S(\level_3_sums[2][21] [1]), .A(n_432), .B(n_501),
     .CI(n_409));
  ADDFX1 g21861(.CO(n_548), .S(\level_3_sums[19][8] [1]), .A(n_444), .B(n_406),
     .CI(n_477));
  AOI21X1 g21862(.Y(n_547), .A0(\level_8_sums[18][5] ), .A1(n_485), .B0(n_535));
  AOI21X1 g21863(.Y(n_546), .A0(n_484), .A1(\level_8_sums[15] [4]), .B0(n_526));
  AOI21X1 g21864(.Y(n_545), .A0(\level_8_sums[8] [4]), .A1(n_482), .B0(n_525));
  AOI21X1 g21865(.Y(n_544), .A0(n_468), .A1(\level_8_sums[1] [4]), .B0(n_528));
  AOI21X1 g21866(.Y(n_543), .A0(n_470), .A1(\level_8_sums[16][5] ), .B0(n_533));
  AOI21X1 g21867(.Y(n_550), .A0(n_465), .A1(n_276), .B0(\level_8_sums[3][8] ));
  AOI21X1 g21868(.Y(n_542), .A0(\level_8_sums[0] [4]), .A1(n_472), .B0(n_530));
  XNOR2X1 g21869(.Y(n_541), .A(n_480), .B(\level_8_sums[9][5] ));
  XNOR2X1 g21870(.Y(n_540), .A(n_466), .B(\level_8_sums[6] [4]));
  XNOR2X1 g21871(.Y(n_539), .A(n_483), .B(\level_8_sums[11] [4]));
  XNOR2X1 g21872(.Y(n_538), .A(n_479), .B(\level_8_sums[7] [4]));
  XNOR2X1 g21873(.Y(n_537), .A(n_425), .B(n_508));
  INVX1 g21874(.Y(n_534), .A(n_533));
  INVX1 g21875(.Y(n_531), .A(n_530));
  INVX1 g21876(.Y(n_529), .A(n_528));
  ADDFX1 g21877(.CO(n_524), .S(\level_3_sums[2][12][1] ), .A(n_420), .B(n_416),
     .CI(n_404));
  ADDFX1 g21878(.CO(n_523), .S(\level_3_sums[2][17] [1]), .A(n_278), .B(n_419),
     .CI(n_257));
  NAND2BX1 g21879(.Y(n_522), .AN(n_481), .B(\level_8_sums[12][6] ));
  NAND2BX1 g21880(.Y(n_536), .AN(\level_8_sums[12][6] ), .B(n_481));
  NOR2X1 g21881(.Y(n_535), .A(\level_8_sums[18][5] ), .B(n_485));
  NOR2X1 g21882(.Y(n_533), .A(n_470), .B(\level_8_sums[16][5] ));
  NOR2BX1 g21883(.Y(n_532), .AN(\level_8_sums[9][5] ), .B(n_480));
  NOR2X1 g21884(.Y(n_530), .A(\level_8_sums[0] [4]), .B(n_472));
  NOR2X1 g21885(.Y(n_528), .A(n_468), .B(\level_8_sums[1] [4]));
  AND2XL g21886(.Y(n_527), .A(n_466), .B(\level_8_sums[6] [4]));
  NOR2X1 g21887(.Y(n_526), .A(n_484), .B(\level_8_sums[15] [4]));
  NOR2X1 g21888(.Y(n_525), .A(\level_8_sums[8] [4]), .B(n_482));
  AOI21X1 g21889(.Y(n_519), .A0(n_391), .A1(n_436), .B0(n_512));
  OR2XL g21890(.Y(\level_3_sums[19][22][4] ), .A(n_513), .B(n_493));
  AO21XL g21891(.Y(\level_2_sums[2][32] [2]), .A0(n_325), .A1(n_506), .B0(
    \level_2_sums[2][32] [6]));
  AO21XL g21892(.Y(\level_2_sums[2][41] [2]), .A0(n_295), .A1(n_507), .B0(
    \level_2_sums[2][41] [6]));
  XNOR2X1 g21893(.Y(\level_3_sums[19][22][1] ), .A(n_381), .B(n_493));
  XNOR2X1 g21894(.Y(\level_3_sums[10][22][0] ), .A(
    \dot_product_and_ReLU[8].product_terms[180][0] ), .B(n_486));
  XNOR2X1 g21895(.Y(n_518), .A(n_436), .B(n_492));
  NAND2BX1 g21896(.Y(n_517), .AN(n_516), .B(n_515));
  NAND2X1 g21897(.Y(n_521), .A(n_479), .B(\level_8_sums[7] [4]));
  AND2XL g21898(.Y(n_520), .A(n_483), .B(\level_8_sums[11] [4]));
  NAND4XL g21899(.Y(n_513), .A(n_263), .B(n_290), .C(n_391), .D(n_492));
  NOR2X1 g21900(.Y(\level_2_sums[2][32] [6]), .A(n_325), .B(n_506));
  NOR2X1 g21901(.Y(n_516), .A(n_440), .B(n_469));
  NAND2X1 g21902(.Y(n_515), .A(n_440), .B(n_469));
  AOI21X1 g21903(.Y(n_514), .A0(n_252), .A1(n_441), .B0(n_304));
  NOR2X1 g21904(.Y(\level_2_sums[2][41] [6]), .A(n_295), .B(n_507));
  XNOR2X1 g21905(.Y(\level_3_sums[10][12] [0]), .A(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .B(n_260));
  XNOR2X1 g21906(.Y(n_511), .A(n_443), .B(n_475));
  XNOR2X1 g21907(.Y(n_510), .A(n_426), .B(n_458));
  XNOR2X1 g21908(.Y(n_509), .A(n_460), .B(n_464));
  XNOR2X1 g21909(.Y(n_508), .A(n_383), .B(n_459));
  OAI22X1 g21910(.Y(n_512), .A0(n_415), .A1(n_463), .B0(n_381), .B1(n_353));
  ADDFX1 g21911(.CO(n_507), .S(\level_2_sums[2][41] [1]), .A(n_305), .B(n_337),
     .CI(n_433));
  ADDFX1 g21912(.CO(n_504), .S(n_505), .A(
    \dot_product_and_ReLU[5].product_terms[96][0] ), .B(
    \dot_product_and_ReLU[7].product_terms[103][0] ), .CI(n_402));
  ADDFX1 g21913(.CO(n_502), .S(n_503), .A(
    \dot_product_and_ReLU[8].product_terms[180][0] ), .B(
    \dot_product_and_ReLU[0].product_terms[179][0] ), .CI(n_375));
  ADDFX1 g21914(.CO(n_506), .S(\level_2_sums[2][32] [1]), .A(
    \dot_product_and_ReLU[2].product_terms[129][0] ), .B(n_358), .CI(n_368));
  ADDFX1 g21915(.CO(n_501), .S(\level_3_sums[2][21] [0]), .A(
    \dot_product_and_ReLU[1].product_terms[171][1] ), .B(
    \dot_product_and_ReLU[8].product_terms[173][1] ), .CI(n_254));
  OAI2BB1X1 g21916(.Y(\level_3_sums[19][14] [2]), .A0N(n_373), .A1N(n_382), .B0(
    n_461));
  AOI21X1 g21917(.Y(n_500), .A0(n_388), .A1(\level_8_sums[1] [3]), .B0(n_467));
  NAND2X1 g21918(.Y(\level_2_sums[10][29] [2]), .A(n_367), .B(n_438));
  AOI21XL g21919(.Y(n_499), .A0(n_400), .A1(\level_8_sums[9][4] ), .B0(n_480));
  AOI21X1 g21920(.Y(n_498), .A0(n_399), .A1(\level_8_sums[12][5] ), .B0(n_481));
  AOI21XL g21921(.Y(n_497), .A0(n_387), .A1(\level_8_sums[7] [3]), .B0(n_478));
  AOI21X1 g21922(.Y(n_496), .A0(\level_8_sums[3][6] ), .A1(n_386), .B0(n_465));
  AO21XL g21923(.Y(\level_2_sums[2][45] [2]), .A0(n_262), .A1(n_455), .B0(
    \level_2_sums[2][45] [6]));
  OAI21X1 g21924(.Y(n_495), .A0(n_284), .A1(n_397), .B0(n_290));
  OAI21X1 g21925(.Y(n_494), .A0(n_296), .A1(n_418), .B0(n_330));
  XNOR2X1 g21926(.Y(n_491), .A(n_392), .B(\level_8_sums[11] [3]));
  XNOR2X1 g21927(.Y(n_490), .A(n_398), .B(\level_8_sums[6] [3]));
  XNOR2X1 g21928(.Y(n_489), .A(\level_8_sums[16][4] ), .B(n_393));
  XNOR2X1 g21929(.Y(\level_3_sums[19][14] [1]), .A(n_437), .B(n_445));
  XNOR2X1 g21930(.Y(n_488), .A(n_384), .B(\level_8_sums[0] [3]));
  XNOR2X1 g21932(.Y(n_487), .A(n_352), .B(n_397));
  MXI2XL g21933(.Y(n_486), .A(n_270), .B(
    \dot_product_and_ReLU[3].product_terms[178][0] ), .S0(n_418));
  XOR2XL g21934(.Y(n_493), .A(n_415), .B(n_353));
  XNOR2X1 g21935(.Y(n_492), .A(n_263), .B(n_415));
  INVX1 g21936(.Y(n_479), .A(n_478));
  ADDFX1 g21937(.CO(n_477), .S(\level_3_sums[19][8] [0]), .A(
    \dot_product_and_ReLU[0].product_terms[66][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[70][0] ), .CI(n_334));
  ADDFX1 g21938(.CO(n_475), .S(n_476), .A(
    \dot_product_and_ReLU[4].product_terms[98][1] ), .B(n_365), .CI(n_255));
  NAND2BX1 g21947(.Y(n_474), .AN(n_394), .B(\level_8_sums[8] [3]));
  NAND2BX1 g21948(.Y(n_473), .AN(n_395), .B(\level_8_sums[15] [3]));
  NOR2X1 g21949(.Y(\level_2_sums[2][45] [6]), .A(n_262), .B(n_455));
  NAND2BX1 g21950(.Y(n_485), .AN(\level_8_sums[18][4] ), .B(n_396));
  NAND2BX1 g21951(.Y(n_484), .AN(\level_8_sums[15] [3]), .B(n_395));
  NOR2BX1 g21952(.Y(n_483), .AN(\level_8_sums[11] [3]), .B(n_392));
  NAND2BX1 g21953(.Y(n_482), .AN(\level_8_sums[8] [3]), .B(n_394));
  NOR2X1 g21954(.Y(n_481), .A(n_399), .B(\level_8_sums[12][5] ));
  NOR2X1 g21955(.Y(n_480), .A(n_400), .B(\level_8_sums[9][4] ));
  NOR2X1 g21956(.Y(n_478), .A(n_387), .B(\level_8_sums[7] [3]));
  INVX1 g21957(.Y(n_468), .A(n_467));
  AND2XL g21958(.Y(n_463), .A(n_381), .B(n_353));
  OR4X1 g21959(.Y(\level_3_sums[19][8] [7]), .A(n_364), .B(n_401), .C(n_256), .D(
    n_383));
  XNOR2X1 g21960(.Y(\level_3_sums[19][14] [0]), .A(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .B(n_403));
  NAND2BX1 g21961(.Y(n_462), .AN(n_396), .B(\level_8_sums[18][4] ));
  OAI211X1 g21962(.Y(n_461), .A0(n_373), .A1(n_382), .B0(n_259), .C0(n_449));
  AND2XL g21963(.Y(n_472), .A(n_384), .B(\level_8_sums[0] [3]));
  OAI2BB1X1 g21964(.Y(n_471), .A0N(n_349), .A1N(n_365), .B0(n_301));
  XNOR2X1 g21965(.Y(n_460), .A(\dot_product_and_ReLU[3].product_terms[181][0] ),
     .B(n_424));
  XNOR2X1 g21966(.Y(n_459), .A(n_256), .B(n_421));
  AND2XL g21968(.Y(n_470), .A(\level_8_sums[16][4] ), .B(n_393));
  XNOR2X1 g21969(.Y(n_469), .A(n_252), .B(n_441));
  XNOR2X1 g21970(.Y(n_458), .A(n_423), .B(n_257));
  NOR2X1 g21971(.Y(n_467), .A(n_388), .B(\level_8_sums[1] [3]));
  AND2XL g21972(.Y(n_466), .A(n_398), .B(\level_8_sums[6] [3]));
  NOR2X1 g21973(.Y(n_465), .A(\level_8_sums[3][6] ), .B(n_386));
  OAI21X1 g21974(.Y(n_457), .A0(n_281), .A1(n_417), .B0(n_1223));
  XNOR2X1 g21975(.Y(n_464), .A(n_270), .B(n_405));
  INVX1 g21976(.Y(n_456), .A(n_391));
  ADDFX1 g21977(.CO(n_455), .S(\level_2_sums[2][45] [1]), .A(
    \dot_product_and_ReLU[8].product_terms[180][0] ), .B(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .CI(n_369));
  NOR2X1 g21978(.Y(n_454), .A(\level_8_sums[13][5] ), .B(n_434));
  AND2XL g21979(.Y(n_453), .A(\final_sums[13][2] ), .B(n_435));
  AND2XL g21980(.Y(n_452), .A(\final_sums[13][3] ), .B(n_435));
  AND2XL g21981(.Y(n_451), .A(\final_sums[13][4] ), .B(n_435));
  NOR2X1 g21982(.Y(n_450), .A(n_343), .B(n_434));
  NAND2XL g21983(.Y(n_449), .A(n_437), .B(n_439));
  AND2XL g21984(.Y(n_448), .A(\final_sums[13][1] ), .B(n_435));
  OAI21X1 g21985(.Y(\level_2_sums[10][29] [1]), .A0(n_372), .A1(n_371), .B0(
    n_438));
  NOR3BX1 g21986(.Y(n_447), .AN(\level_8_sums[13][7] ), .B(n_327), .C(n_434));
  NOR2BX1 g21987(.Y(n_446), .AN(\final_sums[13][0] ), .B(n_434));
  NAND2X1 g21988(.Y(n_445), .A(n_439), .B(n_259));
  MX2XL g21989(.Y(n_444), .A(\dot_product_and_ReLU[0].product_terms[65][0] ), .B(
    n_266), .S0(n_256));
  XNOR2X1 g21990(.Y(n_443), .A(n_255), .B(n_377));
  XOR2XL g21991(.Y(n_442), .A(\dot_product_and_ReLU[17].product_terms[140] [0]),
     .B(n_385));
  INVX1 g21992(.Y(n_434), .A(n_435));
  ADDFX1 g21993(.CO(n_433), .S(\level_2_sums[2][41] [0]), .A(
    \dot_product_and_ReLU[3].product_terms[164][0] ), .B(
    \dot_product_and_ReLU[2].product_terms[165][0] ), .CI(n_1384));
  ADDFX1 g21994(.CO(n_441), .S(n_432), .A(
    \dot_product_and_ReLU[0].product_terms[169][0] ), .B(
    \dot_product_and_ReLU[10].product_terms[172][1] ), .CI(
    \dot_product_and_ReLU[3].product_terms[168][0] ));
  AOI21X1 g21995(.Y(n_431), .A0(n_302), .A1(\level_8_sums[11] [2]), .B0(n_392));
  AOI21X1 g21996(.Y(n_430), .A0(n_299), .A1(\level_8_sums[8] [2]), .B0(n_394));
  XNOR2X1 g21997(.Y(n_429), .A(n_320), .B(\level_8_sums[0] [2]));
  AOI21X1 g21998(.Y(n_428), .A0(n_297), .A1(\level_8_sums[15] [2]), .B0(n_395));
  AOI21X1 g21999(.Y(n_427), .A0(n_300), .A1(\level_8_sums[18][3] ), .B0(n_396));
  AOI21X1 g22000(.Y(n_440), .A0(\dot_product_and_ReLU[2].product_terms[174][1] ),
     .A1(\dot_product_and_ReLU[8].product_terms[173][1] ), .B0(n_390));
  NAND2XL g22001(.Y(n_426), .A(\dot_product_and_ReLU[17].product_terms[140] [0]),
     .B(n_385));
  OAI21X1 g22002(.Y(n_425), .A0(n_308), .A1(n_370), .B0(n_329));
  NAND2BX1 g22003(.Y(n_439), .AN(n_382), .B(n_298));
  NAND2X1 g22005(.Y(n_438), .A(n_372), .B(n_371));
  OAI21X1 g22006(.Y(n_424), .A0(n_296), .A1(n_288), .B0(n_330));
  OAI2BB1X1 g22007(.Y(n_423), .A0N(
    \dot_product_and_ReLU[1].product_terms[137][0] ), .A1N(n_374), .B0(n_291));
  OAI21X1 g22008(.Y(n_422), .A0(n_272), .A1(n_323), .B0(n_291));
  OAI211X1 g22009(.Y(n_421), .A0(n_266), .A1(n_319), .B0(n_1230), .C0(n_366));
  OAI2BB1X1 g22010(.Y(n_420), .A0N(
    \dot_product_and_ReLU[4].product_terms[97][0] ), .A1N(
    \dot_product_and_ReLU[16].product_terms[102][2] ), .B0(n_380));
  OAI21X1 g22011(.Y(n_437), .A0(n_328), .A1(n_356), .B0(n_332));
  OAI21X1 g22012(.Y(n_419), .A0(n_323), .A1(n_355), .B0(n_291));
  OAI211X1 g22013(.Y(n_436), .A0(n_263), .A1(n_261), .B0(n_290), .C0(n_1243));
  AOI21X1 g22014(.Y(n_435), .A0(n_327), .A1(n_268), .B0(\level_8_sums[13][8] ));
  XNOR2X1 g22016(.Y(n_414), .A(n_294), .B(\level_8_sums[1] [2]));
  XNOR2X1 g22017(.Y(n_413), .A(n_289), .B(\level_8_sums[6] [2]));
  XNOR2X1 g22018(.Y(n_412), .A(n_322), .B(\level_8_sums[12][4] ));
  XNOR2X1 g22019(.Y(n_411), .A(n_321), .B(\level_8_sums[9][3] ));
  XNOR2X1 g22020(.Y(\level_3_sums[2][12][0] ), .A(n_354), .B(n_350));
  XNOR2X1 g22021(.Y(\level_3_sums[2][17] [0]), .A(n_355), .B(n_351));
  XNOR2X1 g22022(.Y(n_410), .A(n_293), .B(\level_8_sums[7] [2]));
  XNOR2X1 g22023(.Y(\level_3_sums[19][22][0] ), .A(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .B(n_348));
  XNOR2X1 g22024(.Y(n_409), .A(n_292), .B(n_252));
  XOR2XL g22025(.Y(n_408), .A(n_349), .B(n_365));
  OAI2BB1X1 g22026(.Y(n_407), .A0N(
    \dot_product_and_ReLU[5].product_terms[96][0] ), .A1N(
    \dot_product_and_ReLU[4].product_terms[98][1] ), .B0(n_379));
  XNOR2X1 g22027(.Y(n_406), .A(n_1457), .B(n_370));
  OAI22X1 g22028(.Y(n_405), .A0(n_262), .A1(n_375), .B0(
    \dot_product_and_ReLU[8].product_terms[180][0] ), .B1(n_288));
  XNOR2X1 g22029(.Y(n_404), .A(n_277), .B(n_1231));
  XOR2XL g22030(.Y(n_403), .A(\dot_product_and_ReLU[1].product_terms[115][0] ),
     .B(n_356));
  XNOR2X1 g22031(.Y(n_418), .A(\dot_product_and_ReLU[0].product_terms[177][0] ),
     .B(n_376));
  AO22XL g22032(.Y(n_402), .A0(\dot_product_and_ReLU[4].product_terms[98][1] ),
     .A1(n_301), .B0(\dot_product_and_ReLU[4].product_terms[97][0] ), .B1(
    \dot_product_and_ReLU[7].product_terms[103][0] ));
  XNOR2X1 g22033(.Y(n_417), .A(\dot_product_and_ReLU[4].product_terms[98][1] ),
     .B(n_349));
  XNOR2X1 g22035(.Y(n_416), .A(\dot_product_and_ReLU[4].product_terms[101][1] ),
     .B(n_350));
  XNOR2X1 g22036(.Y(n_415), .A(\dot_product_and_ReLU[1].product_terms[176][0] ),
     .B(n_375));
  INVXL g22037(.Y(n_401), .A(n_366));
  NOR2X1 g22038(.Y(n_390), .A(n_304), .B(n_292));
  NAND2BX1 g22039(.Y(n_389), .AN(n_326), .B(\level_8_sums[16][3] ));
  NOR2BX1 g22040(.Y(n_400), .AN(\level_8_sums[9][3] ), .B(n_321));
  NOR2BX1 g22041(.Y(n_399), .AN(\level_8_sums[12][4] ), .B(n_322));
  NOR2BX1 g22042(.Y(n_398), .AN(\level_8_sums[6] [2]), .B(n_289));
  NAND2X1 g22043(.Y(n_397), .A(\dot_product_and_ReLU[0].product_terms[177][0] ),
     .B(n_376));
  NOR2X1 g22044(.Y(n_396), .A(n_300), .B(\level_8_sums[18][3] ));
  NOR2X1 g22045(.Y(n_395), .A(n_297), .B(\level_8_sums[15] [2]));
  NOR2X1 g22046(.Y(n_394), .A(n_299), .B(\level_8_sums[8] [2]));
  NAND2BX1 g22047(.Y(n_393), .AN(\level_8_sums[16][3] ), .B(n_326));
  NOR2X1 g22048(.Y(n_392), .A(n_302), .B(\level_8_sums[11] [2]));
  NAND2X1 g22049(.Y(n_391), .A(\dot_product_and_ReLU[1].product_terms[176][0] ),
     .B(n_375));
  OAI21X1 g22050(.Y(n_380), .A0(\dot_product_and_ReLU[4].product_terms[97][0] ),
     .A1(\dot_product_and_ReLU[16].product_terms[102][2] ), .B0(n_354));
  OAI211X1 g22051(.Y(n_379), .A0(\dot_product_and_ReLU[5].product_terms[96][0] ),
     .A1(\dot_product_and_ReLU[4].product_terms[98][1] ), .B0(
    \dot_product_and_ReLU[0].product_terms[100][0] ), .C0(
    \dot_product_and_ReLU[14].product_terms[99][0] ));
  NAND2BX1 g22052(.Y(n_378), .AN(n_324), .B(\level_8_sums[3][5] ));
  AND2X1 g22053(.Y(n_388), .A(\level_8_sums[1] [2]), .B(n_294));
  AND2XL g22054(.Y(n_387), .A(n_293), .B(\level_8_sums[7] [2]));
  XNOR2X1 g22055(.Y(n_377), .A(\dot_product_and_ReLU[4].product_terms[98][1] ),
     .B(n_357));
  NAND2BX1 g22056(.Y(n_386), .AN(\level_8_sums[3][5] ), .B(n_324));
  XNOR2X1 g22057(.Y(n_385), .A(\dot_product_and_ReLU[2].product_terms[143][0] ),
     .B(n_336));
  NOR2BX1 g22058(.Y(n_384), .AN(\level_8_sums[0] [2]), .B(n_320));
  XNOR2X1 g22059(.Y(n_383), .A(\dot_product_and_ReLU[16].product_terms[71][0] ),
     .B(n_253));
  XNOR2X1 g22060(.Y(n_382), .A(\dot_product_and_ReLU[4].product_terms[118][0] ),
     .B(n_335));
  NAND2X1 g22061(.Y(n_381), .A(\dot_product_and_ReLU[3].product_terms[181][0] ),
     .B(n_376));
  INVX1 g22062(.Y(n_376), .A(n_348));
  INVX1 g22063(.Y(n_375), .A(n_288));
  INVXL g22067(.Y(n_374), .A(n_323));
  OAI21X1 g22068(.Y(n_373), .A0(n_273), .A1(n_328), .B0(n_332));
  OA21X1 g22069(.Y(n_372), .A0(\dot_product_and_ReLU[2].product_terms[117][0] ),
     .A1(n_1412), .B0(n_367));
  AOI22X1 g22070(.Y(n_371), .A0(n_312), .A1(n_1411), .B0(
    \dot_product_and_ReLU[2].product_terms[116][0] ), .B1(
    \dot_product_and_ReLU[2].product_terms[117][0] ));
  AOI22X1 g22071(.Y(n_370), .A0(n_311), .A1(n_2871_danc), .B0(
    \dot_product_and_ReLU[16].product_terms[71][0] ), .B1(
    \dot_product_and_ReLU[0].product_terms[65][0] ));
  OAI2BB1X1 g22072(.Y(n_369), .A0N(
    \dot_product_and_ReLU[18].product_terms[183][1] ), .A1N(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .B0(n_344));
  OAI2BB1X1 g22073(.Y(n_368), .A0N(
    \dot_product_and_ReLU[0].product_terms[130][0] ), .A1N(
    \dot_product_and_ReLU[9].product_terms[128][1] ), .B0(n_345));
  AOI21X1 g22075(.Y(n_1472), .A0(\dot_product_and_ReLU[14].product_terms[18][0] ),
     .A1(\dot_product_and_ReLU[1].product_terms[19][1] ), .B0(n_331));
  NAND2X1 g22093(.Y(n_364), .A(n_266), .B(n_329));
  AOI21X1 g22094(.Y(n_2794_danc), .A0(
    \dot_product_and_ReLU[4].product_terms[3][0] ), .A1(
    \dot_product_and_ReLU[19].product_terms[2][0] ), .B0(n_333));
  AOI21X1 g22095(.Y(n_363), .A0(\level_8_sums[16][1] ), .A1(
    \level_8_sums[16][2] ), .B0(n_326));
  AOI21X1 g22096(.Y(n_362), .A0(\level_8_sums[12][2] ), .A1(
    \level_8_sums[12][3] ), .B0(n_322));
  AOI21X1 g22097(.Y(n_361), .A0(\level_8_sums[0] [0]), .A1(\level_8_sums[0] [1]),
     .B0(n_320));
  AOI21X1 g22098(.Y(n_360), .A0(\level_8_sums[6] [0]), .A1(\level_8_sums[6] [1]),
     .B0(n_289));
  AOI21XL g22099(.Y(n_359), .A0(\level_8_sums[9][1] ), .A1(\level_8_sums[9][2] ),
     .B0(n_321));
  OAI2BB1X1 g22100(.Y(n_358), .A0N(
    \dot_product_and_ReLU[14].product_terms[131][0] ), .A1N(n_274), .B0(n_325));
  NAND2X1 g22101(.Y(n_367), .A(\dot_product_and_ReLU[2].product_terms[117][0] ),
     .B(n_1412));
  NAND2X1 g22102(.Y(n_366), .A(\dot_product_and_ReLU[0].product_terms[66][0] ),
     .B(n_1410));
  OAI2BB1X1 g22103(.Y(n_357), .A0N(
    \dot_product_and_ReLU[5].product_terms[96][0] ), .A1N(
    \level_2_sums[17][25][4] ), .B0(n_1223));
  OAI2BB1X1 g22104(.Y(n_365), .A0N(
    \dot_product_and_ReLU[4].product_terms[97][0] ), .A1N(
    \level_2_sums[17][25][4] ), .B0(n_1223));
  XNOR2X1 g22105(.Y(n_347), .A(\level_8_sums[15] [0]), .B(\level_8_sums[15] [1]));
  AOI21X1 g22106(.Y(n_1545), .A0(B[219]), .A1(B[218]), .B0(n_303));
  AOI21X1 g22107(.Y(n_346), .A0(\level_8_sums[3][3] ), .A1(\level_8_sums[3][4] ),
     .B0(n_324));
  OAI21X1 g22108(.Y(n_345), .A0(\dot_product_and_ReLU[0].product_terms[130][0] ),
     .A1(\dot_product_and_ReLU[9].product_terms[128][1] ), .B0(
    \dot_product_and_ReLU[2].product_terms[129][0] ));
  OAI21XL g22109(.Y(n_344), .A0(\dot_product_and_ReLU[18].product_terms[183][1] ),
     .A1(\dot_product_and_ReLU[3].product_terms[181][0] ), .B0(
    \dot_product_and_ReLU[8].product_terms[182][0] ));
  AOI21X1 g22110(.Y(n_343), .A0(\level_8_sums[13][5] ), .A1(
    \level_8_sums[13][6] ), .B0(n_327));
  XNOR2X1 g22111(.Y(n_342), .A(\level_8_sums[7] [0]), .B(\level_8_sums[7] [1]));
  XNOR2X1 g22112(.Y(n_341), .A(\level_8_sums[1] [0]), .B(\level_8_sums[1] [1]));
  XNOR2X1 g22113(.Y(n_340), .A(\level_8_sums[18][1] ), .B(\level_8_sums[18][2] ));
  XNOR2X1 g22114(.Y(n_339), .A(\level_8_sums[11] [0]), .B(\level_8_sums[11] [1]));
  XNOR2X1 g22115(.Y(n_338), .A(\level_8_sums[8] [0]), .B(\level_8_sums[8] [1]));
  XOR2XL g22116(.Y(\level_2_sums[2][32] [0]), .A(
    \dot_product_and_ReLU[0].product_terms[130][0] ), .B(n_1396));
  XOR2XL g22117(.Y(\level_2_sums[10][29] [0]), .A(
    \dot_product_and_ReLU[2].product_terms[116][0] ), .B(
    \level_2_sums[17][29][1] ));
  OAI2BB1X1 g22119(.Y(n_337), .A0N(
    \dot_product_and_ReLU[0].product_terms[167][0] ), .A1N(n_267), .B0(n_295));
  XNOR2X1 g22120(.Y(n_336), .A(\dot_product_and_ReLU[4].product_terms[136][1] ),
     .B(\dot_product_and_ReLU[1].product_terms[137][0] ));
  MX2XL g22121(.Y(n_335), .A(n_273), .B(
    \dot_product_and_ReLU[0].product_terms[119][0] ), .S0(
    \dot_product_and_ReLU[1].product_terms[115][0] ));
  XNOR2X1 g22122(.Y(n_356), .A(\dot_product_and_ReLU[2].product_terms[117][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[114][1] ));
  MXI2XL g22124(.Y(n_334), .A(n_264), .B(
    \dot_product_and_ReLU[16].product_terms[71][0] ), .S0(n_1229));
  XNOR2X1 g22125(.Y(n_355), .A(\dot_product_and_ReLU[19].product_terms[138][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[141][0] ));
  XOR2XL g22126(.Y(n_354), .A(\dot_product_and_ReLU[14].product_terms[99][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[100][0] ));
  MXI2XL g22127(.Y(n_353), .A(\dot_product_and_ReLU[3].product_terms[181][0] ),
     .B(n_261), .S0(n_1536));
  OAI22X1 g22128(.Y(n_352), .A0(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .A1(n_261), .B0(\dot_product_and_ReLU[3].product_terms[181][0] ), .B1(
    n_270));
  XOR2XL g22129(.Y(n_351), .A(\dot_product_and_ReLU[4].product_terms[136][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[143][0] ));
  XNOR2X1 g22130(.Y(n_350), .A(\dot_product_and_ReLU[4].product_terms[97][0] ),
     .B(\dot_product_and_ReLU[16].product_terms[102][2] ));
  OAI22X1 g22131(.Y(n_349), .A0(\dot_product_and_ReLU[4].product_terms[97][0] ),
     .A1(n_265), .B0(\dot_product_and_ReLU[7].product_terms[103][0] ), .B1(
    n_271));
  XNOR2X1 g22134(.Y(n_348), .A(\dot_product_and_ReLU[18].product_terms[183][1] ),
     .B(\dot_product_and_ReLU[8].product_terms[182][0] ));
  INVX1 g22135(.Y(n_2793_danc), .A(n_333));
  INVX1 g22136(.Y(n_1473), .A(n_331));
  INVX1 g22137(.Y(n_1410), .A(n_319));
  NOR2BX1 g22138(.Y(n_318), .AN(\final_sums[14] [7]), .B(\final_sums[14] [9]));
  NOR2BX1 g22139(.Y(n_317), .AN(\final_sums[14] [1]), .B(\final_sums[14] [9]));
  NOR2BX1 g22140(.Y(n_316), .AN(\final_sums[17] [6]), .B(\final_sums[17] [9]));
  NOR2BX1 g22141(.Y(n_315), .AN(\final_sums[17] [2]), .B(\final_sums[17] [9]));
  NOR2BX1 g22142(.Y(n_314), .AN(\final_sums[17] [3]), .B(\final_sums[17] [9]));
  NOR2BX1 g22143(.Y(n_313), .AN(\final_sums[14] [0]), .B(\final_sums[14] [9]));
  OR2XL g22144(.Y(n_312), .A(\dot_product_and_ReLU[2].product_terms[116][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[117][0] ));
  NAND2X1 g22145(.Y(n_311), .A(n_264), .B(n_266));
  NOR2BX1 g22146(.Y(n_310), .AN(\final_sums[17] [8]), .B(\final_sums[17] [9]));
  NOR2BX1 g22147(.Y(n_309), .AN(\final_sums[17] [5]), .B(\final_sums[17] [9]));
  NOR2XL g22148(.Y(n_308), .A(\dot_product_and_ReLU[2].product_terms[70][0] ),
     .B(\dot_product_and_ReLU[16].product_terms[71][0] ));
  NOR2BX1 g22149(.Y(n_307), .AN(\final_sums[14] [3]), .B(\final_sums[14] [9]));
  NOR2BX1 g22150(.Y(n_306), .AN(\final_sums[14] [5]), .B(\final_sums[14] [9]));
  NOR2X1 g22151(.Y(n_333), .A(\dot_product_and_ReLU[4].product_terms[3][0] ), .B(
    \dot_product_and_ReLU[19].product_terms[2][0] ));
  NAND2XL g22152(.Y(n_332), .A(\dot_product_and_ReLU[4].product_terms[118][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[115][0] ));
  AND2XL g22153(.Y(n_305), .A(\dot_product_and_ReLU[0].product_terms[167][0] ),
     .B(\dot_product_and_ReLU[4].product_terms[166][0] ));
  NOR2X1 g22154(.Y(n_331), .A(\dot_product_and_ReLU[1].product_terms[19][1] ),
     .B(\dot_product_and_ReLU[14].product_terms[18][0] ));
  NAND2XL g22155(.Y(n_330), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[8].product_terms[180][0] ));
  NAND2XL g22156(.Y(n_329), .A(\dot_product_and_ReLU[2].product_terms[70][0] ),
     .B(\dot_product_and_ReLU[16].product_terms[71][0] ));
  NOR2X1 g22157(.Y(n_328), .A(\dot_product_and_ReLU[4].product_terms[118][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[115][0] ));
  NOR2X1 g22158(.Y(n_327), .A(\level_8_sums[13][5] ), .B(\level_8_sums[13][6] ));
  NOR2X1 g22159(.Y(n_326), .A(\level_8_sums[16][1] ), .B(\level_8_sums[16][2] ));
  OR2X1 g22160(.Y(n_325), .A(\dot_product_and_ReLU[14].product_terms[131][0] ),
     .B(n_274));
  NOR2X1 g22161(.Y(n_324), .A(\level_8_sums[3][3] ), .B(\level_8_sums[3][4] ));
  NOR2X1 g22162(.Y(n_323), .A(\dot_product_and_ReLU[4].product_terms[136][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[143][0] ));
  NOR2X1 g22164(.Y(n_322), .A(\level_8_sums[12][2] ), .B(\level_8_sums[12][3] ));
  NOR2XL g22165(.Y(n_321), .A(\level_8_sums[9][1] ), .B(\level_8_sums[9][2] ));
  NOR2X1 g22166(.Y(n_320), .A(\level_8_sums[0] [0]), .B(\level_8_sums[0] [1]));
  NOR2X1 g22167(.Y(n_319), .A(\dot_product_and_ReLU[4].product_terms[68][0] ),
     .B(\dot_product_and_ReLU[1].product_terms[69][1] ));
  INVX1 g22168(.Y(n_1546), .A(n_303));
  NOR2BX1 g22169(.Y(n_287), .AN(\final_sums[17] [4]), .B(\final_sums[17] [9]));
  NOR2BX1 g22170(.Y(n_286), .AN(\final_sums[17] [7]), .B(\final_sums[17] [9]));
  NOR2BX1 g22171(.Y(n_285), .AN(\final_sums[14] [2]), .B(\final_sums[14] [9]));
  NAND2X1 g22172(.Y(n_1435), .A(n_1190), .B(n_1206));
  NOR2XL g22173(.Y(n_284), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[181][0] ));
  NOR2BX1 g22174(.Y(\level_1_sums[2][73] [1]), .AN(
    \dot_product_and_ReLU[1].product_terms[147][0] ), .B(
    \dot_product_and_ReLU[4].product_terms[146][0] ));
  NOR2BX1 g22175(.Y(n_283), .AN(\final_sums[17] [1]), .B(\final_sums[17] [9]));
  NOR2BX1 g22176(.Y(n_282), .AN(\final_sums[17] [0]), .B(\final_sums[17] [9]));
  NOR2XL g22177(.Y(n_281), .A(\dot_product_and_ReLU[16].product_terms[102][2] ),
     .B(\dot_product_and_ReLU[4].product_terms[101][1] ));
  NOR2BX1 g22178(.Y(n_280), .AN(\final_sums[14] [4]), .B(\final_sums[14] [9]));
  NOR2BX1 g22179(.Y(n_279), .AN(\final_sums[14] [6]), .B(\final_sums[14] [9]));
  OR2XL g22180(.Y(n_1548), .A(B[225]), .B(B[224]));
  AND2XL g22181(.Y(n_278), .A(\dot_product_and_ReLU[19].product_terms[138][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[141][0] ));
  NOR2X1 g22182(.Y(n_304), .A(\dot_product_and_ReLU[2].product_terms[174][1] ),
     .B(\dot_product_and_ReLU[8].product_terms[173][1] ));
  NOR2X1 g22183(.Y(n_303), .A(B[219]), .B(B[218]));
  AND2XL g22184(.Y(n_302), .A(\level_8_sums[11] [0]), .B(\level_8_sums[11] [1]));
  NAND2X1 g22185(.Y(n_301), .A(n_271), .B(n_265));
  AND2X1 g22186(.Y(n_300), .A(\level_8_sums[18][2] ), .B(\level_8_sums[18][1] ));
  AND2XL g22187(.Y(n_299), .A(\level_8_sums[8] [0]), .B(\level_8_sums[8] [1]));
  NAND2X1 g22188(.Y(n_298), .A(\dot_product_and_ReLU[0].product_terms[114][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[117][0] ));
  AND2X1 g22189(.Y(n_297), .A(\level_8_sums[15] [1]), .B(\level_8_sums[15] [0]));
  NOR2X1 g22190(.Y(n_296), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[8].product_terms[180][0] ));
  OR2X1 g22191(.Y(n_295), .A(\dot_product_and_ReLU[0].product_terms[167][0] ),
     .B(n_267));
  AND2XL g22192(.Y(n_294), .A(\level_8_sums[1] [0]), .B(\level_8_sums[1] [1]));
  AND2XL g22193(.Y(n_293), .A(\level_8_sums[7] [0]), .B(\level_8_sums[7] [1]));
  NAND2X1 g22194(.Y(n_292), .A(\dot_product_and_ReLU[2].product_terms[175][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[169][0] ));
  NAND2XL g22195(.Y(n_277), .A(\dot_product_and_ReLU[14].product_terms[99][0] ),
     .B(\dot_product_and_ReLU[0].product_terms[100][0] ));
  NAND2X1 g22196(.Y(n_291), .A(\dot_product_and_ReLU[4].product_terms[136][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[143][0] ));
  NAND2X1 g22197(.Y(n_290), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(\dot_product_and_ReLU[3].product_terms[181][0] ));
  NOR2X1 g22198(.Y(n_289), .A(\level_8_sums[6] [0]), .B(\level_8_sums[6] [1]));
  NOR2X1 g22199(.Y(n_288), .A(\dot_product_and_ReLU[8].product_terms[182][0] ),
     .B(\dot_product_and_ReLU[18].product_terms[183][1] ));
  INVX1 g22200(.Y(n_276), .A(\level_8_sums[3][7] ));
  INVX1 g22201(.Y(n_275), .A(\level_8_sums[15] [7]));
  INVX1 g22202(.Y(n_274), .A(\dot_product_and_ReLU[9].product_terms[128][1] ));
  INVX1 g22203(.Y(n_273), .A(\dot_product_and_ReLU[0].product_terms[119][0] ));
  INVX1 g22204(.Y(n_272), .A(\dot_product_and_ReLU[17].product_terms[140] [0]));
  INVX1 g22208(.Y(n_271), .A(\dot_product_and_ReLU[4].product_terms[97][0] ));
  INVX1 g22209(.Y(n_270), .A(\dot_product_and_ReLU[3].product_terms[178][0] ));
  INVX1 g22210(.Y(n_269), .A(\level_8_sums[16][7] ));
  INVX1 g22211(.Y(n_268), .A(\level_8_sums[13][7] ));
  INVX1 g22212(.Y(n_267), .A(\dot_product_and_ReLU[3].product_terms[164][0] ));
  INVX1 g22214(.Y(n_266), .A(\dot_product_and_ReLU[0].product_terms[65][0] ));
  INVX1 g22215(.Y(n_265), .A(\dot_product_and_ReLU[7].product_terms[103][0] ));
  INVX1 g22217(.Y(n_264), .A(\dot_product_and_ReLU[16].product_terms[71][0] ));
  INVX1 g22218(.Y(n_263), .A(\dot_product_and_ReLU[0].product_terms[179][0] ));
  INVX1 g22220(.Y(n_262), .A(\dot_product_and_ReLU[8].product_terms[180][0] ));
  INVX1 g22221(.Y(n_261), .A(\dot_product_and_ReLU[3].product_terms[181][0] ));
  XOR2XL g18108(.Y(n_260), .A(\dot_product_and_ReLU[16].product_terms[102][2] ),
     .B(n_417));
  NAND2BX1 g22222(.Y(n_259), .AN(n_298), .B(n_382));
  MXI2XL g22223(.Y(n_258), .A(n_391), .B(n_456), .S0(n_352));
  MXI2XL g22224(.Y(n_257), .A(n_272), .B(
    \dot_product_and_ReLU[17].product_terms[140] [0]), .S0(n_351));
  MXI2XL g22225(.Y(n_256), .A(n_319), .B(n_1410), .S0(
    \dot_product_and_ReLU[0].product_terms[66][0] ));
  NAND2BX1 g22226(.Y(n_1412), .AN(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .B(n_273));
  CLKXOR2X1 g22227(.Y(n_255), .A(\dot_product_and_ReLU[5].product_terms[96][0] ),
     .B(\level_2_sums[17][25][0] ));
  XOR2XL g22228(.Y(n_254), .A(\dot_product_and_ReLU[0].product_terms[169][0] ),
     .B(\dot_product_and_ReLU[2].product_terms[175][0] ));
  MXI2XL g22229(.Y(n_253), .A(\dot_product_and_ReLU[0].product_terms[65][0] ),
     .B(n_266), .S0(\dot_product_and_ReLU[2].product_terms[70][0] ));
  CLKXOR2X1 g22230(.Y(n_252), .A(\dot_product_and_ReLU[8].product_terms[173][1] ),
     .B(\dot_product_and_ReLU[2].product_terms[174][1] ));
  DFFRX2 \B_reg[7] (.Q(\dot_product_and_ReLU[7].product_terms[7][0] ), .QN(n_251),
     .D(n_64), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[10] (.Q(\dot_product_and_ReLU[7].product_terms[10][0] ), .D(
    in[10]), .SE(updown), .SI(\dot_product_and_ReLU[7].product_terms[10][0] ),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[13] (.Q(n_250), .D(in[13]), .SE(updown), .SI(
    \dot_product_and_ReLU[0].product_terms[13][0] ), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[17] (.Q(\dot_product_and_ReLU[0].product_terms[17][1] ), .D(
    in[17]), .SE(updown), .SI(\dot_product_and_ReLU[0].product_terms[17][1] ),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[36] (.Q(\dot_product_and_ReLU[8].product_terms[36][0] ), .D(
    in[36]), .SE(updown), .SI(\dot_product_and_ReLU[8].product_terms[36][0] ),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[38] (.Q(\dot_product_and_ReLU[7].product_terms[38][1] ), .D(
    in[38]), .SE(updown), .SI(\dot_product_and_ReLU[7].product_terms[38][1] ),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[59] (.Q(\dot_product_and_ReLU[19].product_terms[59][1] ), .D(
    in[59]), .SE(updown), .SI(\dot_product_and_ReLU[19].product_terms[59][1] ),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[65] (.Q(n_249), .D(in[65]), .SE(updown), .SI(
    \dot_product_and_ReLU[0].product_terms[65][0] ), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[66] (.Q(\dot_product_and_ReLU[0].product_terms[66][0] ), .QN(
    n_248), .D(n_135), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[70] (.Q(\dot_product_and_ReLU[2].product_terms[70][0] ), .QN(
    n_247), .D(n_125), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[71] (.Q(n_246), .D(in[71]), .SE(updown), .SI(
    \dot_product_and_ReLU[16].product_terms[71][0] ), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[74] (.Q(n_245), .D(in[74]), .SE(updown), .SI(
    \level_1_sums[4][37][1] ), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[84] (.Q(n_244), .D(in[84]), .SE(updown), .SI(
    \dot_product_and_ReLU[3].product_terms[84][0] ), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[114] (.Q(n_243), .D(in[114]), .SE(updown), .SI(
    \dot_product_and_ReLU[0].product_terms[114][1] ), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[118] (.Q(n_242), .D(in[118]), .SE(updown), .SI(
    \dot_product_and_ReLU[4].product_terms[118][0] ), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[127] (.Q(\dot_product_and_ReLU[4].product_terms[127][0] ), .QN(
    n_241), .D(n_45), .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[147] (.Q(\dot_product_and_ReLU[1].product_terms[147][0] ), .D(
    \dot_product_and_ReLU[1].product_terms[147][0] ), .SE(updown), .SI(in[19]),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[173] (.Q(n_240), .D(
    \dot_product_and_ReLU[8].product_terms[173][1] ), .SE(updown), .SI(in[45]),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[181] (.Q(n_239), .D(
    \dot_product_and_ReLU[3].product_terms[181][0] ), .SE(updown), .SI(in[53]),
     .RN(rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[194] (.Q(B[194]), .D(B[194]), .SE(updown), .SI(in[66]), .RN(
    rst_n), .CK(clk));
  SDFFRHQX1 \B_reg[232] (.Q(B[232]), .D(B[232]), .SE(updown), .SI(in[104]), .RN(
    rst_n), .CK(clk));
  MX2XL g20489(.Y(n_238), .A(B[241]), .B(in[113]), .S0(updown));
  MX2XL g20490(.Y(n_237), .A(\dot_product_and_ReLU[0].product_terms[159][1] ),
     .B(in[31]), .S0(updown));
  MX2XL g20491(.Y(n_236), .A(\dot_product_and_ReLU[5].product_terms[160][1] ),
     .B(in[32]), .S0(updown));
  MX2XL g20492(.Y(n_235), .A(\dot_product_and_ReLU[3].product_terms[161][0] ),
     .B(in[33]), .S0(updown));
  MX2XL g20493(.Y(n_234), .A(\level_1_sums[1][81][0] ), .B(in[34]), .S0(updown));
  MX2XL g20494(.Y(n_233), .A(\dot_product_and_ReLU[9].product_terms[163][0] ),
     .B(in[35]), .S0(updown));
  MX2XL g20495(.Y(n_232), .A(in[32]), .B(
    \dot_product_and_ReLU[8].product_terms[32][1] ), .S0(updown));
  MX2XL g20496(.Y(n_231), .A(\dot_product_and_ReLU[3].product_terms[164][0] ),
     .B(in[36]), .S0(updown));
  MX2XL g20497(.Y(n_230), .A(in[33]), .B(
    \dot_product_and_ReLU[2].product_terms[33][0] ), .S0(updown));
  MX2XL g20498(.Y(n_229), .A(in[34]), .B(
    \dot_product_and_ReLU[2].product_terms[34][0] ), .S0(updown));
  MX2XL g20499(.Y(n_228), .A(\dot_product_and_ReLU[2].product_terms[165][0] ),
     .B(in[37]), .S0(updown));
  MX2XL g20500(.Y(n_227), .A(\dot_product_and_ReLU[4].product_terms[166][0] ),
     .B(in[38]), .S0(updown));
  MX2XL g20501(.Y(n_226), .A(\dot_product_and_ReLU[0].product_terms[167][0] ),
     .B(in[39]), .S0(updown));
  MX2XL g20502(.Y(n_225), .A(\dot_product_and_ReLU[3].product_terms[168][0] ),
     .B(in[40]), .S0(updown));
  MX2XL g20503(.Y(n_224), .A(B[253]), .B(in[125]), .S0(updown));
  MX2XL g20504(.Y(n_223), .A(in[35]), .B(
    \dot_product_and_ReLU[2].product_terms[35][0] ), .S0(updown));
  MX2XL g20505(.Y(n_222), .A(\dot_product_and_ReLU[0].product_terms[169][0] ),
     .B(in[41]), .S0(updown));
  MX2XL g20506(.Y(n_221), .A(\dot_product_and_ReLU[1].product_terms[170][0] ),
     .B(in[42]), .S0(updown));
  MX2XL g20507(.Y(n_220), .A(in[37]), .B(
    \dot_product_and_ReLU[2].product_terms[37][1] ), .S0(updown));
  MX2XL g20508(.Y(n_219), .A(\dot_product_and_ReLU[1].product_terms[171][1] ),
     .B(in[43]), .S0(updown));
  MX2XL g20509(.Y(n_218), .A(\dot_product_and_ReLU[10].product_terms[172][1] ),
     .B(in[44]), .S0(updown));
  MX2XL g20510(.Y(n_217), .A(\dot_product_and_ReLU[2].product_terms[174][1] ),
     .B(in[46]), .S0(updown));
  MX2XL g20511(.Y(n_216), .A(\dot_product_and_ReLU[2].product_terms[175][0] ),
     .B(in[47]), .S0(updown));
  MX2XL g20512(.Y(n_215), .A(in[39]), .B(
    \dot_product_and_ReLU[0].product_terms[39][0] ), .S0(updown));
  MX2XL g20513(.Y(n_214), .A(\dot_product_and_ReLU[1].product_terms[176][0] ),
     .B(in[48]), .S0(updown));
  MX2XL g20514(.Y(n_213), .A(in[40]), .B(
    \dot_product_and_ReLU[2].product_terms[40][0] ), .S0(updown));
  MX2XL g20515(.Y(n_212), .A(\dot_product_and_ReLU[0].product_terms[177][0] ),
     .B(in[49]), .S0(updown));
  MX2XL g20516(.Y(n_211), .A(\dot_product_and_ReLU[3].product_terms[178][0] ),
     .B(in[50]), .S0(updown));
  MX2XL g20517(.Y(n_210), .A(in[41]), .B(
    \dot_product_and_ReLU[0].product_terms[41][0] ), .S0(updown));
  MX2XL g20518(.Y(n_209), .A(\dot_product_and_ReLU[0].product_terms[179][0] ),
     .B(in[51]), .S0(updown));
  MX2XL g20519(.Y(n_208), .A(\dot_product_and_ReLU[8].product_terms[180][0] ),
     .B(in[52]), .S0(updown));
  MX2XL g20520(.Y(n_207), .A(B[249]), .B(in[121]), .S0(updown));
  MX2XL g20521(.Y(n_206), .A(in[42]), .B(
    \dot_product_and_ReLU[0].product_terms[42][1] ), .S0(updown));
  MX2XL g20522(.Y(n_205), .A(\dot_product_and_ReLU[8].product_terms[182][0] ),
     .B(in[54]), .S0(updown));
  MX2XL g20523(.Y(n_204), .A(B[245]), .B(in[117]), .S0(updown));
  MX2XL g20524(.Y(n_203), .A(\dot_product_and_ReLU[18].product_terms[183][1] ),
     .B(in[55]), .S0(updown));
  MX2XL g20525(.Y(n_202), .A(\dot_product_and_ReLU[3].product_terms[184][1] ),
     .B(in[56]), .S0(updown));
  MX2XL g20526(.Y(n_201), .A(in[43]), .B(
    \dot_product_and_ReLU[6].product_terms[43][0] ), .S0(updown));
  MX2XL g20527(.Y(n_200), .A(in[44]), .B(
    \dot_product_and_ReLU[2].product_terms[44][1] ), .S0(updown));
  MX2XL g20528(.Y(n_199), .A(\dot_product_and_ReLU[5].product_terms[185][0] ),
     .B(in[57]), .S0(updown));
  MX2XL g20529(.Y(n_198), .A(\dot_product_and_ReLU[18].product_terms[186][0] ),
     .B(in[58]), .S0(updown));
  MX2XL g20530(.Y(n_197), .A(in[45]), .B(
    \dot_product_and_ReLU[3].product_terms[45][1] ), .S0(updown));
  MX2XL g20531(.Y(n_196), .A(\dot_product_and_ReLU[0].product_terms[187][0] ),
     .B(in[59]), .S0(updown));
  MX2XL g20532(.Y(n_195), .A(\dot_product_and_ReLU[6].product_terms[188][1] ),
     .B(in[60]), .S0(updown));
  MX2XL g20533(.Y(n_194), .A(in[46]), .B(
    \dot_product_and_ReLU[19].product_terms[46][2] ), .S0(updown));
  MX2XL g20534(.Y(n_193), .A(\dot_product_and_ReLU[0].product_terms[189][0] ),
     .B(in[61]), .S0(updown));
  MX2XL g20535(.Y(n_192), .A(\dot_product_and_ReLU[4].product_terms[190][1] ),
     .B(in[62]), .S0(updown));
  MX2XL g20536(.Y(n_191), .A(\dot_product_and_ReLU[0].product_terms[191][1] ),
     .B(in[63]), .S0(updown));
  MX2XL g20537(.Y(n_190), .A(in[48]), .B(
    \dot_product_and_ReLU[19].product_terms[48][1] ), .S0(updown));
  MX2XL g20538(.Y(n_189), .A(B[192]), .B(in[64]), .S0(updown));
  MX2XL g20539(.Y(n_188), .A(B[193]), .B(in[65]), .S0(updown));
  MX2XL g20540(.Y(n_187), .A(in[49]), .B(
    \dot_product_and_ReLU[0].product_terms[49][0] ), .S0(updown));
  MX2XL g20541(.Y(n_186), .A(B[195]), .B(in[67]), .S0(updown));
  MX2XL g20542(.Y(n_185), .A(B[196]), .B(in[68]), .S0(updown));
  MX2XL g20543(.Y(n_184), .A(in[47]), .B(
    \dot_product_and_ReLU[3].product_terms[47][1] ), .S0(updown));
  MX2XL g20544(.Y(n_183), .A(in[50]), .B(
    \dot_product_and_ReLU[11].product_terms[50][0] ), .S0(updown));
  MX2XL g20545(.Y(n_182), .A(B[197]), .B(in[69]), .S0(updown));
  MX2XL g20546(.Y(n_181), .A(B[198]), .B(in[70]), .S0(updown));
  MX2XL g20547(.Y(n_180), .A(B[199]), .B(in[71]), .S0(updown));
  MX2XL g20548(.Y(n_179), .A(B[200]), .B(in[72]), .S0(updown));
  MX2XL g20549(.Y(n_178), .A(in[51]), .B(
    \dot_product_and_ReLU[5].product_terms[51][1] ), .S0(updown));
  MX2XL g20550(.Y(n_177), .A(in[52]), .B(
    \dot_product_and_ReLU[2].product_terms[52][0] ), .S0(updown));
  MX2XL g20551(.Y(n_176), .A(B[201]), .B(in[73]), .S0(updown));
  MX2XL g20552(.Y(n_175), .A(B[202]), .B(in[74]), .S0(updown));
  MX2XL g20553(.Y(n_174), .A(in[53]), .B(
    \dot_product_and_ReLU[17].product_terms[53][1] ), .S0(updown));
  MX2XL g20554(.Y(n_173), .A(B[203]), .B(in[75]), .S0(updown));
  MX2XL g20555(.Y(n_172), .A(B[204]), .B(in[76]), .S0(updown));
  MX2XL g20556(.Y(n_171), .A(in[54]), .B(
    \dot_product_and_ReLU[3].product_terms[54][0] ), .S0(updown));
  MX2XL g20557(.Y(n_170), .A(B[205]), .B(in[77]), .S0(updown));
  MX2XL g20558(.Y(n_169), .A(B[206]), .B(in[78]), .S0(updown));
  MX2XL g20559(.Y(n_168), .A(B[207]), .B(in[79]), .S0(updown));
  MX2XL g20560(.Y(n_167), .A(in[55]), .B(
    \dot_product_and_ReLU[1].product_terms[55][0] ), .S0(updown));
  MX2XL g20561(.Y(n_166), .A(B[208]), .B(in[80]), .S0(updown));
  MX2XL g20562(.Y(n_165), .A(in[56]), .B(
    \dot_product_and_ReLU[1].product_terms[56][1] ), .S0(updown));
  MX2XL g20563(.Y(n_164), .A(B[209]), .B(in[81]), .S0(updown));
  MX2XL g20564(.Y(n_163), .A(B[210]), .B(in[82]), .S0(updown));
  MX2XL g20565(.Y(n_162), .A(in[57]), .B(
    \dot_product_and_ReLU[7].product_terms[57][2] ), .S0(updown));
  MX2XL g20566(.Y(n_161), .A(B[211]), .B(in[83]), .S0(updown));
  MX2XL g20567(.Y(n_160), .A(B[212]), .B(in[84]), .S0(updown));
  MX2XL g20568(.Y(n_159), .A(B[237]), .B(in[109]), .S0(updown));
  MX2XL g20569(.Y(n_158), .A(in[58]), .B(
    \dot_product_and_ReLU[7].product_terms[58][0] ), .S0(updown));
  MX2XL g20570(.Y(n_157), .A(B[213]), .B(in[85]), .S0(updown));
  MX2XL g20571(.Y(n_156), .A(B[214]), .B(in[86]), .S0(updown));
  MX2XL g20572(.Y(n_155), .A(B[233]), .B(in[105]), .S0(updown));
  MX2XL g20573(.Y(n_154), .A(B[215]), .B(in[87]), .S0(updown));
  MX2XL g20574(.Y(n_153), .A(B[216]), .B(in[88]), .S0(updown));
  MX2XL g20575(.Y(n_152), .A(in[60]), .B(
    \dot_product_and_ReLU[19].product_terms[60][2] ), .S0(updown));
  MX2XL g20576(.Y(n_151), .A(B[217]), .B(in[89]), .S0(updown));
  MX2XL g20577(.Y(n_150), .A(B[218]), .B(in[90]), .S0(updown));
  MX2XL g20578(.Y(n_149), .A(in[61]), .B(
    \dot_product_and_ReLU[15].product_terms[61][1] ), .S0(updown));
  MX2XL g20579(.Y(n_148), .A(B[219]), .B(in[91]), .S0(updown));
  MX2XL g20580(.Y(n_147), .A(B[220]), .B(in[92]), .S0(updown));
  MX2XL g20581(.Y(n_146), .A(in[62]), .B(
    \dot_product_and_ReLU[1].product_terms[62][0] ), .S0(updown));
  MX2XL g20582(.Y(n_145), .A(B[221]), .B(in[93]), .S0(updown));
  MX2XL g20583(.Y(n_144), .A(B[222]), .B(in[94]), .S0(updown));
  MX2XL g20584(.Y(n_143), .A(B[223]), .B(in[95]), .S0(updown));
  MX2XL g20585(.Y(n_142), .A(B[224]), .B(in[96]), .S0(updown));
  MX2XL g20586(.Y(n_141), .A(B[225]), .B(in[97]), .S0(updown));
  MX2XL g20587(.Y(n_140), .A(B[226]), .B(in[98]), .S0(updown));
  MX2XL g20588(.Y(n_139), .A(B[227]), .B(in[99]), .S0(updown));
  MX2XL g20589(.Y(n_138), .A(in[63]), .B(
    \dot_product_and_ReLU[0].product_terms[63][1] ), .S0(updown));
  MX2XL g20590(.Y(n_137), .A(B[228]), .B(in[100]), .S0(updown));
  MX2XL g20591(.Y(n_136), .A(in[64]), .B(
    \dot_product_and_ReLU[7].product_terms[64][1] ), .S0(updown));
  MX2XL g20592(.Y(n_135), .A(in[66]), .B(
    \dot_product_and_ReLU[0].product_terms[66][0] ), .S0(updown));
  MX2XL g20593(.Y(n_134), .A(B[229]), .B(in[101]), .S0(updown));
  MX2XL g20594(.Y(n_133), .A(B[230]), .B(in[102]), .S0(updown));
  MX2XL g20595(.Y(n_132), .A(B[231]), .B(in[103]), .S0(updown));
  MX2XL g20596(.Y(n_131), .A(in[67]), .B(
    \dot_product_and_ReLU[2].product_terms[67][0] ), .S0(updown));
  MX2XL g20597(.Y(n_130), .A(in[68]), .B(
    \dot_product_and_ReLU[4].product_terms[68][0] ), .S0(updown));
  MX2XL g20598(.Y(n_129), .A(B[234]), .B(in[106]), .S0(updown));
  MX2XL g20599(.Y(n_128), .A(in[69]), .B(
    \dot_product_and_ReLU[1].product_terms[69][1] ), .S0(updown));
  MX2XL g20600(.Y(n_127), .A(B[235]), .B(in[107]), .S0(updown));
  MX2XL g20601(.Y(n_126), .A(B[236]), .B(in[108]), .S0(updown));
  MX2XL g20602(.Y(n_125), .A(in[70]), .B(
    \dot_product_and_ReLU[2].product_terms[70][0] ), .S0(updown));
  MX2XL g20603(.Y(n_124), .A(B[238]), .B(in[110]), .S0(updown));
  MX2XL g20604(.Y(n_123), .A(B[239]), .B(in[111]), .S0(updown));
  MX2XL g20605(.Y(n_122), .A(B[240]), .B(in[112]), .S0(updown));
  MX2XL g20606(.Y(n_121), .A(in[72]), .B(
    \dot_product_and_ReLU[5].product_terms[72][0] ), .S0(updown));
  MX2XL g20607(.Y(n_120), .A(in[31]), .B(
    \dot_product_and_ReLU[2].product_terms[31][1] ), .S0(updown));
  MX2XL g20608(.Y(n_119), .A(in[115]), .B(
    \dot_product_and_ReLU[1].product_terms[115][0] ), .S0(updown));
  MX2XL g20609(.Y(n_118), .A(in[73]), .B(
    \dot_product_and_ReLU[1].product_terms[73][0] ), .S0(updown));
  MX2XL g20610(.Y(n_117), .A(B[243]), .B(in[115]), .S0(updown));
  MX2XL g20611(.Y(n_116), .A(B[244]), .B(in[116]), .S0(updown));
  MX2XL g20612(.Y(n_115), .A(B[246]), .B(in[118]), .S0(updown));
  MX2XL g20613(.Y(n_114), .A(B[247]), .B(in[119]), .S0(updown));
  MX2XL g20614(.Y(n_113), .A(B[248]), .B(in[120]), .S0(updown));
  MX2XL g20615(.Y(n_112), .A(in[75]), .B(
    \dot_product_and_ReLU[5].product_terms[75][0] ), .S0(updown));
  MX2XL g20616(.Y(n_111), .A(in[76]), .B(
    \dot_product_and_ReLU[0].product_terms[76][0] ), .S0(updown));
  MX2XL g20617(.Y(n_110), .A(B[250]), .B(in[122]), .S0(updown));
  MX2XL g20618(.Y(n_109), .A(in[77]), .B(
    \dot_product_and_ReLU[1].product_terms[77][0] ), .S0(updown));
  MX2XL g20619(.Y(n_108), .A(B[251]), .B(in[123]), .S0(updown));
  MX2XL g20620(.Y(n_107), .A(B[252]), .B(in[124]), .S0(updown));
  MX2XL g20621(.Y(n_106), .A(in[78]), .B(
    \dot_product_and_ReLU[10].product_terms[78][1] ), .S0(updown));
  MX2XL g20622(.Y(n_105), .A(B[254]), .B(in[126]), .S0(updown));
  MX2XL g20623(.Y(n_104), .A(B[255]), .B(in[127]), .S0(updown));
  MX2XL g20624(.Y(n_103), .A(in[80]), .B(
    \dot_product_and_ReLU[10].product_terms[80][0] ), .S0(updown));
  MX2XL g20625(.Y(n_102), .A(in[81]), .B(
    \dot_product_and_ReLU[3].product_terms[81][0] ), .S0(updown));
  MX2XL g20626(.Y(n_101), .A(in[79]), .B(
    \dot_product_and_ReLU[4].product_terms[79][0] ), .S0(updown));
  MX2XL g20627(.Y(n_100), .A(in[82]), .B(
    \dot_product_and_ReLU[4].product_terms[82][0] ), .S0(updown));
  MX2XL g20628(.Y(n_99), .A(in[83]), .B(
    \dot_product_and_ReLU[3].product_terms[83][0] ), .S0(updown));
  MX2XL g20629(.Y(n_98), .A(in[85]), .B(
    \dot_product_and_ReLU[1].product_terms[85][0] ), .S0(updown));
  MX2XL g20630(.Y(n_97), .A(in[86]), .B(
    \dot_product_and_ReLU[3].product_terms[86][0] ), .S0(updown));
  MX2XL g20631(.Y(n_96), .A(in[87]), .B(
    \dot_product_and_ReLU[12].product_terms[87][0] ), .S0(updown));
  MX2XL g20632(.Y(n_95), .A(in[88]), .B(
    \dot_product_and_ReLU[0].product_terms[88][1] ), .S0(updown));
  MX2XL g20633(.Y(n_94), .A(in[89]), .B(
    \dot_product_and_ReLU[13].product_terms[89][0] ), .S0(updown));
  MX2XL g20634(.Y(n_93), .A(in[90]), .B(
    \dot_product_and_ReLU[0].product_terms[90][0] ), .S0(updown));
  MX2XL g20635(.Y(n_92), .A(in[91]), .B(
    \dot_product_and_ReLU[2].product_terms[91][1] ), .S0(updown));
  MX2XL g20636(.Y(n_91), .A(in[92]), .B(
    \dot_product_and_ReLU[8].product_terms[92][1] ), .S0(updown));
  MX2XL g20637(.Y(n_90), .A(in[93]), .B(
    \dot_product_and_ReLU[0].product_terms[93][0] ), .S0(updown));
  MX2XL g20638(.Y(n_89), .A(in[94]), .B(
    \dot_product_and_ReLU[0].product_terms[94][1] ), .S0(updown));
  MX2XL g20639(.Y(n_88), .A(in[2]), .B(
    \dot_product_and_ReLU[19].product_terms[2][0] ), .S0(updown));
  MX2XL g20640(.Y(n_87), .A(in[95]), .B(
    \dot_product_and_ReLU[2].product_terms[95][0] ), .S0(updown));
  MX2XL g20641(.Y(n_86), .A(in[96]), .B(
    \dot_product_and_ReLU[5].product_terms[96][0] ), .S0(updown));
  MX2XL g20642(.Y(n_85), .A(in[97]), .B(
    \dot_product_and_ReLU[4].product_terms[97][0] ), .S0(updown));
  MX2XL g20643(.Y(n_84), .A(in[98]), .B(
    \dot_product_and_ReLU[4].product_terms[98][1] ), .S0(updown));
  MX2XL g20644(.Y(n_83), .A(in[99]), .B(
    \dot_product_and_ReLU[14].product_terms[99][0] ), .S0(updown));
  MX2XL g20645(.Y(n_82), .A(in[100]), .B(
    \dot_product_and_ReLU[0].product_terms[100][0] ), .S0(updown));
  MX2XL g20646(.Y(n_81), .A(in[101]), .B(
    \dot_product_and_ReLU[4].product_terms[101][1] ), .S0(updown));
  MX2XL g20647(.Y(n_80), .A(in[102]), .B(
    \dot_product_and_ReLU[16].product_terms[102][2] ), .S0(updown));
  MX2XL g20648(.Y(n_79), .A(in[103]), .B(
    \dot_product_and_ReLU[7].product_terms[103][0] ), .S0(updown));
  MX2XL g20649(.Y(n_78), .A(in[1]), .B(
    \dot_product_and_ReLU[4].product_terms[1][0] ), .S0(updown));
  MX2XL g20650(.Y(n_77), .A(in[104]), .B(
    \dot_product_and_ReLU[2].product_terms[104] [1]), .S0(updown));
  MX2XL g20651(.Y(n_76), .A(in[3]), .B(
    \dot_product_and_ReLU[4].product_terms[3][0] ), .S0(updown));
  MX2XL g20652(.Y(n_75), .A(in[4]), .B(
    \dot_product_and_ReLU[2].product_terms[4][0] ), .S0(updown));
  MX2XL g20653(.Y(n_74), .A(in[105]), .B(
    \dot_product_and_ReLU[0].product_terms[105][0] ), .S0(updown));
  MX2XL g20654(.Y(n_73), .A(in[106]), .B(
    \dot_product_and_ReLU[0].product_terms[106][0] ), .S0(updown));
  MX2XL g20655(.Y(n_72), .A(in[5]), .B(
    \dot_product_and_ReLU[0].product_terms[5][0] ), .S0(updown));
  MX2XL g20656(.Y(n_71), .A(in[107]), .B(
    \dot_product_and_ReLU[16].product_terms[107][0] ), .S0(updown));
  MX2XL g20657(.Y(n_70), .A(in[108]), .B(
    \dot_product_and_ReLU[1].product_terms[108][0] ), .S0(updown));
  MX2XL g20658(.Y(n_69), .A(in[0]), .B(
    \dot_product_and_ReLU[0].product_terms[0][0] ), .S0(updown));
  MX2XL g20659(.Y(n_68), .A(in[6]), .B(
    \dot_product_and_ReLU[0].product_terms[6][2] ), .S0(updown));
  MX2XL g20660(.Y(n_67), .A(in[109]), .B(
    \dot_product_and_ReLU[7].product_terms[109][1] ), .S0(updown));
  MX2XL g20661(.Y(n_66), .A(in[110]), .B(
    \dot_product_and_ReLU[3].product_terms[110][0] ), .S0(updown));
  MX2XL g20662(.Y(n_65), .A(in[111]), .B(
    \dot_product_and_ReLU[7].product_terms[111][0] ), .S0(updown));
  MX2XL g20663(.Y(n_64), .A(in[7]), .B(
    \dot_product_and_ReLU[7].product_terms[7][0] ), .S0(updown));
  MX2XL g20664(.Y(n_63), .A(in[112]), .B(
    \dot_product_and_ReLU[17].product_terms[112][2] ), .S0(updown));
  MX2XL g20665(.Y(n_62), .A(in[8]), .B(
    \dot_product_and_ReLU[0].product_terms[8][0] ), .S0(updown));
  MX2XL g20666(.Y(n_61), .A(in[113]), .B(
    \dot_product_and_ReLU[2].product_terms[113][1] ), .S0(updown));
  MX2XL g20667(.Y(n_60), .A(in[9]), .B(
    \dot_product_and_ReLU[6].product_terms[9][0] ), .S0(updown));
  MX2XL g20668(.Y(n_59), .A(B[242]), .B(in[114]), .S0(updown));
  MX2XL g20669(.Y(n_58), .A(in[116]), .B(
    \dot_product_and_ReLU[2].product_terms[116][0] ), .S0(updown));
  MX2XL g20670(.Y(n_57), .A(in[117]), .B(
    \dot_product_and_ReLU[2].product_terms[117][0] ), .S0(updown));
  MX2XL g20671(.Y(n_56), .A(in[119]), .B(
    \dot_product_and_ReLU[0].product_terms[119][0] ), .S0(updown));
  MX2XL g20672(.Y(n_55), .A(in[120]), .B(
    \dot_product_and_ReLU[3].product_terms[120][1] ), .S0(updown));
  MX2XL g20673(.Y(n_54), .A(in[11]), .B(
    \dot_product_and_ReLU[1].product_terms[11][1] ), .S0(updown));
  MX2XL g20674(.Y(n_53), .A(in[12]), .B(
    \dot_product_and_ReLU[16].product_terms[12][0] ), .S0(updown));
  MX2XL g20675(.Y(n_52), .A(in[121]), .B(
    \dot_product_and_ReLU[2].product_terms[121][1] ), .S0(updown));
  MX2XL g20676(.Y(n_51), .A(in[122]), .B(
    \dot_product_and_ReLU[0].product_terms[122][0] ), .S0(updown));
  MX2XL g20677(.Y(n_50), .A(in[123]), .B(
    \dot_product_and_ReLU[3].product_terms[123][1] ), .S0(updown));
  MX2XL g20678(.Y(n_49), .A(in[124]), .B(
    \dot_product_and_ReLU[17].product_terms[124][0] ), .S0(updown));
  MX2XL g20679(.Y(n_48), .A(in[14]), .B(
    \dot_product_and_ReLU[6].product_terms[14][1] ), .S0(updown));
  MX2XL g20680(.Y(n_47), .A(in[125]), .B(
    \dot_product_and_ReLU[4].product_terms[125][1] ), .S0(updown));
  MX2XL g20681(.Y(n_46), .A(in[126]), .B(
    \dot_product_and_ReLU[4].product_terms[126][1] ), .S0(updown));
  MX2XL g20682(.Y(n_45), .A(in[127]), .B(
    \dot_product_and_ReLU[4].product_terms[127][0] ), .S0(updown));
  MX2XL g20683(.Y(n_44), .A(in[16]), .B(
    \dot_product_and_ReLU[7].product_terms[16][0] ), .S0(updown));
  MX2XL g20684(.Y(n_43), .A(\dot_product_and_ReLU[9].product_terms[128][1] ), .B(
    in[0]), .S0(updown));
  MX2XL g20685(.Y(n_42), .A(\dot_product_and_ReLU[2].product_terms[129][0] ), .B(
    in[1]), .S0(updown));
  MX2XL g20686(.Y(n_41), .A(\dot_product_and_ReLU[0].product_terms[130][0] ), .B(
    in[2]), .S0(updown));
  MX2XL g20687(.Y(n_40), .A(\dot_product_and_ReLU[14].product_terms[131][0] ),
     .B(in[3]), .S0(updown));
  MX2XL g20688(.Y(n_39), .A(\dot_product_and_ReLU[1].product_terms[132][1] ), .B(
    in[4]), .S0(updown));
  MX2XL g20689(.Y(n_38), .A(in[15]), .B(
    \dot_product_and_ReLU[4].product_terms[15][0] ), .S0(updown));
  MX2XL g20690(.Y(n_37), .A(in[18]), .B(
    \dot_product_and_ReLU[14].product_terms[18][0] ), .S0(updown));
  MX2XL g20691(.Y(n_36), .A(\dot_product_and_ReLU[4].product_terms[133][0] ), .B(
    in[5]), .S0(updown));
  MX2XL g20692(.Y(n_35), .A(\dot_product_and_ReLU[2].product_terms[134][1] ), .B(
    in[6]), .S0(updown));
  MX2XL g20693(.Y(n_34), .A(\dot_product_and_ReLU[1].product_terms[135][0] ), .B(
    in[7]), .S0(updown));
  MX2XL g20694(.Y(n_33), .A(\dot_product_and_ReLU[4].product_terms[136][1] ), .B(
    in[8]), .S0(updown));
  MX2XL g20695(.Y(n_32), .A(in[19]), .B(
    \dot_product_and_ReLU[1].product_terms[19][1] ), .S0(updown));
  MX2XL g20696(.Y(n_31), .A(in[20]), .B(
    \dot_product_and_ReLU[4].product_terms[20][0] ), .S0(updown));
  MX2XL g20697(.Y(n_30), .A(\dot_product_and_ReLU[1].product_terms[137][0] ), .B(
    in[9]), .S0(updown));
  MX2XL g20698(.Y(n_29), .A(\dot_product_and_ReLU[19].product_terms[138][0] ),
     .B(in[10]), .S0(updown));
  MX2XL g20699(.Y(n_28), .A(in[21]), .B(
    \dot_product_and_ReLU[2].product_terms[21][1] ), .S0(updown));
  MX2XL g20700(.Y(n_27), .A(\dot_product_and_ReLU[8].product_terms[139][0] ), .B(
    in[11]), .S0(updown));
  MX2XL g20701(.Y(n_26), .A(\dot_product_and_ReLU[17].product_terms[140] [0]),
     .B(in[12]), .S0(updown));
  MX2XL g20702(.Y(n_25), .A(in[22]), .B(
    \dot_product_and_ReLU[0].product_terms[22][0] ), .S0(updown));
  MX2XL g20703(.Y(n_24), .A(\dot_product_and_ReLU[0].product_terms[141][0] ), .B(
    in[13]), .S0(updown));
  MX2XL g20704(.Y(n_23), .A(\dot_product_and_ReLU[0].product_terms[142][0] ), .B(
    in[14]), .S0(updown));
  MX2XL g20705(.Y(n_22), .A(\dot_product_and_ReLU[2].product_terms[143][0] ), .B(
    in[15]), .S0(updown));
  MX2XL g20706(.Y(n_21), .A(in[23]), .B(
    \dot_product_and_ReLU[0].product_terms[23][0] ), .S0(updown));
  MX2XL g20707(.Y(n_20), .A(\dot_product_and_ReLU[2].product_terms[144][0] ), .B(
    in[16]), .S0(updown));
  MX2XL g20708(.Y(n_19), .A(in[24]), .B(
    \dot_product_and_ReLU[4].product_terms[24][0] ), .S0(updown));
  MX2XL g20709(.Y(n_18), .A(\dot_product_and_ReLU[0].product_terms[145][1] ), .B(
    in[17]), .S0(updown));
  MX2XL g20710(.Y(n_17), .A(\dot_product_and_ReLU[4].product_terms[146][0] ), .B(
    in[18]), .S0(updown));
  MX2XL g20711(.Y(n_16), .A(in[25]), .B(
    \dot_product_and_ReLU[3].product_terms[25][0] ), .S0(updown));
  MX2XL g20712(.Y(n_15), .A(\dot_product_and_ReLU[1].product_terms[148][0] ), .B(
    in[20]), .S0(updown));
  MX2XL g20713(.Y(n_14), .A(in[26]), .B(
    \dot_product_and_ReLU[19].product_terms[26][2] ), .S0(updown));
  MX2XL g20714(.Y(n_13), .A(\dot_product_and_ReLU[1].product_terms[149][0] ), .B(
    in[21]), .S0(updown));
  MX2XL g20715(.Y(n_12), .A(\dot_product_and_ReLU[0].product_terms[150][0] ), .B(
    in[22]), .S0(updown));
  MX2XL g20716(.Y(n_11), .A(\dot_product_and_ReLU[3].product_terms[151][0] ), .B(
    in[23]), .S0(updown));
  MX2XL g20717(.Y(n_10), .A(\dot_product_and_ReLU[9].product_terms[152][0] ), .B(
    in[24]), .S0(updown));
  MX2XL g20718(.Y(n_9), .A(in[27]), .B(
    \dot_product_and_ReLU[0].product_terms[27][0] ), .S0(updown));
  MX2XL g20719(.Y(n_8), .A(in[28]), .B(
    \dot_product_and_ReLU[0].product_terms[28][0] ), .S0(updown));
  MX2XL g20720(.Y(n_7), .A(\dot_product_and_ReLU[18].product_terms[153][0] ), .B(
    in[25]), .S0(updown));
  MX2XL g20721(.Y(n_6), .A(\dot_product_and_ReLU[14].product_terms[154][0] ), .B(
    in[26]), .S0(updown));
  MX2XL g20722(.Y(n_5), .A(in[29]), .B(
    \dot_product_and_ReLU[0].product_terms[29][0] ), .S0(updown));
  MX2XL g20723(.Y(n_4), .A(\dot_product_and_ReLU[0].product_terms[155][0] ), .B(
    in[27]), .S0(updown));
  MX2XL g20724(.Y(n_3), .A(\dot_product_and_ReLU[17].product_terms[156][2] ), .B(
    in[28]), .S0(updown));
  MX2XL g20725(.Y(n_2), .A(in[30]), .B(
    \dot_product_and_ReLU[1].product_terms[30][1] ), .S0(updown));
  MX2XL g20726(.Y(n_1), .A(\dot_product_and_ReLU[0].product_terms[157][0] ), .B(
    in[29]), .S0(updown));
  MX2XL g20727(.Y(n_0), .A(\dot_product_and_ReLU[1].product_terms[158][0] ), .B(
    in[30]), .S0(updown));
  DFFRX2 \B_reg[0] (.Q(\dot_product_and_ReLU[0].product_terms[0][0] ), .QN(
    UNCONNECTED129), .D(n_69), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[1] (.Q(\dot_product_and_ReLU[4].product_terms[1][0] ), .QN(
    UNCONNECTED130), .D(n_78), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[2] (.Q(\dot_product_and_ReLU[19].product_terms[2][0] ), .QN(
    UNCONNECTED131), .D(n_88), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[3] (.Q(\dot_product_and_ReLU[4].product_terms[3][0] ), .QN(
    UNCONNECTED132), .D(n_76), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[4] (.Q(\dot_product_and_ReLU[2].product_terms[4][0] ), .QN(
    UNCONNECTED133), .D(n_75), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[5] (.Q(\dot_product_and_ReLU[0].product_terms[5][0] ), .QN(
    UNCONNECTED134), .D(n_72), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[6] (.Q(\dot_product_and_ReLU[0].product_terms[6][2] ), .QN(
    UNCONNECTED135), .D(n_68), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[8] (.Q(\dot_product_and_ReLU[0].product_terms[8][0] ), .QN(
    UNCONNECTED136), .D(n_62), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[9] (.Q(\dot_product_and_ReLU[6].product_terms[9][0] ), .QN(
    UNCONNECTED137), .D(n_60), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[11] (.Q(\dot_product_and_ReLU[1].product_terms[11][1] ), .QN(
    UNCONNECTED138), .D(n_54), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[12] (.Q(\dot_product_and_ReLU[16].product_terms[12][0] ), .QN(
    UNCONNECTED139), .D(n_53), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[14] (.Q(\dot_product_and_ReLU[6].product_terms[14][1] ), .QN(
    UNCONNECTED140), .D(n_48), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[15] (.Q(\dot_product_and_ReLU[4].product_terms[15][0] ), .QN(
    UNCONNECTED141), .D(n_38), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[16] (.Q(\dot_product_and_ReLU[7].product_terms[16][0] ), .QN(
    UNCONNECTED142), .D(n_44), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[18] (.Q(\dot_product_and_ReLU[14].product_terms[18][0] ), .QN(
    UNCONNECTED143), .D(n_37), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[19] (.Q(\dot_product_and_ReLU[1].product_terms[19][1] ), .QN(
    UNCONNECTED144), .D(n_32), .RN(rst_n), .CK(clk));
  DFFRHQX1 \B_reg[20] (.Q(\dot_product_and_ReLU[4].product_terms[20][0] ), .D(
    n_31), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[21] (.Q(\dot_product_and_ReLU[2].product_terms[21][1] ), .QN(
    UNCONNECTED145), .D(n_28), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[22] (.Q(\dot_product_and_ReLU[0].product_terms[22][0] ), .QN(
    UNCONNECTED146), .D(n_25), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[23] (.Q(\dot_product_and_ReLU[0].product_terms[23][0] ), .QN(
    UNCONNECTED147), .D(n_21), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[24] (.Q(\dot_product_and_ReLU[4].product_terms[24][0] ), .QN(
    UNCONNECTED148), .D(n_19), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[25] (.Q(\dot_product_and_ReLU[3].product_terms[25][0] ), .QN(
    UNCONNECTED149), .D(n_16), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[26] (.Q(\dot_product_and_ReLU[19].product_terms[26][2] ), .QN(
    UNCONNECTED150), .D(n_14), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[27] (.Q(\dot_product_and_ReLU[0].product_terms[27][0] ), .QN(
    UNCONNECTED151), .D(n_9), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[28] (.Q(\dot_product_and_ReLU[0].product_terms[28][0] ), .QN(
    UNCONNECTED152), .D(n_8), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[29] (.Q(\dot_product_and_ReLU[0].product_terms[29][0] ), .QN(
    UNCONNECTED153), .D(n_5), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[30] (.Q(\dot_product_and_ReLU[1].product_terms[30][1] ), .QN(
    UNCONNECTED154), .D(n_2), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[31] (.Q(\dot_product_and_ReLU[2].product_terms[31][1] ), .QN(
    UNCONNECTED155), .D(n_120), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[32] (.Q(\dot_product_and_ReLU[8].product_terms[32][1] ), .QN(
    UNCONNECTED156), .D(n_232), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[33] (.Q(\dot_product_and_ReLU[2].product_terms[33][0] ), .QN(
    UNCONNECTED157), .D(n_230), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[34] (.Q(\dot_product_and_ReLU[2].product_terms[34][0] ), .QN(
    UNCONNECTED158), .D(n_229), .RN(rst_n), .CK(clk));
  DFFRHQX1 \B_reg[35] (.Q(\dot_product_and_ReLU[2].product_terms[35][0] ), .D(
    n_223), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[37] (.Q(\dot_product_and_ReLU[2].product_terms[37][1] ), .QN(
    UNCONNECTED159), .D(n_220), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[39] (.Q(\dot_product_and_ReLU[0].product_terms[39][0] ), .QN(
    UNCONNECTED160), .D(n_215), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[40] (.Q(\dot_product_and_ReLU[2].product_terms[40][0] ), .QN(
    UNCONNECTED161), .D(n_213), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[41] (.Q(\dot_product_and_ReLU[0].product_terms[41][0] ), .QN(
    UNCONNECTED162), .D(n_210), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[42] (.Q(\dot_product_and_ReLU[0].product_terms[42][1] ), .QN(
    UNCONNECTED163), .D(n_206), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[43] (.Q(\dot_product_and_ReLU[6].product_terms[43][0] ), .QN(
    UNCONNECTED164), .D(n_201), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[44] (.Q(\dot_product_and_ReLU[2].product_terms[44][1] ), .QN(
    UNCONNECTED165), .D(n_200), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[45] (.Q(\dot_product_and_ReLU[3].product_terms[45][1] ), .QN(
    UNCONNECTED166), .D(n_197), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[46] (.Q(\dot_product_and_ReLU[19].product_terms[46][2] ), .QN(
    UNCONNECTED167), .D(n_194), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[47] (.Q(\dot_product_and_ReLU[3].product_terms[47][1] ), .QN(
    UNCONNECTED168), .D(n_184), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[48] (.Q(\dot_product_and_ReLU[19].product_terms[48][1] ), .QN(
    UNCONNECTED169), .D(n_190), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[49] (.Q(\dot_product_and_ReLU[0].product_terms[49][0] ), .QN(
    UNCONNECTED170), .D(n_187), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[50] (.Q(\dot_product_and_ReLU[11].product_terms[50][0] ), .QN(
    UNCONNECTED171), .D(n_183), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[51] (.Q(\dot_product_and_ReLU[5].product_terms[51][1] ), .QN(
    UNCONNECTED172), .D(n_178), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[52] (.Q(\dot_product_and_ReLU[2].product_terms[52][0] ), .QN(
    UNCONNECTED173), .D(n_177), .RN(rst_n), .CK(clk));
  DFFRHQX1 \B_reg[53] (.Q(\dot_product_and_ReLU[17].product_terms[53][1] ), .D(
    n_174), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[54] (.Q(\dot_product_and_ReLU[3].product_terms[54][0] ), .QN(
    UNCONNECTED174), .D(n_171), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[55] (.Q(\dot_product_and_ReLU[1].product_terms[55][0] ), .QN(
    UNCONNECTED175), .D(n_167), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[56] (.Q(\dot_product_and_ReLU[1].product_terms[56][1] ), .QN(
    UNCONNECTED176), .D(n_165), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[57] (.Q(\dot_product_and_ReLU[7].product_terms[57][2] ), .QN(
    UNCONNECTED177), .D(n_162), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[58] (.Q(\dot_product_and_ReLU[7].product_terms[58][0] ), .QN(
    UNCONNECTED178), .D(n_158), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[60] (.Q(\dot_product_and_ReLU[19].product_terms[60][2] ), .QN(
    UNCONNECTED179), .D(n_152), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[61] (.Q(\dot_product_and_ReLU[15].product_terms[61][1] ), .QN(
    UNCONNECTED180), .D(n_149), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[62] (.Q(\dot_product_and_ReLU[1].product_terms[62][0] ), .QN(
    UNCONNECTED181), .D(n_146), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[63] (.Q(\dot_product_and_ReLU[0].product_terms[63][1] ), .QN(
    UNCONNECTED182), .D(n_138), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[64] (.Q(\dot_product_and_ReLU[7].product_terms[64][1] ), .QN(
    UNCONNECTED183), .D(n_136), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[67] (.Q(\dot_product_and_ReLU[2].product_terms[67][0] ), .QN(
    UNCONNECTED184), .D(n_131), .RN(rst_n), .CK(clk));
  DFFRHQX1 \B_reg[68] (.Q(\dot_product_and_ReLU[4].product_terms[68][0] ), .D(
    n_130), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[69] (.Q(\dot_product_and_ReLU[1].product_terms[69][1] ), .QN(
    UNCONNECTED185), .D(n_128), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[72] (.Q(\dot_product_and_ReLU[5].product_terms[72][0] ), .QN(
    UNCONNECTED186), .D(n_121), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[73] (.Q(\dot_product_and_ReLU[1].product_terms[73][0] ), .QN(
    UNCONNECTED187), .D(n_118), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[75] (.Q(\dot_product_and_ReLU[5].product_terms[75][0] ), .QN(
    UNCONNECTED188), .D(n_112), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[76] (.Q(\dot_product_and_ReLU[0].product_terms[76][0] ), .QN(
    UNCONNECTED189), .D(n_111), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[77] (.Q(\dot_product_and_ReLU[1].product_terms[77][0] ), .QN(
    UNCONNECTED190), .D(n_109), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[78] (.Q(\dot_product_and_ReLU[10].product_terms[78][1] ), .QN(
    UNCONNECTED191), .D(n_106), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[79] (.Q(\dot_product_and_ReLU[4].product_terms[79][0] ), .QN(
    UNCONNECTED192), .D(n_101), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[80] (.Q(\dot_product_and_ReLU[10].product_terms[80][0] ), .QN(
    UNCONNECTED193), .D(n_103), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[81] (.Q(\dot_product_and_ReLU[3].product_terms[81][0] ), .QN(
    UNCONNECTED194), .D(n_102), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[82] (.Q(\dot_product_and_ReLU[4].product_terms[82][0] ), .QN(
    UNCONNECTED195), .D(n_100), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[83] (.Q(\dot_product_and_ReLU[3].product_terms[83][0] ), .QN(
    UNCONNECTED196), .D(n_99), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[85] (.Q(\dot_product_and_ReLU[1].product_terms[85][0] ), .QN(
    UNCONNECTED197), .D(n_98), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[86] (.Q(\dot_product_and_ReLU[3].product_terms[86][0] ), .QN(
    UNCONNECTED198), .D(n_97), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[87] (.Q(\dot_product_and_ReLU[12].product_terms[87][0] ), .QN(
    UNCONNECTED199), .D(n_96), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[88] (.Q(\dot_product_and_ReLU[0].product_terms[88][1] ), .QN(
    UNCONNECTED200), .D(n_95), .RN(rst_n), .CK(clk));
  DFFRHQX1 \B_reg[89] (.Q(\dot_product_and_ReLU[13].product_terms[89][0] ), .D(
    n_94), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[90] (.Q(\dot_product_and_ReLU[0].product_terms[90][0] ), .QN(
    UNCONNECTED201), .D(n_93), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[91] (.Q(\dot_product_and_ReLU[2].product_terms[91][1] ), .QN(
    UNCONNECTED202), .D(n_92), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[92] (.Q(\dot_product_and_ReLU[8].product_terms[92][1] ), .QN(
    UNCONNECTED203), .D(n_91), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[93] (.Q(\dot_product_and_ReLU[0].product_terms[93][0] ), .QN(
    UNCONNECTED204), .D(n_90), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[94] (.Q(\dot_product_and_ReLU[0].product_terms[94][1] ), .QN(
    UNCONNECTED205), .D(n_89), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[95] (.Q(\dot_product_and_ReLU[2].product_terms[95][0] ), .QN(
    UNCONNECTED206), .D(n_87), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[96] (.Q(\dot_product_and_ReLU[5].product_terms[96][0] ), .QN(
    UNCONNECTED207), .D(n_86), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[97] (.Q(\dot_product_and_ReLU[4].product_terms[97][0] ), .QN(
    UNCONNECTED208), .D(n_85), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[98] (.Q(\dot_product_and_ReLU[4].product_terms[98][1] ), .QN(
    UNCONNECTED209), .D(n_84), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[99] (.Q(\dot_product_and_ReLU[14].product_terms[99][0] ), .QN(
    UNCONNECTED210), .D(n_83), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[100] (.Q(\dot_product_and_ReLU[0].product_terms[100][0] ), .QN(
    UNCONNECTED211), .D(n_82), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[101] (.Q(\dot_product_and_ReLU[4].product_terms[101][1] ), .QN(
    UNCONNECTED212), .D(n_81), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[102] (.Q(\dot_product_and_ReLU[16].product_terms[102][2] ), .QN(
    UNCONNECTED213), .D(n_80), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[103] (.Q(\dot_product_and_ReLU[7].product_terms[103][0] ), .QN(
    UNCONNECTED214), .D(n_79), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[104] (.Q(\dot_product_and_ReLU[2].product_terms[104] [1]), .QN(
    UNCONNECTED215), .D(n_77), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[105] (.Q(\dot_product_and_ReLU[0].product_terms[105][0] ), .QN(
    UNCONNECTED216), .D(n_74), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[106] (.Q(\dot_product_and_ReLU[0].product_terms[106][0] ), .QN(
    UNCONNECTED217), .D(n_73), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[107] (.Q(\dot_product_and_ReLU[16].product_terms[107][0] ), .QN(
    UNCONNECTED218), .D(n_71), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[108] (.Q(\dot_product_and_ReLU[1].product_terms[108][0] ), .QN(
    UNCONNECTED219), .D(n_70), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[109] (.Q(\dot_product_and_ReLU[7].product_terms[109][1] ), .QN(
    UNCONNECTED220), .D(n_67), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[110] (.Q(\dot_product_and_ReLU[3].product_terms[110][0] ), .QN(
    UNCONNECTED221), .D(n_66), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[111] (.Q(\dot_product_and_ReLU[7].product_terms[111][0] ), .QN(
    UNCONNECTED222), .D(n_65), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[112] (.Q(\dot_product_and_ReLU[17].product_terms[112][2] ), .QN(
    UNCONNECTED223), .D(n_63), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[113] (.Q(\dot_product_and_ReLU[2].product_terms[113][1] ), .QN(
    UNCONNECTED224), .D(n_61), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[115] (.Q(\dot_product_and_ReLU[1].product_terms[115][0] ), .QN(
    UNCONNECTED225), .D(n_119), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[116] (.Q(\dot_product_and_ReLU[2].product_terms[116][0] ), .QN(
    UNCONNECTED226), .D(n_58), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[117] (.Q(\dot_product_and_ReLU[2].product_terms[117][0] ), .QN(
    UNCONNECTED227), .D(n_57), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[119] (.Q(\dot_product_and_ReLU[0].product_terms[119][0] ), .QN(
    UNCONNECTED228), .D(n_56), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[120] (.Q(\dot_product_and_ReLU[3].product_terms[120][1] ), .QN(
    UNCONNECTED229), .D(n_55), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[121] (.Q(\dot_product_and_ReLU[2].product_terms[121][1] ), .QN(
    UNCONNECTED230), .D(n_52), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[122] (.Q(\dot_product_and_ReLU[0].product_terms[122][0] ), .QN(
    UNCONNECTED231), .D(n_51), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[123] (.Q(\dot_product_and_ReLU[3].product_terms[123][1] ), .QN(
    UNCONNECTED232), .D(n_50), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[124] (.Q(\dot_product_and_ReLU[17].product_terms[124][0] ), .QN(
    UNCONNECTED233), .D(n_49), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[125] (.Q(\dot_product_and_ReLU[4].product_terms[125][1] ), .QN(
    UNCONNECTED234), .D(n_47), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[126] (.Q(\dot_product_and_ReLU[4].product_terms[126][1] ), .QN(
    UNCONNECTED235), .D(n_46), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[128] (.Q(\dot_product_and_ReLU[9].product_terms[128][1] ), .QN(
    UNCONNECTED236), .D(n_43), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[129] (.Q(\dot_product_and_ReLU[2].product_terms[129][0] ), .QN(
    UNCONNECTED237), .D(n_42), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[130] (.Q(\dot_product_and_ReLU[0].product_terms[130][0] ), .QN(
    UNCONNECTED238), .D(n_41), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[131] (.Q(\dot_product_and_ReLU[14].product_terms[131][0] ), .QN(
    UNCONNECTED239), .D(n_40), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[132] (.Q(\dot_product_and_ReLU[1].product_terms[132][1] ), .QN(
    UNCONNECTED240), .D(n_39), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[133] (.Q(\dot_product_and_ReLU[4].product_terms[133][0] ), .QN(
    UNCONNECTED241), .D(n_36), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[134] (.Q(\dot_product_and_ReLU[2].product_terms[134][1] ), .QN(
    UNCONNECTED242), .D(n_35), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[135] (.Q(\dot_product_and_ReLU[1].product_terms[135][0] ), .QN(
    UNCONNECTED243), .D(n_34), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[136] (.Q(\dot_product_and_ReLU[4].product_terms[136][1] ), .QN(
    UNCONNECTED244), .D(n_33), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[137] (.Q(\dot_product_and_ReLU[1].product_terms[137][0] ), .QN(
    UNCONNECTED245), .D(n_30), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[138] (.Q(\dot_product_and_ReLU[19].product_terms[138][0] ), .QN(
    UNCONNECTED246), .D(n_29), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[139] (.Q(\dot_product_and_ReLU[8].product_terms[139][0] ), .QN(
    UNCONNECTED247), .D(n_27), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[140] (.Q(\dot_product_and_ReLU[17].product_terms[140] [0]), .QN(
    UNCONNECTED248), .D(n_26), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[141] (.Q(\dot_product_and_ReLU[0].product_terms[141][0] ), .QN(
    UNCONNECTED249), .D(n_24), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[142] (.Q(\dot_product_and_ReLU[0].product_terms[142][0] ), .QN(
    UNCONNECTED250), .D(n_23), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[143] (.Q(\dot_product_and_ReLU[2].product_terms[143][0] ), .QN(
    UNCONNECTED251), .D(n_22), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[144] (.Q(\dot_product_and_ReLU[2].product_terms[144][0] ), .QN(
    UNCONNECTED252), .D(n_20), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[145] (.Q(\dot_product_and_ReLU[0].product_terms[145][1] ), .QN(
    UNCONNECTED253), .D(n_18), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[146] (.Q(\dot_product_and_ReLU[4].product_terms[146][0] ), .QN(
    UNCONNECTED254), .D(n_17), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[148] (.Q(\dot_product_and_ReLU[1].product_terms[148][0] ), .QN(
    UNCONNECTED255), .D(n_15), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[149] (.Q(\dot_product_and_ReLU[1].product_terms[149][0] ), .QN(
    UNCONNECTED256), .D(n_13), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[150] (.Q(\dot_product_and_ReLU[0].product_terms[150][0] ), .QN(
    UNCONNECTED257), .D(n_12), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[151] (.Q(\dot_product_and_ReLU[3].product_terms[151][0] ), .QN(
    UNCONNECTED258), .D(n_11), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[152] (.Q(\dot_product_and_ReLU[9].product_terms[152][0] ), .QN(
    UNCONNECTED259), .D(n_10), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[153] (.Q(\dot_product_and_ReLU[18].product_terms[153][0] ), .QN(
    UNCONNECTED260), .D(n_7), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[154] (.Q(\dot_product_and_ReLU[14].product_terms[154][0] ), .QN(
    UNCONNECTED261), .D(n_6), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[155] (.Q(\dot_product_and_ReLU[0].product_terms[155][0] ), .QN(
    UNCONNECTED262), .D(n_4), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[156] (.Q(\dot_product_and_ReLU[17].product_terms[156][2] ), .QN(
    UNCONNECTED263), .D(n_3), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[157] (.Q(\dot_product_and_ReLU[0].product_terms[157][0] ), .QN(
    UNCONNECTED264), .D(n_1), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[158] (.Q(\dot_product_and_ReLU[1].product_terms[158][0] ), .QN(
    UNCONNECTED265), .D(n_0), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[159] (.Q(\dot_product_and_ReLU[0].product_terms[159][1] ), .QN(
    UNCONNECTED266), .D(n_237), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[160] (.Q(\dot_product_and_ReLU[5].product_terms[160][1] ), .QN(
    UNCONNECTED267), .D(n_236), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[161] (.Q(\dot_product_and_ReLU[3].product_terms[161][0] ), .QN(
    UNCONNECTED268), .D(n_235), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[162] (.Q(\level_1_sums[1][81][0] ), .QN(UNCONNECTED269), .D(
    n_234), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[163] (.Q(\dot_product_and_ReLU[9].product_terms[163][0] ), .QN(
    UNCONNECTED270), .D(n_233), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[164] (.Q(\dot_product_and_ReLU[3].product_terms[164][0] ), .QN(
    UNCONNECTED271), .D(n_231), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[165] (.Q(\dot_product_and_ReLU[2].product_terms[165][0] ), .QN(
    UNCONNECTED272), .D(n_228), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[166] (.Q(\dot_product_and_ReLU[4].product_terms[166][0] ), .QN(
    UNCONNECTED273), .D(n_227), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[167] (.Q(\dot_product_and_ReLU[0].product_terms[167][0] ), .QN(
    UNCONNECTED274), .D(n_226), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[168] (.Q(\dot_product_and_ReLU[3].product_terms[168][0] ), .QN(
    UNCONNECTED275), .D(n_225), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[169] (.Q(\dot_product_and_ReLU[0].product_terms[169][0] ), .QN(
    UNCONNECTED276), .D(n_222), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[170] (.Q(\dot_product_and_ReLU[1].product_terms[170][0] ), .QN(
    UNCONNECTED277), .D(n_221), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[171] (.Q(\dot_product_and_ReLU[1].product_terms[171][1] ), .QN(
    UNCONNECTED278), .D(n_219), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[172] (.Q(\dot_product_and_ReLU[10].product_terms[172][1] ), .QN(
    UNCONNECTED279), .D(n_218), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[174] (.Q(\dot_product_and_ReLU[2].product_terms[174][1] ), .QN(
    UNCONNECTED280), .D(n_217), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[175] (.Q(\dot_product_and_ReLU[2].product_terms[175][0] ), .QN(
    UNCONNECTED281), .D(n_216), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[176] (.Q(\dot_product_and_ReLU[1].product_terms[176][0] ), .QN(
    UNCONNECTED282), .D(n_214), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[177] (.Q(\dot_product_and_ReLU[0].product_terms[177][0] ), .QN(
    UNCONNECTED283), .D(n_212), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[178] (.Q(\dot_product_and_ReLU[3].product_terms[178][0] ), .QN(
    UNCONNECTED284), .D(n_211), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[179] (.Q(\dot_product_and_ReLU[0].product_terms[179][0] ), .QN(
    UNCONNECTED285), .D(n_209), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[180] (.Q(\dot_product_and_ReLU[8].product_terms[180][0] ), .QN(
    UNCONNECTED286), .D(n_208), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[182] (.Q(\dot_product_and_ReLU[8].product_terms[182][0] ), .QN(
    UNCONNECTED287), .D(n_205), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[183] (.Q(\dot_product_and_ReLU[18].product_terms[183][1] ), .QN(
    UNCONNECTED288), .D(n_203), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[184] (.Q(\dot_product_and_ReLU[3].product_terms[184][1] ), .QN(
    UNCONNECTED289), .D(n_202), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[185] (.Q(\dot_product_and_ReLU[5].product_terms[185][0] ), .QN(
    UNCONNECTED290), .D(n_199), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[186] (.Q(\dot_product_and_ReLU[18].product_terms[186][0] ), .QN(
    UNCONNECTED291), .D(n_198), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[187] (.Q(\dot_product_and_ReLU[0].product_terms[187][0] ), .QN(
    UNCONNECTED292), .D(n_196), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[188] (.Q(\dot_product_and_ReLU[6].product_terms[188][1] ), .QN(
    UNCONNECTED293), .D(n_195), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[189] (.Q(\dot_product_and_ReLU[0].product_terms[189][0] ), .QN(
    UNCONNECTED294), .D(n_193), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[190] (.Q(\dot_product_and_ReLU[4].product_terms[190][1] ), .QN(
    UNCONNECTED295), .D(n_192), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[191] (.Q(\dot_product_and_ReLU[0].product_terms[191][1] ), .QN(
    UNCONNECTED296), .D(n_191), .RN(rst_n), .CK(clk));
  DFFRX2 \B_reg[192] (.Q(B[192]), .QN(UNCONNECTED297), .D(n_189), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[193] (.Q(B[193]), .QN(UNCONNECTED298), .D(n_188), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[195] (.Q(B[195]), .QN(UNCONNECTED299), .D(n_186), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[196] (.Q(B[196]), .QN(UNCONNECTED300), .D(n_185), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[197] (.Q(B[197]), .QN(UNCONNECTED301), .D(n_182), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[198] (.Q(B[198]), .QN(UNCONNECTED302), .D(n_181), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[199] (.Q(B[199]), .QN(UNCONNECTED303), .D(n_180), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[200] (.Q(B[200]), .QN(UNCONNECTED304), .D(n_179), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[201] (.Q(B[201]), .QN(UNCONNECTED305), .D(n_176), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[202] (.Q(B[202]), .QN(UNCONNECTED306), .D(n_175), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[203] (.Q(B[203]), .QN(UNCONNECTED307), .D(n_173), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[204] (.Q(B[204]), .QN(UNCONNECTED308), .D(n_172), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[205] (.Q(B[205]), .QN(UNCONNECTED309), .D(n_170), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[206] (.Q(B[206]), .QN(UNCONNECTED310), .D(n_169), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[207] (.Q(B[207]), .QN(UNCONNECTED311), .D(n_168), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[208] (.Q(B[208]), .QN(UNCONNECTED312), .D(n_166), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[209] (.Q(B[209]), .QN(UNCONNECTED313), .D(n_164), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[210] (.Q(B[210]), .QN(UNCONNECTED314), .D(n_163), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[211] (.Q(B[211]), .QN(UNCONNECTED315), .D(n_161), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[212] (.Q(B[212]), .QN(UNCONNECTED316), .D(n_160), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[213] (.Q(B[213]), .QN(UNCONNECTED317), .D(n_157), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[214] (.Q(B[214]), .QN(UNCONNECTED318), .D(n_156), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[215] (.Q(B[215]), .QN(UNCONNECTED319), .D(n_154), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[216] (.Q(B[216]), .QN(UNCONNECTED320), .D(n_153), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[217] (.Q(B[217]), .QN(UNCONNECTED321), .D(n_151), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[218] (.Q(B[218]), .QN(UNCONNECTED322), .D(n_150), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[219] (.Q(B[219]), .QN(UNCONNECTED323), .D(n_148), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[220] (.Q(B[220]), .QN(UNCONNECTED324), .D(n_147), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[221] (.Q(B[221]), .QN(UNCONNECTED325), .D(n_145), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[222] (.Q(B[222]), .QN(UNCONNECTED326), .D(n_144), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[223] (.Q(B[223]), .QN(UNCONNECTED327), .D(n_143), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[224] (.Q(B[224]), .QN(UNCONNECTED328), .D(n_142), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[225] (.Q(B[225]), .QN(UNCONNECTED329), .D(n_141), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[226] (.Q(B[226]), .QN(UNCONNECTED330), .D(n_140), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[227] (.Q(B[227]), .QN(UNCONNECTED331), .D(n_139), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[228] (.Q(B[228]), .QN(UNCONNECTED332), .D(n_137), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[229] (.Q(B[229]), .QN(UNCONNECTED333), .D(n_134), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[230] (.Q(B[230]), .QN(UNCONNECTED334), .D(n_133), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[231] (.Q(B[231]), .QN(UNCONNECTED335), .D(n_132), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[233] (.Q(B[233]), .QN(UNCONNECTED336), .D(n_155), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[234] (.Q(B[234]), .QN(UNCONNECTED337), .D(n_129), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[235] (.Q(B[235]), .QN(UNCONNECTED338), .D(n_127), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[236] (.Q(B[236]), .QN(UNCONNECTED339), .D(n_126), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[237] (.Q(B[237]), .QN(UNCONNECTED340), .D(n_159), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[238] (.Q(B[238]), .QN(UNCONNECTED341), .D(n_124), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[239] (.Q(B[239]), .QN(UNCONNECTED342), .D(n_123), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[240] (.Q(B[240]), .QN(UNCONNECTED343), .D(n_122), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[241] (.Q(B[241]), .QN(UNCONNECTED344), .D(n_238), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[242] (.Q(B[242]), .QN(UNCONNECTED345), .D(n_59), .RN(rst_n), .CK(
    clk));
  DFFRX2 \B_reg[243] (.Q(B[243]), .QN(UNCONNECTED346), .D(n_117), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[244] (.Q(B[244]), .QN(UNCONNECTED347), .D(n_116), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[245] (.Q(B[245]), .QN(UNCONNECTED348), .D(n_204), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[246] (.Q(B[246]), .QN(UNCONNECTED349), .D(n_115), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[247] (.Q(B[247]), .QN(UNCONNECTED350), .D(n_114), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[248] (.Q(B[248]), .QN(UNCONNECTED351), .D(n_113), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[249] (.Q(B[249]), .QN(UNCONNECTED352), .D(n_207), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[250] (.Q(B[250]), .QN(UNCONNECTED353), .D(n_110), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[251] (.Q(B[251]), .QN(UNCONNECTED354), .D(n_108), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[252] (.Q(B[252]), .QN(UNCONNECTED355), .D(n_107), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[253] (.Q(B[253]), .QN(UNCONNECTED356), .D(n_224), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[254] (.Q(B[254]), .QN(UNCONNECTED357), .D(n_105), .RN(rst_n),
     .CK(clk));
  DFFRX2 \B_reg[255] (.Q(B[255]), .QN(UNCONNECTED358), .D(n_104), .RN(rst_n),
     .CK(clk));
  BUFX8 g21207(.Y(\dot_product_and_ReLU[0].product_terms[13][0] ), .A(n_250));
  BUFX8 g21208(.Y(\dot_product_and_ReLU[0].product_terms[65][0] ), .A(n_249));
  BUFX8 g21209(.Y(\dot_product_and_ReLU[16].product_terms[71][0] ), .A(n_246));
  BUFX8 g21210(.Y(\level_1_sums[4][37][1] ), .A(n_245));
  BUFX8 g21211(.Y(\dot_product_and_ReLU[3].product_terms[84][0] ), .A(n_244));
  BUFX8 g21212(.Y(\dot_product_and_ReLU[0].product_terms[114][1] ), .A(n_243));
  BUFX8 g21213(.Y(\dot_product_and_ReLU[4].product_terms[118][0] ), .A(n_242));
  BUFX8 g21214(.Y(\dot_product_and_ReLU[8].product_terms[173][1] ), .A(n_240));
  BUFX8 g21215(.Y(\dot_product_and_ReLU[3].product_terms[181][0] ), .A(n_239));
endmodule

module csa_tree_ADD_TC_OP_19_group_17897(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_435, n_434, n_431, n_429, n_427, n_425, n_423, n_421, n_419, n_417, 
    n_416, n_415, n_413, n_412, n_411, n_410, n_409, n_408, n_407, n_406, 
    n_405, n_404, n_403, n_401, n_400, n_399, n_398, n_397, n_396, n_395, 
    n_394, n_393, n_392, n_391, n_390, n_389, n_388, n_387, n_386, n_385, 
    n_384, n_383, n_382, n_380, n_379, n_378, n_377, n_376, n_375, n_374, 
    n_373, n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_364, n_363, 
    n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, 
    n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, 
    n_342, n_341, n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, 
    n_332, n_331, n_330, n_329, n_327, n_326, n_325, n_324, n_323, n_322, 
    n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, n_312, 
    n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, 
    n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, 
    n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, n_282, 
    n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, 
    n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, 
    n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, 
    n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, n_242, 
    n_241, n_240, n_239, n_238, n_237, n_236, n_234, n_233, n_232, n_231, 
    n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, 
    n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, 
    n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, 
    n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, 
    n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, 
    n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, 
    n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, 
    n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, 
    n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, 
    n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
    n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = out_0[18];
  AND3XL g14971(.Y(out_0[18]), .A(n_318), .B(n_385), .C(n_435));
  XNOR2X1 g14972(.Y(out_0[15]), .A(n_394), .B(n_434));
  NAND2BX1 g14973(.Y(n_435), .AN(n_384), .B(n_434));
  ADDFX1 g14974(.CO(n_434), .S(out_0[14]), .A(n_378), .B(n_397), .CI(n_431));
  ADDFX1 g14975(.CO(n_431), .S(out_0[13]), .A(n_407), .B(n_398), .CI(n_429));
  ADDFX1 g14976(.CO(n_429), .S(out_0[12]), .A(n_415), .B(n_408), .CI(n_427));
  ADDFX1 g14977(.CO(n_427), .S(out_0[11]), .A(n_409), .B(n_416), .CI(n_425));
  ADDFX1 g14978(.CO(n_425), .S(out_0[10]), .A(n_411), .B(n_410), .CI(n_423));
  ADDFX1 g14979(.CO(n_423), .S(out_0[9]), .A(n_403), .B(n_412), .CI(n_421));
  ADDFX1 g14980(.CO(n_421), .S(out_0[8]), .A(n_405), .B(n_404), .CI(n_419));
  ADDFX1 g14981(.CO(n_419), .S(out_0[7]), .A(n_399), .B(n_406), .CI(n_417));
  ADDFX1 g14982(.CO(n_417), .S(out_0[6]), .A(n_395), .B(n_400), .CI(n_413));
  ADDFX1 g14983(.CO(n_415), .S(n_416), .A(n_392), .B(n_391), .CI(n_363));
  ADDFX1 g14984(.CO(n_413), .S(out_0[5]), .A(n_374), .B(n_396), .CI(n_401));
  ADDFX1 g14985(.CO(n_411), .S(n_412), .A(n_358), .B(n_386), .CI(n_389));
  ADDFX1 g14986(.CO(n_409), .S(n_410), .A(n_388), .B(n_357), .CI(n_393));
  ADDFX1 g14987(.CO(n_407), .S(n_408), .A(n_362), .B(n_390), .CI(n_377));
  ADDFX1 g14988(.CO(n_405), .S(n_406), .A(n_382), .B(n_369), .CI(n_373));
  ADDFX1 g14989(.CO(n_403), .S(n_404), .A(n_359), .B(n_372), .CI(n_387));
  ADDFX1 g14990(.CO(n_401), .S(out_0[4]), .A(n_350), .B(n_380), .CI(n_375));
  ADDFX1 g14991(.CO(n_399), .S(n_400), .A(n_366), .B(n_341), .CI(n_383));
  ADDFX1 g14992(.CO(n_397), .S(n_398), .A(n_352), .B(n_361), .CI(n_376));
  ADDFX1 g14993(.CO(n_395), .S(n_396), .A(n_354), .B(n_343), .CI(n_367));
  NAND2BX1 g14994(.Y(n_394), .AN(n_384), .B(n_385));
  ADDFX1 g14995(.CO(n_392), .S(n_393), .A(n_336), .B(n_370), .CI(n_345));
  ADDFX1 g14996(.CO(n_390), .S(n_391), .A(n_344), .B(n_347), .CI(n_356));
  ADDFX1 g14997(.CO(n_388), .S(n_389), .A(n_337), .B(n_301), .CI(n_371));
  ADDFX1 g14998(.CO(n_386), .S(n_387), .A(n_295), .B(n_349), .CI(n_368));
  NAND2X1 g14999(.Y(n_385), .A(n_331), .B(n_379));
  NOR2X1 g15000(.Y(n_384), .A(n_331), .B(n_379));
  ADDFX1 g15001(.CO(n_382), .S(n_383), .A(n_322), .B(n_342), .CI(n_320));
  ADDFX1 g15002(.CO(n_380), .S(out_0[3]), .A(n_339), .B(n_364), .CI(n_351));
  ADDFX1 g15003(.CO(n_379), .S(n_378), .A(n_332), .B(n_306), .CI(n_360));
  ADDFX1 g15004(.CO(n_376), .S(n_377), .A(n_346), .B(n_305), .CI(n_353));
  ADDFX1 g15005(.CO(n_374), .S(n_375), .A(n_338), .B(n_308), .CI(n_355));
  ADDFX1 g15006(.CO(n_372), .S(n_373), .A(n_303), .B(n_335), .CI(n_340));
  ADDFX1 g15007(.CO(n_370), .S(n_371), .A(n_294), .B(n_314), .CI(n_348));
  ADDFX1 g15008(.CO(n_368), .S(n_369), .A(n_321), .B(n_319), .CI(n_293));
  ADDFX1 g15009(.CO(n_366), .S(n_367), .A(n_312), .B(n_289), .CI(n_307));
  ADDFX1 g15010(.CO(n_364), .S(out_0[2]), .A(n_327), .B(n_261), .CI(n_330));
  ADDFX1 g15011(.CO(n_362), .S(n_363), .A(n_323), .B(n_316), .CI(n_299));
  ADDFX1 g15012(.CO(n_360), .S(n_361), .A(n_285), .B(n_333), .CI(n_304));
  ADDFX1 g15013(.CO(n_358), .S(n_359), .A(n_302), .B(n_281), .CI(n_334));
  ADDFX1 g15014(.CO(n_356), .S(n_357), .A(n_326), .B(n_300), .CI(n_324));
  ADDFX1 g15015(.CO(n_354), .S(n_355), .A(n_275), .B(n_278), .CI(n_310));
  ADDFX1 g15016(.CO(n_352), .S(n_353), .A(n_297), .B(n_315), .CI(n_298));
  ADDFX1 g15017(.CO(n_350), .S(n_351), .A(n_269), .B(n_329), .CI(n_279));
  ADDFX1 g15018(.CO(n_348), .S(n_349), .A(n_287), .B(n_292), .CI(n_267));
  ADDFX1 g15019(.CO(n_346), .S(n_347), .A(n_245), .B(n_264), .CI(n_325));
  ADDFX1 g15020(.CO(n_344), .S(n_345), .A(n_241), .B(n_313), .CI(n_265));
  ADDFX1 g15021(.CO(n_342), .S(n_343), .A(n_233), .B(n_283), .CI(n_309));
  ADDFX1 g15022(.CO(n_340), .S(n_341), .A(n_282), .B(n_311), .CI(n_277));
  ADDFX1 g15023(.CO(n_338), .S(n_339), .A(n_262), .B(n_257), .CI(n_260));
  ADDFX1 g15024(.CO(n_336), .S(n_337), .A(n_280), .B(n_266), .CI(n_291));
  ADDFX1 g15025(.CO(n_334), .S(n_335), .A(n_227), .B(n_276), .CI(n_255));
  ADDFX1 g15026(.CO(n_332), .S(n_333), .A(n_213), .B(n_296), .CI(n_220));
  CLKXOR2X1 g15027(.Y(n_331), .A(n_209), .B(n_317));
  ADDFX1 g15028(.CO(n_329), .S(n_330), .A(n_258), .B(n_263), .CI(n_195));
  ADDFX1 g15029(.CO(n_327), .S(out_0[1]), .A(n_234), .B(n_259), .CI(n_189));
  ADDFX1 g15030(.CO(n_325), .S(n_326), .A(n_236), .B(n_250), .CI(n_273));
  ADDFX1 g15031(.CO(n_323), .S(n_324), .A(n_154), .B(n_167), .CI(n_290));
  ADDFX1 g15032(.CO(n_321), .S(n_322), .A(n_223), .B(n_252), .CI(n_249));
  ADDFX1 g15033(.CO(n_319), .S(n_320), .A(n_232), .B(n_288), .CI(n_247));
  NAND2XL g15034(.Y(n_318), .A(n_209), .B(n_317));
  ADDFX1 g15035(.CO(n_315), .S(n_316), .A(n_240), .B(n_159), .CI(n_271));
  ADDFX1 g15036(.CO(n_313), .S(n_314), .A(n_230), .B(n_185), .CI(n_286));
  ADDFX1 g15037(.CO(n_311), .S(n_312), .A(n_274), .B(n_253), .CI(n_242));
  ADDFX1 g15038(.CO(n_309), .S(n_310), .A(n_256), .B(n_215), .CI(n_217));
  ADDFX1 g15039(.CO(n_307), .S(n_308), .A(n_224), .B(n_268), .CI(n_243));
  ADDFX1 g15040(.CO(n_317), .S(n_306), .A(n_212), .B(n_284), .CI(n_202));
  ADDFX1 g15041(.CO(n_304), .S(n_305), .A(n_239), .B(n_244), .CI(n_221));
  ADDFX1 g15042(.CO(n_302), .S(n_303), .A(n_248), .B(n_187), .CI(n_246));
  ADDFX1 g15043(.CO(n_300), .S(n_301), .A(n_237), .B(n_251), .CI(n_155));
  ADDFX1 g15044(.CO(n_298), .S(n_299), .A(n_272), .B(n_66), .CI(n_163));
  ADDFX1 g15045(.CO(n_296), .S(n_297), .A(n_20), .B(n_158), .CI(n_270));
  ADDFX1 g15046(.CO(n_294), .S(n_295), .A(n_231), .B(n_254), .CI(n_219));
  ADDFX1 g15047(.CO(n_292), .S(n_293), .A(n_222), .B(n_179), .CI(n_197));
  ADDFX1 g15048(.CO(n_290), .S(n_291), .A(n_229), .B(n_218), .CI(n_127));
  ADDFX1 g15049(.CO(n_288), .S(n_289), .A(n_216), .B(n_161), .CI(n_211));
  ADDFX1 g15050(.CO(n_286), .S(n_287), .A(n_207), .B(n_113), .CI(n_178));
  ADDFX1 g15051(.CO(n_284), .S(n_285), .A(n_12), .B(n_238), .CI(n_89));
  ADDFX1 g15052(.CO(n_282), .S(n_283), .A(n_182), .B(n_214), .CI(n_26));
  ADDFX1 g15053(.CO(n_280), .S(n_281), .A(n_186), .B(n_151), .CI(n_226));
  ADDFX1 g15054(.CO(n_278), .S(n_279), .A(n_204), .B(n_194), .CI(n_225));
  ADDFX1 g15055(.CO(n_276), .S(n_277), .A(n_210), .B(n_135), .CI(n_175));
  ADDFX1 g15056(.CO(n_274), .S(n_275), .A(n_180), .B(n_203), .CI(n_183));
  ADDFX1 g15057(.CO(n_272), .S(n_273), .A(n_146), .B(n_228), .CI(in_11[10]));
  ADDFX1 g15058(.CO(n_270), .S(n_271), .A(n_44), .B(n_114), .CI(n_205));
  ADDFX1 g15059(.CO(n_268), .S(n_269), .A(n_200), .B(n_198), .CI(n_181));
  ADDFX1 g15060(.CO(n_266), .S(n_267), .A(n_193), .B(n_196), .CI(n_169));
  ADDFX1 g15061(.CO(n_264), .S(n_265), .A(n_206), .B(n_115), .CI(n_145));
  ADDFX1 g15062(.CO(n_262), .S(n_263), .A(n_172), .B(n_177), .CI(n_190));
  ADDFX1 g15063(.CO(n_260), .S(n_261), .A(n_188), .B(n_201), .CI(n_199));
  ADDFX1 g15064(.CO(n_258), .S(n_259), .A(n_152), .B(n_173), .CI(n_191));
  ADDFX1 g15065(.CO(n_256), .S(n_257), .A(n_176), .B(n_42), .CI(n_74));
  ADDFX1 g15066(.CO(n_254), .S(n_255), .A(n_174), .B(n_208), .CI(n_133));
  ADDFX1 g15067(.CO(n_252), .S(n_253), .A(n_156), .B(n_96), .CI(n_40));
  ADDFX1 g15068(.CO(n_250), .S(n_251), .A(n_147), .B(n_168), .CI(n_150));
  ADDFX1 g15069(.CO(n_248), .S(n_249), .A(n_139), .B(n_25), .CI(n_164));
  ADDFX1 g15070(.CO(n_246), .S(n_247), .A(n_160), .B(n_50), .CI(n_141));
  ADDFX1 g15071(.CO(n_244), .S(n_245), .A(n_149), .B(n_144), .CI(n_166));
  ADDFX1 g15072(.CO(n_242), .S(n_243), .A(n_143), .B(n_157), .CI(n_97));
  ADDFX1 g15073(.CO(n_240), .S(n_241), .A(n_56), .B(n_126), .CI(n_184));
  ADDFX1 g15074(.CO(n_238), .S(n_239), .A(n_148), .B(n_43), .CI(n_14));
  ADDFX1 g15075(.CO(n_236), .S(n_237), .A(n_192), .B(in_1[9]), .CI(n_46));
  ADDFX1 g15076(.CO(n_234), .S(out_0[0]), .A(n_119), .B(n_48), .CI(n_153));
  ADDFX1 g15077(.CO(n_232), .S(n_233), .A(n_142), .B(n_137), .CI(n_165));
  ADDFX1 g15078(.CO(n_230), .S(n_231), .A(n_110), .B(n_68), .CI(n_132));
  ADDFX1 g15079(.CO(n_228), .S(n_229), .A(n_24), .B(n_130), .CI(in_5[9]));
  ADDFX1 g15080(.CO(n_226), .S(n_227), .A(n_140), .B(n_111), .CI(n_134));
  ADDFX1 g15081(.CO(n_224), .S(n_225), .A(n_123), .B(n_80), .CI(n_171));
  ADDFX1 g15082(.CO(n_222), .S(n_223), .A(n_136), .B(n_38), .CI(n_39));
  ADDFX1 g15083(.CO(n_220), .S(n_221), .A(n_85), .B(n_65), .CI(n_162));
  ADDFX1 g15084(.CO(n_218), .S(n_219), .A(n_131), .B(in_11[8]), .CI(in_0[8]));
  ADDFX1 g15085(.CO(n_216), .S(n_217), .A(n_170), .B(n_95), .CI(n_36));
  ADDFX1 g15086(.CO(n_214), .S(n_215), .A(n_122), .B(n_125), .CI(n_73));
  ADDFX1 g15087(.CO(n_212), .S(n_213), .A(n_13), .B(n_129), .CI(n_23));
  ADDFX1 g15088(.CO(n_210), .S(n_211), .A(n_94), .B(n_52), .CI(in_0[5]));
  ADDFX1 g15089(.CO(n_207), .S(n_208), .A(n_100), .B(in_1[7]), .CI(in_7[7]));
  ADDFX1 g15090(.CO(n_205), .S(n_206), .A(n_22), .B(n_107), .CI(in_7[10]));
  ADDFX1 g15091(.CO(n_203), .S(n_204), .A(n_78), .B(n_69), .CI(n_61));
  ADDFX1 g15092(.CO(n_209), .S(n_202), .A(n_128), .B(n_9), .CI(n_88));
  ADDFX1 g15093(.CO(n_200), .S(n_201), .A(n_28), .B(n_31), .CI(n_116));
  ADDFX1 g15094(.CO(n_198), .S(n_199), .A(n_84), .B(n_64), .CI(n_62));
  ADDFX1 g15095(.CO(n_196), .S(n_197), .A(n_37), .B(n_138), .CI(in_0[7]));
  ADDFX1 g15096(.CO(n_194), .S(n_195), .A(n_108), .B(n_58), .CI(n_70));
  ADDFX1 g15097(.CO(n_192), .S(n_193), .A(in_16[8]), .B(n_104), .CI(in_4[8]));
  ADDFX1 g15098(.CO(n_190), .S(n_191), .A(n_118), .B(n_121), .CI(n_60));
  ADDFX1 g15099(.CO(n_188), .S(n_189), .A(n_32), .B(n_109), .CI(n_117));
  ADDFX1 g15100(.CO(n_186), .S(n_187), .A(n_105), .B(n_99), .CI(n_49));
  ADDFX1 g15101(.CO(n_184), .S(n_185), .A(n_103), .B(n_67), .CI(in_15[9]));
  ADDFX1 g15102(.CO(n_182), .S(n_183), .A(n_77), .B(n_41), .CI(n_79));
  ADDFX1 g15103(.CO(n_180), .S(n_181), .A(n_30), .B(n_63), .CI(n_57));
  ADDFX1 g15104(.CO(n_178), .S(n_179), .A(n_87), .B(in_17[7]), .CI(in_11[7]));
  ADDFX1 g15105(.CO(n_176), .S(n_177), .A(n_18), .B(n_120), .CI(n_59));
  ADDFX1 g15106(.CO(n_174), .S(n_175), .A(n_51), .B(n_101), .CI(in_0[6]));
  ADDFX1 g15107(.CO(n_172), .S(n_173), .A(n_19), .B(n_47), .CI(n_81));
  ADDFX1 g15108(.CO(n_170), .S(n_171), .A(n_27), .B(n_83), .CI(in_0[3]));
  ADDFX1 g15109(.CO(n_168), .S(n_169), .A(n_86), .B(n_98), .CI(in_7[8]));
  ADDFX1 g15110(.CO(n_166), .S(n_167), .A(n_34), .B(n_45), .CI(in_0[10]));
  ADDFX1 g15111(.CO(n_164), .S(n_165), .A(n_8), .B(n_124), .CI(in_7[5]));
  ADDFX1 g15112(.CO(n_162), .S(n_163), .A(n_55), .B(in_0[11]), .CI(in_11[11]));
  ADDFX1 g15113(.CO(n_160), .S(n_161), .A(n_72), .B(n_35), .CI(in_11[5]));
  ADDFX1 g15114(.CO(n_158), .S(n_159), .A(n_33), .B(in_15[11]), .CI(in_1[11]));
  ADDFX1 g15115(.CO(n_156), .S(n_157), .A(n_29), .B(in_15[4]), .CI(in_17[4]));
  ADDFX1 g15116(.CO(n_154), .S(n_155), .A(n_112), .B(in_11[9]), .CI(in_0[9]));
  ADDFX1 g15117(.CO(n_152), .S(n_153), .A(in_10[0]), .B(n_11), .CI(n_82));
  ADDFX1 g15118(.CO(n_150), .S(n_151), .A(n_93), .B(in_15[8]), .CI(in_1[8]));
  ADDHX1 g15119(.CO(n_148), .S(n_149), .A(in_4[11]), .B(n_106));
  ADDFX1 g15120(.CO(n_146), .S(n_147), .A(n_92), .B(in_3[9]), .CI(in_4[9]));
  ADDFX1 g15121(.CO(n_144), .S(n_145), .A(n_102), .B(in_1[10]), .CI(in_15[10]));
  ADDFX1 g15122(.CO(n_142), .S(n_143), .A(n_76), .B(in_1[4]), .CI(in_7[4]));
  ADDFX1 g15123(.CO(n_140), .S(n_141), .A(n_54), .B(in_14[6]), .CI(in_15[6]));
  ADDFX1 g15124(.CO(n_138), .S(n_139), .A(n_7), .B(in_16[6]), .CI(in_2[6]));
  ADDFX1 g15125(.CO(n_136), .S(n_137), .A(n_75), .B(in_19[5]), .CI(in_5[5]));
  ADDFX1 g15126(.CO(n_134), .S(n_135), .A(n_71), .B(in_1[6]), .CI(in_11[6]));
  ADDFX1 g15127(.CO(n_132), .S(n_133), .A(n_53), .B(in_5[7]), .CI(in_15[7]));
  ADDFX1 g15128(.CO(n_130), .S(n_131), .A(n_16), .B(in_18[8]), .CI(in_12[8]));
  INVX1 g15129(.Y(n_129), .A(n_91));
  INVX1 g15130(.Y(n_128), .A(n_90));
  ADDFX1 g15131(.CO(n_126), .S(n_127), .A(in_16[9]), .B(in_17[9]), .CI(in_7[9]));
  ADDFX1 g15132(.CO(n_124), .S(n_125), .A(in_18[4]), .B(in_12[4]), .CI(in_3[4]));
  ADDFX1 g15133(.CO(n_122), .S(n_123), .A(in_12[3]), .B(in_7[3]), .CI(in_17[3]));
  ADDFX1 g15134(.CO(n_120), .S(n_121), .A(in_10[1]), .B(in_16[1]), .CI(in_6[1]));
  ADDFX1 g15135(.CO(n_118), .S(n_119), .A(in_1[0]), .B(in_14[0]), .CI(in_17[0]));
  ADDFX1 g15136(.CO(n_116), .S(n_117), .A(in_11[1]), .B(in_15[1]), .CI(in_14[1]));
  ADDFX1 g15137(.CO(n_114), .S(n_115), .A(in_5[10]), .B(in_4[10]), .CI(in_17[10]));
  ADDFX1 g15138(.CO(n_112), .S(n_113), .A(in_2[8]), .B(in_5[8]), .CI(in_17[8]));
  ADDFX1 g15139(.CO(n_110), .S(n_111), .A(in_6[7]), .B(in_2[7]), .CI(in_14[7]));
  ADDFX1 g15140(.CO(n_108), .S(n_109), .A(n_10), .B(in_0[1]), .CI(in_2[1]));
  ADDFX1 g15141(.CO(n_106), .S(n_107), .A(in_13[10]), .B(in_13[9]), .CI(
    in_18[10]));
  ADDFX1 g15142(.CO(n_104), .S(n_105), .A(in_10[7]), .B(n_17), .CI(in_12[7]));
  ADDFX1 g15143(.CO(n_102), .S(n_103), .A(in_12[9]), .B(n_3), .CI(in_18[9]));
  ADDFX1 g15144(.CO(n_100), .S(n_101), .A(n_2), .B(in_3[6]), .CI(in_19[6]));
  ADDFX1 g15145(.CO(n_98), .S(n_99), .A(in_19[7]), .B(in_4[7]), .CI(in_16[7]));
  ADDFX1 g15146(.CO(n_96), .S(n_97), .A(in_5[4]), .B(in_0[4]), .CI(in_11[4]));
  ADDFX1 g15147(.CO(n_94), .S(n_95), .A(in_16[4]), .B(in_19[4]), .CI(in_2[4]));
  ADDFX1 g15148(.CO(n_92), .S(n_93), .A(in_10[8]), .B(n_15), .CI(in_6[8]));
  ADDFX1 g15149(.CO(n_90), .S(n_91), .A(in_7[12]), .B(in_11[12]), .CI(in_17[13]));
  INVX1 g15150(.Y(n_89), .A(n_88));
  ADDFX1 g15151(.CO(n_86), .S(n_87), .A(in_10[6]), .B(in_18[7]), .CI(in_3[7]));
  ADDFX1 g15152(.CO(n_88), .S(n_85), .A(n_5), .B(in_7[12]), .CI(in_17[12]));
  ADDFX1 g15153(.CO(n_83), .S(n_84), .A(in_3[2]), .B(in_16[2]), .CI(in_13[2]));
  ADDFX1 g15154(.CO(n_81), .S(n_82), .A(in_11[0]), .B(in_5[0]), .CI(in_16[0]));
  ADDFX1 g15155(.CO(n_79), .S(n_80), .A(in_2[3]), .B(in_19[3]), .CI(in_15[3]));
  ADDFX1 g15156(.CO(n_77), .S(n_78), .A(in_18[3]), .B(in_3[3]), .CI(in_4[3]));
  ADDFX1 g15157(.CO(n_75), .S(n_76), .A(in_9[4]), .B(in_10[4]), .CI(in_13[4]));
  ADDFX1 g15158(.CO(n_73), .S(n_74), .A(in_1[3]), .B(in_14[3]), .CI(in_11[3]));
  ADDFX1 g15159(.CO(n_71), .S(n_72), .A(in_9[5]), .B(in_18[5]), .CI(in_6[5]));
  ADDFX1 g15160(.CO(n_69), .S(n_70), .A(in_1[2]), .B(in_2[2]), .CI(in_11[2]));
  ADDFX1 g15161(.CO(n_67), .S(n_68), .A(in_14[8]), .B(in_3[8]), .CI(in_19[8]));
  ADDFX1 g15162(.CO(n_65), .S(n_66), .A(n_4), .B(in_7[11]), .CI(in_17[11]));
  ADDFX1 g15163(.CO(n_63), .S(n_64), .A(in_9[2]), .B(in_6[2]), .CI(in_7[2]));
  ADDFX1 g15164(.CO(n_61), .S(n_62), .A(in_15[2]), .B(in_19[2]), .CI(in_0[2]));
  ADDFX1 g15165(.CO(n_59), .S(n_60), .A(in_9[1]), .B(in_19[1]), .CI(in_3[1]));
  ADDFX1 g15166(.CO(n_57), .S(n_58), .A(in_5[2]), .B(in_17[2]), .CI(in_14[2]));
  ADDFX1 g15167(.CO(n_55), .S(n_56), .A(in_19[10]), .B(in_3[10]), .CI(in_16[10]));
  ADDFX1 g15168(.CO(n_53), .S(n_54), .A(in_9[6]), .B(in_13[6]), .CI(in_12[6]));
  ADDFX1 g15169(.CO(n_51), .S(n_52), .A(in_16[5]), .B(in_12[5]), .CI(in_3[5]));
  ADDFX1 g15170(.CO(n_49), .S(n_50), .A(in_6[6]), .B(in_7[6]), .CI(in_17[6]));
  ADDFX1 g15171(.CO(n_47), .S(n_48), .A(in_7[0]), .B(n_0), .CI(in_15[0]));
  ADDFX1 g15172(.CO(n_45), .S(n_46), .A(in_6[9]), .B(in_19[9]), .CI(in_2[9]));
  ADDFX1 g15173(.CO(n_43), .S(n_44), .A(in_3[11]), .B(in_18[11]), .CI(in_16[11]));
  ADDFX1 g15174(.CO(n_41), .S(n_42), .A(in_16[3]), .B(in_6[3]), .CI(in_5[3]));
  ADDFX1 g15175(.CO(n_39), .S(n_40), .A(in_4[5]), .B(in_2[5]), .CI(in_14[5]));
  ADDFX1 g15176(.CO(n_37), .S(n_38), .A(in_18[6]), .B(in_4[6]), .CI(in_5[6]));
  ADDFX1 g15177(.CO(n_35), .S(n_36), .A(in_4[4]), .B(in_6[4]), .CI(in_14[4]));
  ADDFX1 g15178(.CO(n_33), .S(n_34), .A(in_12[10]), .B(n_1), .CI(in_2[10]));
  ADDFX1 g15179(.CO(n_31), .S(n_32), .A(in_1[1]), .B(in_7[1]), .CI(in_17[1]));
  ADDFX1 g15180(.CO(n_29), .S(n_30), .A(in_9[3]), .B(in_10[3]), .CI(in_13[3]));
  ADDFX1 g15181(.CO(n_27), .S(n_28), .A(in_4[2]), .B(in_10[2]), .CI(in_12[2]));
  ADDFX1 g15182(.CO(n_25), .S(n_26), .A(in_15[5]), .B(in_1[5]), .CI(in_17[5]));
  XNOR2X1 g15183(.Y(n_24), .A(in_13[9]), .B(n_21));
  XNOR2X1 g15184(.Y(n_23), .A(in_1[12]), .B(n_20));
  NOR2BX1 g15185(.Y(n_22), .AN(n_21), .B(in_13[9]));
  ADDHX1 g15186(.CO(n_18), .S(n_19), .A(in_4[1]), .B(in_5[1]));
  ADDHX1 g15187(.CO(n_16), .S(n_17), .A(in_9[7]), .B(in_13[7]));
  ADDHX1 g15188(.CO(n_21), .S(n_15), .A(in_9[8]), .B(in_13[8]));
  ADDHX1 g15189(.CO(n_13), .S(n_14), .A(in_1[12]), .B(in_11[12]));
  ADDHX1 g15190(.CO(n_12), .S(n_20), .A(in_15[12]), .B(in_0[11]));
  ADDHX1 g15191(.CO(n_10), .S(n_11), .A(in_0[0]), .B(in_4[0]));
  OAI22X1 g15192(.Y(n_9), .A0(in_15[12]), .A1(n_6), .B0(in_1[12]), .B1(in_0[11]));
  OAI2BB1X1 g15193(.Y(n_8), .A0N(in_10[5]), .A1N(in_13[5]), .B0(n_7));
  OR2X1 g15194(.Y(n_7), .A(in_10[5]), .B(in_13[5]));
  AND2XL g15195(.Y(n_6), .A(in_1[12]), .B(in_0[11]));
  INVX1 g15196(.Y(n_5), .A(in_18[11]));
  INVX1 g15197(.Y(n_4), .A(in_12[10]));
  INVX1 g15198(.Y(n_3), .A(in_14[8]));
  INVX1 g15199(.Y(n_2), .A(in_10[6]));
  INVX1 g15200(.Y(n_1), .A(in_6[9]));
  BUFX2 drc_bufs(.Y(n_0), .A(in_2[0]));
endmodule

module csa_tree_ADD_TC_OP_19_group_8228_1(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_352, n_350, n_348, n_346, n_344, n_342, n_340, n_338, n_336, n_334, 
    n_333, n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, 
    n_322, n_321, n_320, n_319, n_318, n_316, n_315, n_314, n_313, n_312, 
    n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, 
    n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, 
    n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, n_282, 
    n_281, n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, 
    n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, 
    n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, 
    n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, 
    n_240, n_239, n_238, n_237, n_236, n_234, n_233, n_232, n_231, n_230, 
    n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, 
    n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, 
    n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, 
    n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, 
    n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, 
    n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, 
    n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, 
    n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_150, n_149, 
    n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  assign out_0[14] = 1'b0;
  OR2X1 g4397(.Y(out_0[18]), .A(n_236), .B(n_352));
  AOI222X1 g4398(.Y(n_352), .A0(n_108), .A1(n_232), .B0(n_301), .B1(n_350), .C0(
    n_233), .C1(n_300));
  ADDFX1 g4399(.CO(n_350), .S(out_0[13]), .A(n_299), .B(n_318), .CI(n_348));
  ADDFX1 g4400(.CO(n_348), .S(out_0[12]), .A(n_326), .B(n_319), .CI(n_346));
  ADDFX1 g4401(.CO(n_346), .S(out_0[11]), .A(n_332), .B(n_327), .CI(n_344));
  ADDFX1 g4402(.CO(n_344), .S(out_0[10]), .A(n_330), .B(n_333), .CI(n_342));
  ADDFX1 g4403(.CO(n_342), .S(out_0[9]), .A(n_328), .B(n_331), .CI(n_340));
  ADDFX1 g4404(.CO(n_340), .S(out_0[8]), .A(n_324), .B(n_329), .CI(n_338));
  ADDFX1 g4405(.CO(n_338), .S(out_0[7]), .A(n_320), .B(n_325), .CI(n_336));
  ADDFX1 g4406(.CO(n_336), .S(out_0[6]), .A(n_312), .B(n_334), .CI(n_321));
  ADDFX1 g4407(.CO(n_334), .S(out_0[5]), .A(n_297), .B(n_313), .CI(n_322));
  ADDFX1 g4408(.CO(n_332), .S(n_333), .A(n_292), .B(n_314), .CI(n_305));
  ADDFX1 g4409(.CO(n_330), .S(n_331), .A(n_295), .B(n_310), .CI(n_315));
  ADDFX1 g4410(.CO(n_328), .S(n_329), .A(n_296), .B(n_308), .CI(n_311));
  ADDFX1 g4411(.CO(n_326), .S(n_327), .A(n_286), .B(n_304), .CI(n_307));
  ADDFX1 g4412(.CO(n_324), .S(n_325), .A(n_302), .B(n_290), .CI(n_309));
  ADDFX1 g4413(.CO(n_322), .S(out_0[4]), .A(n_275), .B(n_316), .CI(n_298));
  ADDFX1 g4414(.CO(n_320), .S(n_321), .A(n_293), .B(n_284), .CI(n_303));
  ADDFX1 g4415(.CO(n_318), .S(n_319), .A(n_285), .B(n_306), .CI(n_282));
  ADDFX1 g4416(.CO(n_316), .S(out_0[3]), .A(n_279), .B(n_254), .CI(n_276));
  ADDFX1 g4417(.CO(n_314), .S(n_315), .A(n_265), .B(n_258), .CI(n_288));
  ADDFX1 g4418(.CO(n_312), .S(n_313), .A(n_277), .B(n_272), .CI(n_294));
  ADDFX1 g4419(.CO(n_310), .S(n_311), .A(n_262), .B(n_289), .CI(n_266));
  ADDFX1 g4420(.CO(n_308), .S(n_309), .A(n_273), .B(n_283), .CI(n_270));
  ADDFX1 g4421(.CO(n_306), .S(n_307), .A(n_246), .B(n_267), .CI(n_291));
  ADDFX1 g4422(.CO(n_304), .S(n_305), .A(n_257), .B(n_268), .CI(n_287));
  ADDFX1 g4423(.CO(n_302), .S(n_303), .A(n_271), .B(n_250), .CI(n_274));
  OR2XL g4424(.Y(n_301), .A(n_233), .B(n_300));
  ADDFX1 g4425(.CO(n_300), .S(n_299), .A(n_199), .B(n_208), .CI(n_281));
  ADDFX1 g4426(.CO(n_297), .S(n_298), .A(n_253), .B(n_252), .CI(n_278));
  ADDFX1 g4427(.CO(n_295), .S(n_296), .A(n_263), .B(n_161), .CI(n_269));
  ADDFX1 g4428(.CO(n_293), .S(n_294), .A(n_251), .B(n_240), .CI(n_256));
  ADDFX1 g4429(.CO(n_291), .S(n_292), .A(n_247), .B(n_260), .CI(n_241));
  ADDFX1 g4430(.CO(n_289), .S(n_290), .A(n_249), .B(n_193), .CI(n_264));
  ADDFX1 g4431(.CO(n_287), .S(n_288), .A(n_261), .B(n_248), .CI(n_242));
  ADDFX1 g4432(.CO(n_285), .S(n_286), .A(n_228), .B(n_259), .CI(n_219));
  ADDFX1 g4433(.CO(n_283), .S(n_284), .A(n_239), .B(n_255), .CI(n_231));
  ADDFX1 g4434(.CO(n_281), .S(n_282), .A(n_218), .B(n_209), .CI(n_245));
  ADDFX1 g4435(.CO(n_279), .S(out_0[2]), .A(n_223), .B(n_234), .CI(n_244));
  ADDFX1 g4436(.CO(n_277), .S(n_278), .A(n_224), .B(n_238), .CI(n_221));
  ADDFX1 g4437(.CO(n_275), .S(n_276), .A(n_222), .B(n_217), .CI(n_243));
  ADDFX1 g4438(.CO(n_273), .S(n_274), .A(n_172), .B(n_226), .CI(n_187));
  ADDFX1 g4439(.CO(n_271), .S(n_272), .A(n_237), .B(n_227), .CI(n_173));
  ADDFX1 g4440(.CO(n_269), .S(n_270), .A(n_207), .B(n_230), .CI(n_215));
  ADDFX1 g4441(.CO(n_267), .S(n_268), .A(n_127), .B(n_191), .CI(n_229));
  ADDFX1 g4442(.CO(n_265), .S(n_266), .A(n_213), .B(n_211), .CI(n_192));
  ADDFX1 g4443(.CO(n_263), .S(n_264), .A(n_202), .B(n_186), .CI(n_165));
  ADDFX1 g4444(.CO(n_261), .S(n_262), .A(n_206), .B(n_214), .CI(n_189));
  ADDFX1 g4445(.CO(n_259), .S(n_260), .A(n_105), .B(n_196), .CI(n_204));
  ADDFX1 g4446(.CO(n_257), .S(n_258), .A(n_205), .B(n_197), .CI(n_160));
  ADDFX1 g4447(.CO(n_255), .S(n_256), .A(n_185), .B(n_194), .CI(n_220));
  ADDFX1 g4448(.CO(n_253), .S(n_254), .A(n_200), .B(n_181), .CI(n_225));
  ADDFX1 g4449(.CO(n_251), .S(n_252), .A(n_183), .B(n_216), .CI(n_195));
  ADDFX1 g4450(.CO(n_249), .S(n_250), .A(n_184), .B(n_117), .CI(n_203));
  ADDFX1 g4451(.CO(n_247), .S(n_248), .A(n_63), .B(n_212), .CI(n_188));
  ADDFX1 g4452(.CO(n_245), .S(n_246), .A(n_131), .B(n_190), .CI(n_95));
  ADDFX1 g4453(.CO(n_243), .S(n_244), .A(n_167), .B(n_178), .CI(n_201));
  ADDFX1 g4454(.CO(n_241), .S(n_242), .A(n_210), .B(n_91), .CI(n_163));
  ADDFX1 g4455(.CO(n_239), .S(n_240), .A(n_182), .B(n_37), .CI(n_177));
  ADDFX1 g4456(.CO(n_237), .S(n_238), .A(n_175), .B(n_170), .CI(n_180));
  NOR2XL g4457(.Y(n_236), .A(n_108), .B(n_232));
  ADDFX1 g4458(.CO(n_234), .S(out_0[1]), .A(n_150), .B(n_153), .CI(n_179));
  ADDFX1 g4459(.CO(n_232), .S(n_233), .A(n_109), .B(n_136), .CI(n_198));
  ADDFX1 g4460(.CO(n_230), .S(n_231), .A(n_176), .B(n_93), .CI(n_143));
  ADDFX1 g4461(.CO(n_228), .S(n_229), .A(n_90), .B(n_159), .CI(n_162));
  ADDFX1 g4462(.CO(n_226), .S(n_227), .A(n_174), .B(n_154), .CI(n_139));
  ADDFX1 g4463(.CO(n_224), .S(n_225), .A(n_157), .B(n_166), .CI(n_171));
  ADDFX1 g4464(.CO(n_222), .S(n_223), .A(n_140), .B(n_152), .CI(n_169));
  ADDFX1 g4465(.CO(n_220), .S(n_221), .A(n_77), .B(n_89), .CI(n_155));
  ADDFX1 g4466(.CO(n_218), .S(n_219), .A(n_104), .B(n_158), .CI(n_126));
  ADDFX1 g4467(.CO(n_216), .S(n_217), .A(n_134), .B(n_168), .CI(n_123));
  ADDFX1 g4468(.CO(n_214), .S(n_215), .A(n_149), .B(n_142), .CI(n_116));
  ADDFX1 g4469(.CO(n_212), .S(n_213), .A(n_147), .B(n_112), .CI(in_0[8]));
  ADDFX1 g4470(.CO(n_210), .S(n_211), .A(n_50), .B(n_133), .CI(n_164));
  ADDFX1 g4471(.CO(n_208), .S(n_209), .A(n_130), .B(n_129), .CI(n_94));
  ADDFX1 g4472(.CO(n_206), .S(n_207), .A(in_11[7]), .B(n_144), .CI(n_92));
  ADDFX1 g4473(.CO(n_204), .S(n_205), .A(n_125), .B(n_146), .CI(n_32));
  ADDFX1 g4474(.CO(n_202), .S(n_203), .A(n_42), .B(n_138), .CI(n_102));
  ADDFX1 g4475(.CO(n_200), .S(n_201), .A(n_111), .B(n_35), .CI(n_135));
  ADDFX1 g4476(.CO(n_198), .S(n_199), .A(n_98), .B(n_128), .CI(n_137));
  ADDFX1 g4477(.CO(n_196), .S(n_197), .A(n_72), .B(n_132), .CI(in_0[9]));
  ADDFX1 g4478(.CO(n_194), .S(n_195), .A(n_119), .B(n_122), .CI(n_156));
  ADDFX1 g4479(.CO(n_192), .S(n_193), .A(n_51), .B(n_113), .CI(n_81));
  ADDFX1 g4480(.CO(n_190), .S(n_191), .A(n_124), .B(n_62), .CI(in_1[10]));
  ADDFX1 g4481(.CO(n_188), .S(n_189), .A(n_148), .B(in_5[8]), .CI(in_1[8]));
  ADDFX1 g4482(.CO(n_186), .S(n_187), .A(n_145), .B(n_57), .CI(n_36));
  ADDFX1 g4483(.CO(n_184), .S(n_185), .A(n_39), .B(n_118), .CI(n_76));
  ADDFX1 g4484(.CO(n_182), .S(n_183), .A(n_97), .B(n_86), .CI(n_114));
  ADDFX1 g4485(.CO(n_180), .S(n_181), .A(n_75), .B(n_87), .CI(n_115));
  ADDFX1 g4486(.CO(n_178), .S(n_179), .A(n_41), .B(n_141), .CI(n_53));
  ADDFX1 g4487(.CO(n_176), .S(n_177), .A(n_69), .B(n_96), .CI(in_0[5]));
  ADDFX1 g4488(.CO(n_174), .S(n_175), .A(n_101), .B(n_106), .CI(n_74));
  ADDFX1 g4489(.CO(n_172), .S(n_173), .A(n_43), .B(n_88), .CI(n_103));
  ADDFX1 g4490(.CO(n_170), .S(n_171), .A(n_79), .B(n_107), .CI(n_110));
  ADDFX1 g4491(.CO(n_168), .S(n_169), .A(n_71), .B(n_59), .CI(n_44));
  ADDFX1 g4492(.CO(n_166), .S(n_167), .A(n_82), .B(n_85), .CI(n_52));
  ADDFX1 g4493(.CO(n_164), .S(n_165), .A(n_61), .B(n_56), .CI(in_5[7]));
  ADDFX1 g4494(.CO(n_162), .S(n_163), .A(in_4[9]), .B(n_121), .CI(in_1[9]));
  ADDFX1 g4495(.CO(n_160), .S(n_161), .A(n_73), .B(n_80), .CI(n_33));
  ADDFX1 g4496(.CO(n_158), .S(n_159), .A(in_4[10]), .B(in_8[10]), .CI(n_120));
  ADDFX1 g4497(.CO(n_156), .S(n_157), .A(n_84), .B(n_58), .CI(n_34));
  ADDFX1 g4498(.CO(n_154), .S(n_155), .A(n_15), .B(n_78), .CI(in_5[4]));
  ADDFX1 g4499(.CO(n_152), .S(n_153), .A(n_54), .B(n_83), .CI(n_45));
  ADDFX1 g4500(.CO(n_150), .S(out_0[0]), .A(n_18), .B(n_55), .CI(n_49));
  ADDFX1 g4501(.CO(n_148), .S(n_149), .A(n_46), .B(n_64), .CI(in_12[7]));
  ADDFX1 g4502(.CO(n_146), .S(n_147), .A(n_30), .B(n_60), .CI(in_2[8]));
  ADDFX1 g4503(.CO(n_144), .S(n_145), .A(n_38), .B(n_68), .CI(in_2[6]));
  ADDFX1 g4504(.CO(n_142), .S(n_143), .A(n_47), .B(in_3[6]), .CI(in_5[6]));
  ADDFX1 g4505(.CO(n_140), .S(n_141), .A(n_17), .B(n_24), .CI(n_48));
  ADDFX1 g4506(.CO(n_138), .S(n_139), .A(n_10), .B(n_100), .CI(in_2[5]));
  ADDHX1 g4507(.CO(n_136), .S(n_137), .A(n_29), .B(n_28));
  ADDFX1 g4508(.CO(n_134), .S(n_135), .A(n_23), .B(n_40), .CI(in_0[2]));
  ADDFX1 g4509(.CO(n_132), .S(n_133), .A(n_12), .B(n_67), .CI(in_3[8]));
  ADDFX1 g4510(.CO(n_130), .S(n_131), .A(n_14), .B(n_5), .CI(n_9));
  ADDFX1 g4511(.CO(n_128), .S(n_129), .A(n_11), .B(n_21), .CI(n_99));
  ADDFX1 g4512(.CO(n_126), .S(n_127), .A(n_13), .B(in_18[10]), .CI(in_0[10]));
  ADDFX1 g4513(.CO(n_124), .S(n_125), .A(n_8), .B(n_6), .CI(in_17[9]));
  ADDFX1 g4514(.CO(n_122), .S(n_123), .A(n_70), .B(in_4[3]), .CI(in_5[3]));
  ADDFX1 g4515(.CO(n_120), .S(n_121), .A(in_19[9]), .B(n_66), .CI(in_3[8]));
  ADDFX1 g4516(.CO(n_118), .S(n_119), .A(n_19), .B(in_12[4]), .CI(in_4[4]));
  ADDFX1 g4517(.CO(n_116), .S(n_117), .A(n_65), .B(in_0[6]), .CI(in_1[6]));
  ADDFX1 g4518(.CO(n_114), .S(n_115), .A(n_25), .B(in_2[3]), .CI(in_3[3]));
  ADDFX1 g4519(.CO(n_112), .S(n_113), .A(n_31), .B(in_4[7]), .CI(in_2[7]));
  ADDFX1 g4520(.CO(n_110), .S(n_111), .A(n_26), .B(in_4[2]), .CI(in_11[2]));
  OAI2BB1X1 g4521(.Y(n_109), .A0N(n_27), .A1N(n_16), .B0(n_108));
  OR2X1 g4522(.Y(n_108), .A(n_27), .B(n_16));
  ADDFX1 g4523(.CO(n_106), .S(n_107), .A(in_8[3]), .B(in_14[3]), .CI(in_18[3]));
  ADDFX1 g4524(.CO(n_104), .S(n_105), .A(in_12[10]), .B(in_17[10]), .CI(
    in_11[10]));
  ADDFX1 g4525(.CO(n_102), .S(n_103), .A(in_4[5]), .B(in_5[5]), .CI(in_11[5]));
  ADDFX1 g4526(.CO(n_100), .S(n_101), .A(in_6[4]), .B(in_10[4]), .CI(in_19[4]));
  ADDFX1 g4527(.CO(n_98), .S(n_99), .A(in_8[12]), .B(in_0[12]), .CI(n_1));
  ADDFX1 g4528(.CO(n_96), .S(n_97), .A(in_14[4]), .B(in_8[4]), .CI(in_17[4]));
  ADDFX1 g4529(.CO(n_94), .S(n_95), .A(n_22), .B(in_8[11]), .CI(in_0[11]));
  ADDFX1 g4530(.CO(n_92), .S(n_93), .A(in_4[6]), .B(in_11[6]), .CI(in_18[6]));
  ADDFX1 g4531(.CO(n_90), .S(n_91), .A(in_5[9]), .B(in_11[9]), .CI(in_18[9]));
  ADDFX1 g4532(.CO(n_88), .S(n_89), .A(in_11[4]), .B(in_1[4]), .CI(in_0[4]));
  ADDFX1 g4533(.CO(n_86), .S(n_87), .A(n_20), .B(in_0[3]), .CI(in_11[3]));
  ADDFX1 g4534(.CO(n_84), .S(n_85), .A(in_12[2]), .B(in_18[2]), .CI(in_16[2]));
  ADDFX1 g4535(.CO(n_82), .S(n_83), .A(in_5[1]), .B(in_10[1]), .CI(in_4[1]));
  ADDFX1 g4536(.CO(n_80), .S(n_81), .A(in_18[7]), .B(in_0[7]), .CI(in_1[7]));
  ADDFX1 g4537(.CO(n_78), .S(n_79), .A(in_6[3]), .B(in_10[3]), .CI(in_19[3]));
  ADDFX1 g4538(.CO(n_76), .S(n_77), .A(in_2[4]), .B(in_3[4]), .CI(in_18[4]));
  ADDFX1 g4539(.CO(n_74), .S(n_75), .A(in_1[3]), .B(in_12[3]), .CI(in_17[3]));
  ADDFX1 g4540(.CO(n_72), .S(n_73), .A(in_8[8]), .B(in_17[8]), .CI(in_12[8]));
  ADDFX1 g4541(.CO(n_70), .S(n_71), .A(in_1[2]), .B(in_6[2]), .CI(in_14[2]));
  ADDFX1 g4542(.CO(n_68), .S(n_69), .A(in_13[5]), .B(in_10[5]), .CI(in_16[5]));
  ADDFX1 g4543(.CO(n_66), .S(n_67), .A(in_10[8]), .B(in_6[8]), .CI(in_19[8]));
  ADDFX1 g4544(.CO(n_64), .S(n_65), .A(in_10[6]), .B(in_13[6]), .CI(in_16[6]));
  ADDFX1 g4545(.CO(n_62), .S(n_63), .A(in_13[9]), .B(in_8[9]), .CI(in_12[9]));
  ADDFX1 g4546(.CO(n_60), .S(n_61), .A(in_13[7]), .B(in_10[7]), .CI(in_16[7]));
  ADDFX1 g4547(.CO(n_58), .S(n_59), .A(in_8[2]), .B(in_10[2]), .CI(in_19[2]));
  ADDFX1 g4548(.CO(n_56), .S(n_57), .A(in_8[6]), .B(in_12[6]), .CI(in_17[6]));
  ADDFX1 g4549(.CO(n_54), .S(n_55), .A(in_10[0]), .B(in_18[0]), .CI(in_5[0]));
  ADDFX1 g4550(.CO(n_52), .S(n_53), .A(in_11[1]), .B(in_0[1]), .CI(in_3[1]));
  ADDFX1 g4551(.CO(n_50), .S(n_51), .A(in_8[7]), .B(in_17[7]), .CI(in_3[7]));
  ADDFX1 g4552(.CO(n_48), .S(n_49), .A(in_3[0]), .B(in_0[0]), .CI(in_11[0]));
  ADDFX1 g4553(.CO(n_46), .S(n_47), .A(in_6[6]), .B(in_14[6]), .CI(in_19[6]));
  ADDFX1 g4554(.CO(n_44), .S(n_45), .A(in_1[1]), .B(in_14[1]), .CI(in_2[1]));
  ADDFX1 g4555(.CO(n_42), .S(n_43), .A(in_8[5]), .B(in_12[5]), .CI(in_17[5]));
  ADDFX1 g4556(.CO(n_40), .S(n_41), .A(in_16[1]), .B(in_18[1]), .CI(in_12[1]));
  ADDFX1 g4557(.CO(n_38), .S(n_39), .A(in_6[5]), .B(in_14[5]), .CI(in_19[5]));
  ADDFX1 g4558(.CO(n_36), .S(n_37), .A(in_3[5]), .B(in_18[5]), .CI(in_1[5]));
  ADDFX1 g4559(.CO(n_34), .S(n_35), .A(in_5[2]), .B(in_3[2]), .CI(in_2[2]));
  ADDFX1 g4560(.CO(n_32), .S(n_33), .A(in_4[8]), .B(in_11[8]), .CI(in_18[8]));
  ADDFX1 g4561(.CO(n_30), .S(n_31), .A(in_14[7]), .B(in_6[7]), .CI(in_19[7]));
  OAI21X1 g4562(.Y(n_29), .A0(in_8[12]), .A1(n_7), .B0(n_27));
  XNOR2X1 g4563(.Y(n_28), .A(in_0[12]), .B(n_1));
  NAND2X1 g4564(.Y(n_27), .A(in_8[12]), .B(n_7));
  ADDHX1 g4565(.CO(n_25), .S(n_26), .A(in_13[2]), .B(in_17[2]));
  ADDHX1 g4566(.CO(n_23), .S(n_24), .A(in_6[1]), .B(in_13[1]));
  ADDHX1 g4567(.CO(n_21), .S(n_22), .A(in_12[11]), .B(in_18[11]));
  ADDHX1 g4568(.CO(n_19), .S(n_20), .A(in_13[3]), .B(in_16[3]));
  ADDHX1 g4569(.CO(n_17), .S(n_18), .A(n_2), .B(in_14[0]));
  OAI22X1 g4570(.Y(n_16), .A0(in_18[11]), .A1(n_0), .B0(in_1[11]), .B1(in_0[12]));
  OAI2BB1X1 g4571(.Y(n_15), .A0N(in_16[4]), .A1N(in_13[4]), .B0(n_10));
  OAI21X1 g4572(.Y(n_14), .A0(in_5[10]), .A1(n_4), .B0(n_11));
  XNOR2X1 g4573(.Y(n_13), .A(in_5[10]), .B(in_3[8]));
  XNOR2X1 g4574(.Y(n_12), .A(in_16[8]), .B(in_13[8]));
  NAND2X1 g4576(.Y(n_11), .A(in_5[10]), .B(n_4));
  OR2X1 g4577(.Y(n_10), .A(in_16[4]), .B(in_13[4]));
  NOR2BX1 g4579(.Y(n_9), .AN(in_5[10]), .B(in_3[8]));
  OR2X1 g4580(.Y(n_8), .A(in_16[8]), .B(in_13[8]));
  NAND2X1 g4581(.Y(n_7), .A(in_1[11]), .B(in_18[11]));
  INVX1 g4582(.Y(n_6), .A(in_2[9]));
  INVX1 g4583(.Y(n_5), .A(in_17[11]));
  INVX1 g4585(.Y(n_4), .A(in_1[11]));
  BUFX2 drc_bufs(.Y(n_2), .A(in_2[0]));
  MXI2XL g2(.Y(n_1), .A(n_4), .B(in_1[11]), .S0(in_18[11]));
  NOR2BX1 g4589(.Y(n_0), .AN(in_0[12]), .B(n_4));
endmodule

module csa_tree_ADD_TC_OP_19_group_14031(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_363, n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, 
    n_353, n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, 
    n_343, n_342, n_341, n_340, n_339, n_338, n_337, n_336, n_335, n_334, 
    n_333, n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, 
    n_323, n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, 
    n_313, n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, 
    n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, 
    n_293, n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, 
    n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, 
    n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, 
    n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
    n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, 
    n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, 
    n_223, n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, 
    n_213, n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, 
    n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 
    n_193, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, 
    n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, 
    n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, 
    n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, 
    n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, 
    n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
    n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, 
    n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, 
    n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, 
    n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, 
    n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, 
    n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
    n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  ADDFX1 cdnfadd(.CO(n_49), .S(out_0[0]), .A(n_349), .B(n_333), .CI(n_332));
  ADDFX1 cdnfadd1(.CO(n_48), .S(out_0[1]), .A(n_350), .B(n_334), .CI(n_49));
  ADDFX1 cdnfadd2(.CO(n_47), .S(out_0[2]), .A(n_351), .B(n_335), .CI(n_48));
  ADDFX1 cdnfadd3(.CO(n_46), .S(out_0[3]), .A(n_352), .B(n_336), .CI(n_47));
  ADDFX1 cdnfadd4(.CO(n_45), .S(out_0[4]), .A(n_353), .B(n_337), .CI(n_46));
  ADDFX1 cdnfadd5(.CO(n_44), .S(out_0[5]), .A(n_354), .B(n_338), .CI(n_45));
  ADDFX1 cdnfadd6(.CO(n_43), .S(out_0[6]), .A(n_355), .B(n_339), .CI(n_44));
  ADDFX1 cdnfadd7(.CO(n_42), .S(out_0[7]), .A(n_356), .B(n_340), .CI(n_43));
  ADDFX1 cdnfadd8(.CO(n_41), .S(out_0[8]), .A(n_357), .B(n_341), .CI(n_42));
  ADDFX1 cdnfadd9(.CO(n_40), .S(out_0[9]), .A(n_358), .B(n_342), .CI(n_41));
  ADDFX1 cdnfadd10(.CO(n_39), .S(out_0[10]), .A(n_359), .B(n_343), .CI(n_40));
  ADDFX1 cdnfadd11(.CO(n_38), .S(out_0[11]), .A(n_360), .B(n_344), .CI(n_39));
  ADDFX1 cdnfadd12(.CO(n_37), .S(out_0[12]), .A(n_361), .B(n_345), .CI(n_38));
  ADDFX1 cdnfadd13(.CO(n_36), .S(out_0[13]), .A(n_362), .B(n_346), .CI(n_37));
  ADDFX1 cdnfadd14(.CO(n_35), .S(out_0[14]), .A(n_363), .B(n_347), .CI(n_36));
  ADDFX1 cdnfadd15(.CO(n_34), .S(out_0[15]), .A(n_31), .B(n_348), .CI(n_35));
  ADDFX1 cdnfadd_000_0(.CO(n_331), .S(n_332), .A(in_14[0]), .B(in_15[0]), .CI(
    in_1[0]));
  ADDFX1 cdnfadd_000_1(.CO(n_330), .S(n_329), .A(in_16[0]), .B(in_11[0]), .CI(
    in_4[0]));
  ADDFX1 cdnfadd_000_2(.CO(n_328), .S(n_349), .A(in_5[0]), .B(in_19[0]), .CI(
    in_17[0]));
  ADDFX1 cdnfadd_000_3(.CO(n_225), .S(n_333), .A(in_10[0]), .B(n_25), .CI(n_329));
  ADDFX1 cdnfadd_001_0(.CO(n_327), .S(n_326), .A(in_19[1]), .B(in_14[1]), .CI(
    in_10[1]));
  ADDFX1 cdnfadd_001_1(.CO(n_325), .S(n_324), .A(in_11[1]), .B(in_5[1]), .CI(
    in_15[1]));
  ADDFX1 cdnfadd_001_2(.CO(n_323), .S(n_322), .A(in_8[1]), .B(in_7[1]), .CI(
    in_13[1]));
  ADDFX1 cdnfadd_001_3(.CO(n_321), .S(n_320), .A(in_2[1]), .B(in_1[1]), .CI(
    in_12[1]));
  ADDFX1 cdnfadd_001_4(.CO(n_319), .S(n_318), .A(in_4[1]), .B(in_17[1]), .CI(
    in_16[1]));
  ADDFX1 cdnfadd_001_5(.CO(n_223), .S(n_222), .A(n_20), .B(n_330), .CI(n_328));
  ADDFX1 cdnfadd_001_6(.CO(n_221), .S(n_220), .A(n_331), .B(n_322), .CI(n_326));
  ADDFX1 cdnfadd_001_7(.CO(n_219), .S(n_350), .A(n_324), .B(n_318), .CI(n_320));
  ADDFX1 cdnfadd_001_8(.CO(n_149), .S(n_334), .A(n_225), .B(n_222), .CI(n_220));
  ADDFX1 cdnfadd_002_0(.CO(n_317), .S(n_316), .A(in_5[2]), .B(in_3[2]), .CI(
    in_10[2]));
  ADDFX1 cdnfadd_002_1(.CO(n_315), .S(n_314), .A(in_15[2]), .B(in_14[2]), .CI(
    in_4[2]));
  ADDFX1 cdnfadd_002_2(.CO(n_313), .S(n_312), .A(in_17[2]), .B(in_2[2]), .CI(
    in_12[2]));
  ADDFX1 cdnfadd_002_3(.CO(n_311), .S(n_310), .A(in_8[2]), .B(in_7[2]), .CI(
    in_16[2]));
  ADDFX1 cdnfadd_002_4(.CO(n_309), .S(n_308), .A(in_11[2]), .B(in_1[2]), .CI(
    n_23));
  ADDFX1 cdnfadd_002_5(.CO(n_218), .S(n_217), .A(n_323), .B(n_327), .CI(n_325));
  ADDFX1 cdnfadd_002_6(.CO(n_216), .S(n_215), .A(n_314), .B(n_321), .CI(n_316));
  ADDFX1 cdnfadd_002_7(.CO(n_214), .S(n_213), .A(n_319), .B(n_310), .CI(n_312));
  ADDFX1 cdnfadd_002_8(.CO(n_148), .S(n_147), .A(n_223), .B(n_308), .CI(n_217));
  ADDFX1 cdnfadd_002_9(.CO(n_146), .S(n_351), .A(n_221), .B(n_219), .CI(n_215));
  ADDFX1 cdnfadd_002_10(.CO(n_90), .S(n_335), .A(n_213), .B(n_147), .CI(n_149));
  ADDFX1 cdnfadd_003_0(.CO(n_307), .S(n_306), .A(in_5[3]), .B(in_3[3]), .CI(
    in_8[3]));
  ADDFX1 cdnfadd_003_1(.CO(n_305), .S(n_304), .A(in_15[3]), .B(in_10[3]), .CI(
    in_14[3]));
  ADDFX1 cdnfadd_003_2(.CO(n_303), .S(n_302), .A(in_19[3]), .B(in_13[3]), .CI(
    in_2[3]));
  ADDFX1 cdnfadd_003_3(.CO(n_301), .S(n_300), .A(in_11[3]), .B(in_7[3]), .CI(
    n_16));
  ADDFX1 cdnfadd_003_4(.CO(n_299), .S(n_298), .A(in_17[3]), .B(in_12[3]), .CI(
    in_16[3]));
  ADDFX1 cdnfadd_003_5(.CO(n_212), .S(n_211), .A(in_1[3]), .B(in_4[3]), .CI(
    n_317));
  ADDFX1 cdnfadd_003_6(.CO(n_210), .S(n_209), .A(n_306), .B(n_315), .CI(n_313));
  ADDFX1 cdnfadd_003_7(.CO(n_208), .S(n_207), .A(n_311), .B(n_302), .CI(n_304));
  ADDFX1 cdnfadd_003_8(.CO(n_145), .S(n_144), .A(n_309), .B(n_211), .CI(n_218));
  ADDFX1 cdnfadd_003_9(.CO(n_143), .S(n_142), .A(n_300), .B(n_298), .CI(n_216));
  ADDFX1 cdnfadd_003_10(.CO(n_141), .S(n_140), .A(n_209), .B(n_214), .CI(n_207));
  ADDFX1 cdnfadd_003_11(.CO(n_89), .S(n_352), .A(n_142), .B(n_148), .CI(n_144));
  ADDFX1 cdnfadd_003_12(.CO(n_353), .S(n_336), .A(n_146), .B(n_140), .CI(n_90));
  ADDFX1 cdnfadd_004_0(.CO(n_297), .S(n_296), .A(in_17[4]), .B(in_19[4]), .CI(
    in_11[4]));
  ADDFX1 cdnfadd_004_1(.CO(n_295), .S(n_294), .A(in_1[4]), .B(in_7[4]), .CI(
    in_12[4]));
  ADDFX1 cdnfadd_004_2(.CO(n_293), .S(n_292), .A(in_8[4]), .B(in_10[4]), .CI(
    n_27));
  ADDFX1 cdnfadd_004_3(.CO(n_291), .S(n_290), .A(in_14[4]), .B(in_16[4]), .CI(
    in_13[4]));
  ADDFX1 cdnfadd_004_4(.CO(n_289), .S(n_288), .A(in_4[4]), .B(in_15[4]), .CI(
    in_2[4]));
  ADDFX1 cdnfadd_004_5(.CO(n_206), .S(n_200), .A(n_307), .B(n_305), .CI(n_303));
  ADDFX1 cdnfadd_004_6(.CO(n_199), .S(n_198), .A(n_301), .B(n_299), .CI(n_296));
  ADDFX1 cdnfadd_004_7(.CO(n_139), .S(n_138), .A(n_212), .B(n_292), .CI(n_294));
  ADDFX1 cdnfadd_004_8(.CO(n_137), .S(n_136), .A(n_288), .B(n_210), .CI(n_290));
  ADDFX1 cdnfadd_004_9(.CO(n_88), .S(n_87), .A(n_200), .B(n_208), .CI(n_145));
  ADDFX1 cdnfadd_004_10(.CO(n_86), .S(n_85), .A(n_198), .B(n_143), .CI(n_138));
  ADDFX1 cdnfadd_004_11(.CO(n_63), .S(n_62), .A(n_136), .B(n_141), .CI(n_87));
  ADDFX1 cdnfadd_004_12(.CO(n_354), .S(n_337), .A(n_89), .B(n_85), .CI(n_62));
  ADDFX1 cdnfadd_005_0(.CO(n_287), .S(n_286), .A(in_3[5]), .B(n_17), .CI(
    in_10[5]));
  ADDFX1 cdnfadd_005_1(.CO(n_285), .S(n_284), .A(in_19[5]), .B(n_10), .CI(
    in_12[5]));
  ADDFX1 cdnfadd_005_2(.CO(n_283), .S(n_282), .A(in_11[5]), .B(in_8[5]), .CI(
    in_17[5]));
  ADDFX1 cdnfadd_005_3(.CO(n_281), .S(n_280), .A(in_7[5]), .B(in_1[5]), .CI(
    in_14[5]));
  ADDFX1 cdnfadd_005_4(.CO(n_279), .S(n_278), .A(in_15[5]), .B(in_2[5]), .CI(
    in_4[5]));
  ADDFX1 cdnfadd_005_5(.CO(n_197), .S(n_196), .A(in_13[5]), .B(in_16[5]), .CI(
    n_297));
  ADDFX1 cdnfadd_005_6(.CO(n_195), .S(n_194), .A(n_295), .B(n_293), .CI(n_284));
  ADDFX1 cdnfadd_005_7(.CO(n_193), .S(n_192), .A(n_291), .B(n_289), .CI(n_286));
  ADDFX1 cdnfadd_005_8(.CO(n_135), .S(n_134), .A(n_280), .B(n_282), .CI(n_206));
  ADDFX1 cdnfadd_005_9(.CO(n_133), .S(n_132), .A(n_196), .B(n_278), .CI(n_194));
  ADDFX1 cdnfadd_005_10(.CO(n_84), .S(n_83), .A(n_199), .B(n_139), .CI(n_137));
  ADDFX1 cdnfadd_005_11(.CO(n_61), .S(n_60), .A(n_192), .B(n_134), .CI(n_88));
  ADDFX1 cdnfadd_005_12(.CO(n_59), .S(n_58), .A(n_132), .B(n_86), .CI(n_83));
  ADDFX1 cdnfadd_005_13(.CO(n_355), .S(n_338), .A(n_63), .B(n_60), .CI(n_58));
  ADDFX1 cdnfadd_006_1(.CO(n_277), .S(n_276), .A(in_5[5]), .B(in_10[6]), .CI(
    in_12[6]));
  ADDFX1 cdnfadd_006_2(.CO(n_275), .S(n_274), .A(in_19[6]), .B(in_8[6]), .CI(
    in_1[6]));
  ADDFX1 cdnfadd_006_3(.CO(n_273), .S(n_272), .A(in_14[6]), .B(in_17[6]), .CI(
    in_11[6]));
  ADDFX1 cdnfadd_006_4(.CO(n_271), .S(n_270), .A(n_22), .B(in_13[6]), .CI(
    in_4[6]));
  ADDFX1 cdnfadd_006_5(.CO(n_269), .S(n_268), .A(in_16[6]), .B(in_7[6]), .CI(
    in_15[6]));
  ADDFX1 cdnfadd_006_6(.CO(n_191), .S(n_190), .A(in_2[6]), .B(n_287), .CI(n_285));
  ADDFX1 cdnfadd_006_7(.CO(n_187), .S(n_185), .A(n_283), .B(n_281), .CI(n_279));
  ADDFX1 cdnfadd_006_8(.CO(n_184), .S(n_183), .A(n_274), .B(n_276), .CI(n_268));
  ADDFX1 cdnfadd_006_9(.CO(n_131), .S(n_130), .A(n_197), .B(n_272), .CI(n_270));
  ADDFX1 cdnfadd_006_10(.CO(n_129), .S(n_128), .A(n_195), .B(n_190), .CI(n_193));
  ADDFX1 cdnfadd_006_11(.CO(n_82), .S(n_81), .A(n_185), .B(n_135), .CI(n_183));
  ADDFX1 cdnfadd_006_12(.CO(n_113), .S(n_112), .A(n_130), .B(n_133), .CI(n_128));
  ADDFX1 cdnfadd_006_13(.CO(n_51), .S(n_50), .A(n_84), .B(n_81), .CI(n_61));
  ADDFX1 cdnfadd_006_14(.CO(n_356), .S(n_339), .A(n_112), .B(n_59), .CI(n_50));
  ADDFX1 cdnfadd_007_0(.CO(n_267), .S(n_266), .A(n_21), .B(in_8[7]), .CI(n_15));
  ADDFX1 cdnfadd_007_1(.CO(n_265), .S(n_264), .A(in_12[7]), .B(in_17[7]), .CI(
    in_7[7]));
  ADDFX1 cdnfadd_007_2(.CO(n_263), .S(n_262), .A(in_19[7]), .B(in_11[7]), .CI(
    in_10[7]));
  ADDFX1 cdnfadd_007_3(.CO(n_261), .S(n_260), .A(in_15[7]), .B(in_4[7]), .CI(
    in_14[7]));
  ADDFX1 cdnfadd_007_4(.CO(n_259), .S(n_258), .A(in_16[7]), .B(in_1[7]), .CI(
    in_13[7]));
  ADDFX1 cdnfadd_007_5(.CO(n_238), .S(n_237), .A(in_2[7]), .B(n_277), .CI(n_266));
  ADDFX1 cdnfadd_007_6(.CO(n_182), .S(n_181), .A(n_275), .B(n_271), .CI(n_273));
  ADDFX1 cdnfadd_007_7(.CO(n_180), .S(n_179), .A(n_269), .B(n_262), .CI(n_264));
  ADDFX1 cdnfadd_007_8(.CO(n_161), .S(n_160), .A(n_258), .B(n_260), .CI(n_191));
  ADDFX1 cdnfadd_007_9(.CO(n_127), .S(n_126), .A(n_187), .B(n_237), .CI(n_181));
  ADDFX1 cdnfadd_007_10(.CO(n_111), .S(n_110), .A(n_184), .B(n_131), .CI(n_129));
  ADDFX1 cdnfadd_007_11(.CO(n_65), .S(n_64), .A(n_179), .B(n_160), .CI(n_82));
  ADDFX1 cdnfadd_007_12(.CO(n_79), .S(n_78), .A(n_126), .B(n_110), .CI(n_113));
  ADDFX1 cdnfadd_007_13(.CO(n_357), .S(n_340), .A(n_64), .B(n_51), .CI(n_78));
  ADDFX1 cdnfadd_008_1(.CO(n_257), .S(n_256), .A(in_12[8]), .B(n_19), .CI(
    in_8[8]));
  ADDFX1 cdnfadd_008_2(.CO(n_255), .S(n_254), .A(n_9), .B(in_19[8]), .CI(
    in_13[8]));
  ADDFX1 cdnfadd_008_3(.CO(n_253), .S(n_252), .A(in_10[8]), .B(in_17[8]), .CI(
    in_14[8]));
  ADDFX1 cdnfadd_008_4(.CO(n_177), .S(n_176), .A(in_7[8]), .B(in_11[8]), .CI(
    n_256));
  ADDFX1 cdnfadd_008_5(.CO(n_251), .S(n_250), .A(in_4[8]), .B(in_15[8]), .CI(
    in_2[8]));
  ADDFX1 cdnfadd_008_6(.CO(n_236), .S(n_235), .A(in_16[8]), .B(n_267), .CI(
    in_1[8]));
  ADDFX1 cdnfadd_008_7(.CO(n_175), .S(n_174), .A(n_265), .B(n_263), .CI(n_259));
  ADDFX1 cdnfadd_008_8(.CO(n_125), .S(n_124), .A(n_261), .B(n_254), .CI(n_176));
  ADDFX1 cdnfadd_008_9(.CO(n_159), .S(n_158), .A(n_252), .B(n_238), .CI(n_235));
  ADDFX1 cdnfadd_008_10(.CO(n_123), .S(n_122), .A(n_182), .B(n_250), .CI(n_174));
  ADDFX1 cdnfadd_008_11(.CO(n_92), .S(n_91), .A(n_180), .B(n_161), .CI(n_124));
  ADDFX1 cdnfadd_008_12(.CO(n_109), .S(n_108), .A(n_122), .B(n_158), .CI(n_127));
  ADDFX1 cdnfadd_008_13(.CO(n_57), .S(n_56), .A(n_111), .B(n_91), .CI(n_65));
  ADDFX1 cdnfadd_008_14(.CO(n_358), .S(n_341), .A(n_108), .B(n_79), .CI(n_56));
  ADDFX1 cdnfadd_009_0(.CO(n_249), .S(n_248), .A(in_3[9]), .B(in_12[8]), .CI(
    in_8[9]));
  ADDFX1 cdnfadd_009_1(.CO(n_247), .S(n_246), .A(in_3[8]), .B(n_11), .CI(
    in_19[9]));
  ADDFX1 cdnfadd_009_2(.CO(n_234), .S(n_233), .A(in_1[9]), .B(in_10[9]), .CI(
    n_248));
  ADDFX1 cdnfadd_009_3(.CO(n_173), .S(n_172), .A(in_13[9]), .B(in_14[9]), .CI(
    n_257));
  ADDFX1 cdnfadd_009_4(.CO(n_245), .S(n_244), .A(in_11[9]), .B(in_7[9]), .CI(
    in_4[9]));
  ADDFX1 cdnfadd_009_5(.CO(n_243), .S(n_242), .A(in_15[9]), .B(in_16[9]), .CI(
    in_2[9]));
  ADDFX1 cdnfadd_009_6(.CO(n_171), .S(n_170), .A(n_255), .B(n_253), .CI(n_246));
  ADDFX1 cdnfadd_009_7(.CO(n_121), .S(n_120), .A(n_236), .B(n_251), .CI(n_177));
  ADDFX1 cdnfadd_009_8(.CO(n_119), .S(n_118), .A(n_233), .B(n_244), .CI(n_172));
  ADDFX1 cdnfadd_009_9(.CO(n_117), .S(n_116), .A(n_175), .B(n_242), .CI(n_170));
  ADDFX1 cdnfadd_009_10(.CO(n_107), .S(n_106), .A(n_125), .B(n_159), .CI(n_120));
  ADDFX1 cdnfadd_009_11(.CO(n_105), .S(n_104), .A(n_123), .B(n_118), .CI(n_116));
  ADDFX1 cdnfadd_009_12(.CO(n_77), .S(n_76), .A(n_92), .B(n_106), .CI(n_109));
  ADDFX1 cdnfadd_009_13(.CO(n_359), .S(n_342), .A(n_104), .B(n_57), .CI(n_76));
  ADDFX1 cdnfadd_010_1(.CO(n_232), .S(n_241), .A(n_8), .B(in_12[8]), .CI(
    in_7[10]));
  ADDFX1 cdnfadd_010_2(.CO(n_229), .S(n_231), .A(n_249), .B(in_10[10]), .CI(
    in_11[10]));
  ADDFX1 cdnfadd_010_3(.CO(n_226), .S(n_240), .A(in_19[10]), .B(in_4[10]), .CI(
    in_15[10]));
  ADDFX1 cdnfadd_010_4(.CO(n_228), .S(n_239), .A(in_16[10]), .B(in_14[10]), .CI(
    in_2[10]));
  ADDFX1 cdnfadd_010_5(.CO(n_165), .S(n_164), .A(in_13[10]), .B(n_247), .CI(
    n_234));
  ADDFX1 cdnfadd_010_6(.CO(n_115), .S(n_114), .A(n_241), .B(n_173), .CI(n_243));
  ADDFX1 cdnfadd_010_7(.CO(n_157), .S(n_156), .A(n_231), .B(n_245), .CI(n_239));
  ADDFX1 cdnfadd_010_8(.CO(n_96), .S(n_95), .A(n_171), .B(n_240), .CI(n_164));
  ADDFX1 cdnfadd_010_9(.CO(n_103), .S(n_102), .A(n_121), .B(n_119), .CI(n_114));
  ADDFX1 cdnfadd_010_10(.CO(n_75), .S(n_74), .A(n_156), .B(n_95), .CI(n_117));
  ADDFX1 cdnfadd_010_11(.CO(n_73), .S(n_72), .A(n_107), .B(n_102), .CI(n_105));
  ADDFX1 cdnfadd_010_12(.CO(n_360), .S(n_343), .A(n_74), .B(n_77), .CI(n_72));
  ADDFX1 cdnfadd_011_1(.CO(n_204), .S(n_230), .A(in_14[11]), .B(in_15[11]), .CI(
    in_11[11]));
  ADDFX1 cdnfadd_011_2(.CO(n_203), .S(n_227), .A(in_10[11]), .B(n_5), .CI(
    in_19[11]));
  ADDFX1 cdnfadd_011_3(.CO(n_202), .S(n_224), .A(in_2[11]), .B(in_16[11]), .CI(
    in_13[11]));
  ADDFX1 cdnfadd_011_4(.CO(n_169), .S(n_168), .A(n_232), .B(in_4[11]), .CI(n_230));
  ADDFX1 cdnfadd_011_5(.CO(n_155), .S(n_154), .A(n_229), .B(n_228), .CI(n_227));
  ADDFX1 cdnfadd_011_6(.CO(n_94), .S(n_93), .A(n_226), .B(n_165), .CI(n_224));
  ADDFX1 cdnfadd_011_7(.CO(n_101), .S(n_100), .A(n_168), .B(n_115), .CI(n_154));
  ADDFX1 cdnfadd_011_8(.CO(n_71), .S(n_70), .A(n_157), .B(n_93), .CI(n_96));
  ADDFX1 cdnfadd_011_9(.CO(n_55), .S(n_54), .A(n_103), .B(n_100), .CI(n_75));
  ADDFX1 cdnfadd_011_10(.CO(n_361), .S(n_344), .A(n_70), .B(n_54), .CI(n_73));
  ADDFX1 cdnfadd_012_1(.CO(n_188), .S(n_205), .A(in_14[11]), .B(n_4), .CI(
    in_10[12]));
  ADDFX1 cdnfadd_012_3(.CO(n_186), .S(n_201), .A(in_16[12]), .B(in_2[12]), .CI(
    n_205));
  ADDFX1 cdnfadd_012_4(.CO(n_153), .S(n_152), .A(n_204), .B(n_203), .CI(n_24));
  ADDFX1 cdnfadd_012_5(.CO(n_151), .S(n_150), .A(n_202), .B(n_201), .CI(n_169));
  ADDFX1 cdnfadd_012_6(.CO(n_69), .S(n_68), .A(n_155), .B(n_152), .CI(n_94));
  ADDFX1 cdnfadd_012_7(.CO(n_53), .S(n_52), .A(n_150), .B(n_101), .CI(n_68));
  ADDFX1 cdnfadd_012_8(.CO(n_362), .S(n_345), .A(n_71), .B(n_52), .CI(n_55));
  ADDFX1 cdnfadd_013_0(.CO(n_178), .S(n_189), .A(n_6), .B(n_3), .CI(n_4));
  ADDFX1 cdnfadd_013_2(.CO(n_167), .S(n_166), .A(n_189), .B(n_26), .CI(n_7));
  ADDFX1 cdnfadd_013_3(.CO(n_163), .S(n_162), .A(n_12), .B(n_188), .CI(n_166));
  ADDFX1 cdnfadd_013_4(.CO(n_99), .S(n_98), .A(n_18), .B(n_186), .CI(n_162));
  ADDFX1 cdnfadd_013_5(.CO(n_67), .S(n_66), .A(n_153), .B(n_98), .CI(n_151));
  ADDFX1 cdnfadd_013_6(.CO(n_347), .S(n_346), .A(n_69), .B(n_66), .CI(n_53));
  ADDFX1 cdnfadd_014_0(.CO(n_80), .S(n_97), .A(n_29), .B(n_167), .CI(n_163));
  ADDFX1 cdnfadd_014_1(.CO(n_348), .S(n_363), .A(n_97), .B(n_99), .CI(n_67));
  OA21X1 g338(.Y(out_0[18]), .A0(n_28), .A1(n_30), .B0(n_32));
  INVX1 g339(.Y(n_32), .A(n_34));
  XOR2XL g340(.Y(n_31), .A(n_28), .B(n_30));
  INVX1 g341(.Y(n_30), .A(n_80));
  XNOR2X1 g342(.Y(n_29), .A(n_14), .B(n_178));
  NAND2BX1 g343(.Y(n_28), .AN(n_14), .B(n_178));
  AOI2BB1X1 g344(.Y(n_27), .A0N(in_5[4]), .A1N(in_3[4]), .B0(n_17));
  OAI21X1 g345(.Y(n_26), .A0(in_14[11]), .A1(n_4), .B0(n_13));
  AOI2BB1X1 g346(.Y(n_25), .A0N(in_12[0]), .A1N(n_1), .B0(n_20));
  AOI21X1 g347(.Y(n_24), .A0(n_7), .A1(n_6), .B0(n_18));
  AOI2BB1X1 g348(.Y(n_23), .A0N(in_19[2]), .A1N(in_13[2]), .B0(n_16));
  OAI2BB1X1 g349(.Y(n_22), .A0N(in_5[6]), .A1N(in_3[6]), .B0(n_15));
  AOI2BB1X1 g350(.Y(n_21), .A0N(in_5[7]), .A1N(in_3[7]), .B0(n_19));
  AND2XL g351(.Y(n_20), .A(in_12[0]), .B(n_1));
  AND2XL g352(.Y(n_19), .A(in_5[7]), .B(in_3[7]));
  NOR2X1 g353(.Y(n_18), .A(n_7), .B(n_6));
  AND2X1 g354(.Y(n_17), .A(in_5[4]), .B(in_3[4]));
  AND2XL g355(.Y(n_16), .A(in_19[2]), .B(in_13[2]));
  OR2X1 g356(.Y(n_15), .A(in_5[6]), .B(in_3[6]));
  INVX1 g357(.Y(n_14), .A(n_13));
  NAND2X1 g358(.Y(n_13), .A(in_14[11]), .B(n_4));
  INVX1 g359(.Y(n_12), .A(in_2[13]));
  INVX1 g360(.Y(n_11), .A(in_17[9]));
  INVX1 g361(.Y(n_10), .A(in_5[5]));
  INVX1 g362(.Y(n_9), .A(in_3[8]));
  INVX1 g363(.Y(n_8), .A(in_8[9]));
  INVX1 g364(.Y(n_7), .A(in_13[12]));
  INVX1 g365(.Y(n_6), .A(in_4[12]));
  INVX1 g366(.Y(n_5), .A(in_12[8]));
  INVX1 g367(.Y(n_4), .A(in_15[11]));
  INVX1 g368(.Y(n_3), .A(in_16[12]));
  INVXL drc_bufs(.Y(n_1), .A(n_0));
  INVXL drc_bufs370(.Y(n_0), .A(in_2[0]));
endmodule

module csa_tree_ADD_TC_OP_19_group_12094(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_401, n_399, n_397, n_395, n_393, n_391, n_389, n_387, n_385, n_383, 
    n_382, n_381, n_379, n_378, n_377, n_376, n_375, n_374, n_373, n_372, 
    n_371, n_370, n_369, n_367, n_366, n_365, n_364, n_363, n_362, n_361, 
    n_360, n_359, n_358, n_357, n_356, n_355, n_353, n_352, n_351, n_350, 
    n_349, n_348, n_347, n_346, n_345, n_344, n_343, n_342, n_341, n_340, 
    n_339, n_338, n_337, n_335, n_334, n_333, n_332, n_331, n_330, n_329, 
    n_328, n_327, n_326, n_325, n_324, n_323, n_322, n_321, n_320, n_319, 
    n_318, n_317, n_316, n_315, n_314, n_313, n_312, n_311, n_310, n_309, 
    n_308, n_307, n_306, n_305, n_304, n_303, n_302, n_301, n_299, n_298, 
    n_297, n_296, n_295, n_294, n_293, n_292, n_291, n_290, n_289, n_288, 
    n_287, n_286, n_285, n_284, n_283, n_282, n_281, n_280, n_279, n_278, 
    n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, n_268, 
    n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
    n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, n_249, n_248, 
    n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, 
    n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, 
    n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, n_217, 
    n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, n_207, 
    n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
    n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, n_187, 
    n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, 
    n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
    n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, 
    n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, 
    n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
    n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, 
    n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
    n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, 
    n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, 
    n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
    n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
    n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
    n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  AOI21X2 g5087(.Y(out_0[18]), .A0(n_9), .A1(n_193), .B0(n_401));
  ADDFX1 g5088(.CO(n_401), .S(out_0[15]), .A(n_198), .B(n_281), .CI(n_399));
  ADDFX1 g5089(.CO(n_399), .S(out_0[14]), .A(n_282), .B(n_357), .CI(n_397));
  ADDFX1 g5090(.CO(n_397), .S(out_0[13]), .A(n_358), .B(n_369), .CI(n_395));
  ADDFX1 g5091(.CO(n_395), .S(out_0[12]), .A(n_370), .B(n_381), .CI(n_393));
  ADDFX1 g5092(.CO(n_393), .S(out_0[11]), .A(n_377), .B(n_382), .CI(n_391));
  ADDFX1 g5093(.CO(n_391), .S(out_0[10]), .A(n_375), .B(n_378), .CI(n_389));
  ADDFX1 g5094(.CO(n_389), .S(out_0[9]), .A(n_373), .B(n_376), .CI(n_387));
  ADDFX1 g5095(.CO(n_387), .S(out_0[8]), .A(n_371), .B(n_374), .CI(n_385));
  ADDFX1 g5096(.CO(n_385), .S(out_0[7]), .A(n_372), .B(n_363), .CI(n_383));
  ADDFX1 g5097(.CO(n_383), .S(out_0[6]), .A(n_355), .B(n_379), .CI(n_364));
  ADDFX1 g5098(.CO(n_381), .S(n_382), .A(n_345), .B(n_365), .CI(n_360));
  ADDFX1 g5099(.CO(n_379), .S(out_0[5]), .A(n_337), .B(n_367), .CI(n_356));
  ADDFX1 g5100(.CO(n_377), .S(n_378), .A(n_346), .B(n_361), .CI(n_366));
  ADDFX1 g5101(.CO(n_375), .S(n_376), .A(n_349), .B(n_340), .CI(n_362));
  ADDFX1 g5102(.CO(n_373), .S(n_374), .A(n_334), .B(n_351), .CI(n_350));
  ADDFX1 g5103(.CO(n_371), .S(n_372), .A(n_328), .B(n_341), .CI(n_352));
  ADDFX1 g5104(.CO(n_369), .S(n_370), .A(n_343), .B(n_348), .CI(n_359));
  ADDFX1 g5105(.CO(n_367), .S(out_0[4]), .A(n_322), .B(n_338), .CI(n_353));
  ADDFX1 g5106(.CO(n_365), .S(n_366), .A(n_331), .B(n_312), .CI(n_339));
  ADDFX1 g5107(.CO(n_363), .S(n_364), .A(n_329), .B(n_326), .CI(n_342));
  ADDFX1 g5108(.CO(n_361), .S(n_362), .A(n_313), .B(n_332), .CI(n_333));
  ADDFX1 g5109(.CO(n_359), .S(n_360), .A(n_311), .B(n_316), .CI(n_344));
  ADDFX1 g5110(.CO(n_357), .S(n_358), .A(n_289), .B(n_258), .CI(n_347));
  ADDFX1 g5111(.CO(n_355), .S(n_356), .A(n_321), .B(n_318), .CI(n_330));
  ADDFX1 g5112(.CO(n_353), .S(out_0[3]), .A(n_302), .B(n_335), .CI(n_320));
  ADDFX1 g5113(.CO(n_351), .S(n_352), .A(n_291), .B(n_325), .CI(n_308));
  ADDFX1 g5114(.CO(n_349), .S(n_350), .A(n_307), .B(n_314), .CI(n_327));
  ADDFX1 g5115(.CO(n_347), .S(n_348), .A(n_221), .B(n_315), .CI(n_290));
  ADDFX1 g5116(.CO(n_345), .S(n_346), .A(n_309), .B(n_246), .CI(n_324));
  ADDFX1 g5117(.CO(n_343), .S(n_344), .A(n_230), .B(n_323), .CI(n_222));
  ADDFX1 g5118(.CO(n_341), .S(n_342), .A(n_287), .B(n_317), .CI(n_292));
  ADDFX1 g5119(.CO(n_339), .S(n_340), .A(n_267), .B(n_272), .CI(n_310));
  ADDFX1 g5120(.CO(n_337), .S(n_338), .A(n_301), .B(n_304), .CI(n_319));
  ADDFX1 g5121(.CO(n_335), .S(out_0[2]), .A(n_299), .B(n_250), .CI(n_306));
  ADDFX1 g5122(.CO(n_333), .S(n_334), .A(n_296), .B(n_294), .CI(n_268));
  ADDFX1 g5123(.CO(n_331), .S(n_332), .A(n_274), .B(n_284), .CI(n_295));
  ADDFX1 g5124(.CO(n_329), .S(n_330), .A(n_278), .B(n_303), .CI(n_288));
  ADDFX1 g5125(.CO(n_327), .S(n_328), .A(n_279), .B(n_260), .CI(n_298));
  ADDFX1 g5126(.CO(n_325), .S(n_326), .A(n_277), .B(n_280), .CI(n_266));
  ADDFX1 g5127(.CO(n_323), .S(n_324), .A(n_283), .B(n_39), .CI(n_188));
  ADDFX1 g5128(.CO(n_321), .S(n_322), .A(n_275), .B(n_270), .CI(n_286));
  ADDFX1 g5129(.CO(n_319), .S(n_320), .A(n_254), .B(n_305), .CI(n_276));
  ADDFX1 g5130(.CO(n_317), .S(n_318), .A(n_269), .B(n_256), .CI(n_285));
  ADDFX1 g5131(.CO(n_315), .S(n_316), .A(n_263), .B(n_159), .CI(n_245));
  ADDFX1 g5132(.CO(n_313), .S(n_314), .A(n_261), .B(n_259), .CI(n_297));
  ADDFX1 g5133(.CO(n_311), .S(n_312), .A(n_273), .B(n_264), .CI(n_271));
  ADDFX1 g5134(.CO(n_309), .S(n_310), .A(n_201), .B(n_169), .CI(n_293));
  ADDFX1 g5135(.CO(n_307), .S(n_308), .A(n_226), .B(n_265), .CI(n_262));
  ADDFX1 g5136(.CO(n_305), .S(n_306), .A(n_247), .B(n_252), .CI(n_206));
  ADDFX1 g5137(.CO(n_303), .S(n_304), .A(n_215), .B(n_253), .CI(n_244));
  ADDFX1 g5138(.CO(n_301), .S(n_302), .A(n_228), .B(n_249), .CI(n_216));
  ADDFX1 g5139(.CO(n_299), .S(out_0[1]), .A(n_217), .B(n_180), .CI(n_248));
  ADDFX1 g5140(.CO(n_297), .S(n_298), .A(n_177), .B(n_242), .CI(n_237));
  ADDFX1 g5141(.CO(n_295), .S(n_296), .A(n_225), .B(n_103), .CI(n_241));
  ADDFX1 g5142(.CO(n_293), .S(n_294), .A(n_194), .B(n_123), .CI(n_240));
  ADDFX1 g5143(.CO(n_291), .S(n_292), .A(n_255), .B(n_220), .CI(n_238));
  ADDFX1 g5144(.CO(n_289), .S(n_290), .A(n_229), .B(n_143), .CI(n_208));
  ADDFX1 g5145(.CO(n_287), .S(n_288), .A(n_243), .B(n_234), .CI(n_236));
  ADDFX1 g5146(.CO(n_285), .S(n_286), .A(n_227), .B(n_165), .CI(n_232));
  ADDFX1 g5147(.CO(n_283), .S(n_284), .A(n_87), .B(n_37), .CI(n_239));
  ADDFX1 g5148(.CO(n_281), .S(n_282), .A(n_174), .B(n_196), .CI(n_257));
  ADDFX1 g5149(.CO(n_279), .S(n_280), .A(n_204), .B(n_233), .CI(n_178));
  ADDFX1 g5150(.CO(n_277), .S(n_278), .A(n_171), .B(n_192), .CI(n_231));
  ADDFX1 g5151(.CO(n_275), .S(n_276), .A(n_251), .B(n_210), .CI(n_205));
  ADDFX1 g5152(.CO(n_273), .S(n_274), .A(n_212), .B(n_102), .CI(n_213));
  ADDFX1 g5153(.CO(n_271), .S(n_272), .A(n_223), .B(n_111), .CI(n_45));
  ADDFX1 g5154(.CO(n_269), .S(n_270), .A(n_209), .B(n_151), .CI(n_200));
  ADDFX1 g5155(.CO(n_267), .S(n_268), .A(n_214), .B(n_202), .CI(n_224));
  ADDFX1 g5156(.CO(n_265), .S(n_266), .A(n_191), .B(n_75), .CI(n_235));
  ADDFX1 g5157(.CO(n_263), .S(n_264), .A(n_211), .B(n_73), .CI(n_44));
  ADDFX1 g5158(.CO(n_261), .S(n_262), .A(n_203), .B(n_125), .CI(n_157));
  ADDFX1 g5159(.CO(n_259), .S(n_260), .A(n_219), .B(n_195), .CI(n_79));
  ADDFX1 g5160(.CO(n_257), .S(n_258), .A(n_142), .B(n_197), .CI(n_207));
  ADDFX1 g5161(.CO(n_255), .S(n_256), .A(n_199), .B(n_164), .CI(n_107));
  ADDFX1 g5162(.CO(n_253), .S(n_254), .A(n_185), .B(n_147), .CI(n_183));
  ADDFX1 g5163(.CO(n_251), .S(n_252), .A(n_181), .B(n_173), .CI(n_160));
  ADDFX1 g5164(.CO(n_249), .S(n_250), .A(n_184), .B(n_179), .CI(n_186));
  ADDFX1 g5165(.CO(n_247), .S(n_248), .A(n_144), .B(n_182), .CI(n_161));
  ADDFX1 g5166(.CO(n_245), .S(n_246), .A(n_28), .B(n_168), .CI(n_167));
  ADDFX1 g5167(.CO(n_243), .S(n_244), .A(n_146), .B(n_97), .CI(n_153));
  ADDFX1 g5168(.CO(n_241), .S(n_242), .A(n_74), .B(n_189), .CI(n_131));
  ADDFX1 g5169(.CO(n_239), .S(n_240), .A(n_175), .B(in_14[8]), .CI(in_6[8]));
  ADDFX1 g5170(.CO(n_237), .S(n_238), .A(n_170), .B(n_190), .CI(n_33));
  ADDFX1 g5171(.CO(n_235), .S(n_236), .A(n_96), .B(n_152), .CI(n_137));
  ADDFX1 g5172(.CO(n_233), .S(n_234), .A(n_163), .B(n_150), .CI(n_95));
  ADDFX1 g5173(.CO(n_231), .S(n_232), .A(n_154), .B(n_133), .CI(n_77));
  ADDFX1 g5174(.CO(n_229), .S(n_230), .A(n_22), .B(n_27), .CI(n_166));
  ADDFX1 g5175(.CO(n_227), .S(n_228), .A(n_172), .B(n_67), .CI(n_83));
  ADDFX1 g5176(.CO(n_225), .S(n_226), .A(n_176), .B(n_148), .CI(n_32));
  ADDFX1 g5177(.CO(n_223), .S(n_224), .A(n_156), .B(n_78), .CI(n_91));
  ADDFX1 g5178(.CO(n_221), .S(n_222), .A(n_38), .B(n_187), .CI(n_121));
  ADDFX1 g5179(.CO(n_219), .S(n_220), .A(n_149), .B(n_136), .CI(n_106));
  ADDFX1 g5180(.CO(n_217), .S(out_0[0]), .A(n_81), .B(n_41), .CI(n_145));
  ADDFX1 g5181(.CO(n_215), .S(n_216), .A(n_155), .B(n_127), .CI(n_93));
  ADDFX1 g5182(.CO(n_213), .S(n_214), .A(n_141), .B(n_18), .CI(in_17[8]));
  ADDFX1 g5183(.CO(n_211), .S(n_212), .A(n_140), .B(n_7), .CI(in_11[9]));
  ADDFX1 g5184(.CO(n_209), .S(n_210), .A(n_85), .B(n_138), .CI(n_30));
  ADDFX1 g5185(.CO(n_207), .S(n_208), .A(n_113), .B(n_120), .CI(n_158));
  ADDFX1 g5186(.CO(n_205), .S(n_206), .A(n_139), .B(n_99), .CI(n_31));
  ADDFX1 g5187(.CO(n_203), .S(n_204), .A(n_57), .B(n_58), .CI(n_162));
  ADDFX1 g5188(.CO(n_201), .S(n_202), .A(n_128), .B(n_124), .CI(n_130));
  ADDFX1 g5189(.CO(n_199), .S(n_200), .A(n_84), .B(n_66), .CI(n_126));
  MXI2XL g5190(.Y(n_198), .A(n_29), .B(n_9), .S0(n_193));
  ADDFX1 g5191(.CO(n_196), .S(n_197), .A(n_48), .B(n_112), .CI(n_135));
  ADDFX1 g5192(.CO(n_194), .S(n_195), .A(n_88), .B(n_129), .CI(in_17[7]));
  ADDFX1 g5193(.CO(n_191), .S(n_192), .A(n_100), .B(n_76), .CI(n_47));
  ADDFX1 g5194(.CO(n_189), .S(n_190), .A(n_109), .B(in_7[6]), .CI(in_17[6]));
  ADDFX1 g5195(.CO(n_187), .S(n_188), .A(n_36), .B(in_7[10]), .CI(n_110));
  ADDFX1 g5196(.CO(n_185), .S(n_186), .A(n_51), .B(n_34), .CI(n_116));
  ADDFX1 g5197(.CO(n_183), .S(n_184), .A(n_71), .B(n_114), .CI(n_61));
  ADDFX1 g5198(.CO(n_181), .S(n_182), .A(n_62), .B(n_80), .CI(n_40));
  ADDFX1 g5199(.CO(n_179), .S(n_180), .A(n_105), .B(n_115), .CI(n_117));
  ADDFX1 g5200(.CO(n_177), .S(n_178), .A(n_94), .B(n_46), .CI(n_89));
  ADDFX1 g5201(.CO(n_175), .S(n_176), .A(in_16[6]), .B(n_108), .CI(in_2[7]));
  ADDFX1 g5202(.CO(n_193), .S(n_174), .A(n_13), .B(n_29), .CI(n_134));
  ADDFX1 g5203(.CO(n_172), .S(n_173), .A(n_104), .B(n_64), .CI(n_118));
  ADDFX1 g5204(.CO(n_170), .S(n_171), .A(n_59), .B(in_14[5]), .CI(n_132));
  ADDFX1 g5205(.CO(n_168), .S(n_169), .A(n_90), .B(in_14[9]), .CI(n_122));
  ADDFX1 g5206(.CO(n_166), .S(n_167), .A(n_86), .B(in_9[10]), .CI(in_14[10]));
  ADDFX1 g5207(.CO(n_164), .S(n_165), .A(n_82), .B(n_92), .CI(n_101));
  ADDFX1 g5208(.CO(n_162), .S(n_163), .A(n_10), .B(n_54), .CI(in_3[5]));
  ADDFX1 g5209(.CO(n_160), .S(n_161), .A(n_119), .B(n_65), .CI(n_35));
  ADDFX1 g5210(.CO(n_158), .S(n_159), .A(n_72), .B(in_17[11]), .CI(in_14[11]));
  ADDFX1 g5211(.CO(n_156), .S(n_157), .A(n_56), .B(in_7[7]), .CI(in_4[7]));
  ADDFX1 g5212(.CO(n_154), .S(n_155), .A(n_25), .B(n_50), .CI(n_70));
  ADDFX1 g5213(.CO(n_152), .S(n_153), .A(n_68), .B(in_4[4]), .CI(in_14[4]));
  ADDFX1 g5214(.CO(n_150), .S(n_151), .A(n_16), .B(n_55), .CI(in_9[4]));
  ADDFX1 g5215(.CO(n_148), .S(n_149), .A(n_42), .B(in_8[6]), .CI(in_12[6]));
  ADDFX1 g5216(.CO(n_146), .S(n_147), .A(n_69), .B(n_60), .CI(n_98));
  ADDFX1 g5217(.CO(n_144), .S(n_145), .A(in_16[0]), .B(n_24), .CI(n_63));
  ADDFX1 g5218(.CO(n_142), .S(n_143), .A(n_21), .B(n_49), .CI(in_17[12]));
  ADDFX1 g5219(.CO(n_140), .S(n_141), .A(in_18[8]), .B(n_12), .CI(n_52));
  ADDFX1 g5220(.CO(n_138), .S(n_139), .A(n_26), .B(in_8[2]), .CI(in_6[2]));
  ADDFX1 g5221(.CO(n_136), .S(n_137), .A(n_43), .B(in_17[5]), .CI(in_11[5]));
  ADDFX1 g5222(.CO(n_134), .S(n_135), .A(n_0), .B(n_1), .CI(n_5));
  ADDFX1 g5223(.CO(n_132), .S(n_133), .A(n_19), .B(in_8[4]), .CI(in_6[4]));
  ADDFX1 g5224(.CO(n_130), .S(n_131), .A(n_15), .B(in_19[7]), .CI(in_3[7]));
  ADDFX1 g5225(.CO(n_128), .S(n_129), .A(n_53), .B(in_5[7]), .CI(in_10[7]));
  ADDFX1 g5226(.CO(n_126), .S(n_127), .A(n_20), .B(in_6[3]), .CI(in_9[3]));
  ADDFX1 g5227(.CO(n_124), .S(n_125), .A(in_8[7]), .B(in_11[7]), .CI(in_12[7]));
  ADDFX1 g5228(.CO(n_122), .S(n_123), .A(in_12[8]), .B(in_19[8]), .CI(in_11[8]));
  ADDFX1 g5229(.CO(n_120), .S(n_121), .A(n_14), .B(in_4[11]), .CI(in_9[11]));
  ADDFX1 g5230(.CO(n_118), .S(n_119), .A(in_0[1]), .B(in_1[1]), .CI(n_2));
  ADDFX1 g5231(.CO(n_116), .S(n_117), .A(in_12[1]), .B(in_3[1]), .CI(in_4[1]));
  ADDFX1 g5232(.CO(n_114), .S(n_115), .A(n_23), .B(in_6[1]), .CI(in_11[1]));
  ADDFX1 g5233(.CO(n_112), .S(n_113), .A(n_11), .B(in_14[12]), .CI(in_9[12]));
  ADDFX1 g5234(.CO(n_110), .S(n_111), .A(n_17), .B(in_8[9]), .CI(in_4[9]));
  ADDFX1 g5235(.CO(n_108), .S(n_109), .A(in_1[6]), .B(in_15[6]), .CI(in_18[6]));
  ADDFX1 g5236(.CO(n_106), .S(n_107), .A(in_7[5]), .B(in_4[5]), .CI(in_9[5]));
  ADDFX1 g5237(.CO(n_104), .S(n_105), .A(in_7[1]), .B(in_16[1]), .CI(in_15[1]));
  ADDFX1 g5238(.CO(n_102), .S(n_103), .A(in_8[8]), .B(in_4[8]), .CI(in_9[8]));
  ADDFX1 g5239(.CO(n_100), .S(n_101), .A(in_10[4]), .B(in_19[4]), .CI(in_2[4]));
  ADDFX1 g5240(.CO(n_98), .S(n_99), .A(in_2[2]), .B(in_9[2]), .CI(in_3[2]));
  ADDFX1 g5241(.CO(n_96), .S(n_97), .A(in_11[4]), .B(in_7[4]), .CI(in_17[4]));
  ADDFX1 g5242(.CO(n_94), .S(n_95), .A(in_8[5]), .B(in_2[5]), .CI(in_12[5]));
  ADDFX1 g5243(.CO(n_92), .S(n_93), .A(in_17[3]), .B(in_8[3]), .CI(in_3[3]));
  ADDFX1 g5244(.CO(n_90), .S(n_91), .A(in_2[8]), .B(in_3[8]), .CI(in_7[8]));
  ADDFX1 g5245(.CO(n_88), .S(n_89), .A(in_5[6]), .B(in_19[6]), .CI(in_2[6]));
  ADDFX1 g5246(.CO(n_86), .S(n_87), .A(in_5[9]), .B(in_2[9]), .CI(in_10[9]));
  ADDFX1 g5247(.CO(n_84), .S(n_85), .A(in_7[3]), .B(in_5[3]), .CI(in_14[3]));
  ADDFX1 g5248(.CO(n_82), .S(n_83), .A(in_12[3]), .B(in_11[3]), .CI(in_4[3]));
  ADDFX1 g5249(.CO(n_80), .S(n_81), .A(in_3[0]), .B(in_7[0]), .CI(in_9[0]));
  ADDFX1 g5250(.CO(n_78), .S(n_79), .A(in_6[7]), .B(in_9[7]), .CI(in_14[7]));
  ADDFX1 g5251(.CO(n_76), .S(n_77), .A(in_5[4]), .B(in_12[4]), .CI(in_3[4]));
  ADDFX1 g5252(.CO(n_74), .S(n_75), .A(in_4[6]), .B(in_6[6]), .CI(in_9[6]));
  ADDFX1 g5253(.CO(n_72), .S(n_73), .A(in_5[10]), .B(in_8[10]), .CI(in_11[10]));
  ADDFX1 g5254(.CO(n_70), .S(n_71), .A(in_15[2]), .B(in_7[2]), .CI(in_18[2]));
  ADDFX1 g5255(.CO(n_68), .S(n_69), .A(in_1[3]), .B(in_15[3]), .CI(in_18[3]));
  ADDFX1 g5256(.CO(n_66), .S(n_67), .A(in_19[3]), .B(in_10[3]), .CI(in_2[3]));
  ADDFX1 g5257(.CO(n_64), .S(n_65), .A(in_14[1]), .B(in_19[1]), .CI(in_17[1]));
  ADDFX1 g5258(.CO(n_62), .S(n_63), .A(in_4[0]), .B(in_6[0]), .CI(in_11[0]));
  ADDFX1 g5259(.CO(n_60), .S(n_61), .A(in_16[2]), .B(in_14[2]), .CI(in_17[2]));
  ADDFX1 g5260(.CO(n_58), .S(n_59), .A(in_15[5]), .B(in_18[5]), .CI(in_5[5]));
  ADDFX1 g5261(.CO(n_56), .S(n_57), .A(in_0[6]), .B(n_4), .CI(in_10[6]));
  ADDFX1 g5262(.CO(n_54), .S(n_55), .A(in_0[4]), .B(in_1[4]), .CI(in_18[4]));
  ADDFX1 g5263(.CO(n_52), .S(n_53), .A(in_0[7]), .B(in_1[7]), .CI(in_18[7]));
  ADDFX1 g5264(.CO(n_50), .S(n_51), .A(in_5[2]), .B(in_1[2]), .CI(in_10[2]));
  ADDFX1 g5265(.CO(n_48), .S(n_49), .A(n_6), .B(in_7[11]), .CI(in_4[12]));
  ADDFX1 g5266(.CO(n_46), .S(n_47), .A(in_10[5]), .B(in_19[5]), .CI(in_6[5]));
  ADDFX1 g5267(.CO(n_44), .S(n_45), .A(in_7[9]), .B(in_9[9]), .CI(in_17[9]));
  ADDFX1 g5268(.CO(n_42), .S(n_43), .A(in_0[5]), .B(in_1[5]), .CI(in_16[5]));
  ADDFX1 g5269(.CO(n_40), .S(n_41), .A(in_1[0]), .B(in_12[0]), .CI(in_0[0]));
  ADDFX1 g5270(.CO(n_38), .S(n_39), .A(n_8), .B(in_4[10]), .CI(in_17[10]));
  ADDFX1 g5271(.CO(n_36), .S(n_37), .A(in_12[9]), .B(in_6[9]), .CI(in_19[9]));
  ADDFX1 g5272(.CO(n_34), .S(n_35), .A(in_8[1]), .B(in_18[1]), .CI(in_9[1]));
  ADDFX1 g5273(.CO(n_32), .S(n_33), .A(in_11[6]), .B(in_3[6]), .CI(in_14[6]));
  ADDFX1 g5274(.CO(n_30), .S(n_31), .A(in_12[2]), .B(in_11[2]), .CI(in_4[2]));
  INVX1 g5275(.Y(n_29), .A(n_9));
  ADDHX1 g5276(.CO(n_27), .S(n_28), .A(in_10[10]), .B(in_19[10]));
  ADDHX1 g5277(.CO(n_25), .S(n_26), .A(in_0[2]), .B(in_19[2]));
  ADDHX1 g5278(.CO(n_23), .S(n_24), .A(in_15[0]), .B(in_19[0]));
  ADDHX1 g5279(.CO(n_21), .S(n_22), .A(in_7[11]), .B(in_19[11]));
  ADDHX1 g5280(.CO(n_19), .S(n_20), .A(in_16[3]), .B(in_0[3]));
  ADDHX1 g5281(.CO(n_17), .S(n_18), .A(in_5[8]), .B(in_10[8]));
  OAI2BB1X1 g5282(.Y(n_16), .A0N(in_16[4]), .A1N(in_15[4]), .B0(n_10));
  OAI2BB1X1 g5283(.Y(n_15), .A0N(in_16[7]), .A1N(in_15[7]), .B0(n_12));
  MX2XL g5284(.Y(n_14), .A(n_6), .B(in_5[10]), .S0(in_10[11]));
  NOR2X1 g5287(.Y(n_13), .A(in_4[12]), .B(in_9[12]));
  OR2X1 g5288(.Y(n_12), .A(in_16[7]), .B(in_15[7]));
  NOR2X1 g5289(.Y(n_11), .A(n_6), .B(in_10[11]));
  OR2X1 g5290(.Y(n_10), .A(in_16[4]), .B(in_15[4]));
  NOR2X1 g5291(.Y(n_9), .A(in_7[11]), .B(in_14[12]));
  INVX1 g5292(.Y(n_8), .A(in_2[10]));
  INVX1 g5294(.Y(n_7), .A(in_3[8]));
  INVX1 g5296(.Y(n_6), .A(in_5[10]));
  INVX1 g5297(.Y(n_5), .A(in_17[13]));
  INVX1 g5299(.Y(n_4), .A(in_16[6]));
  BUFX2 drc_bufs(.Y(n_2), .A(in_2[1]));
  CLKXOR2X1 g2(.Y(n_1), .A(in_4[12]), .B(in_9[12]));
  CLKXOR2X1 g5303(.Y(n_0), .A(in_7[11]), .B(in_14[12]));
endmodule

module csa_tree_ADD_TC_OP_19_group_10152(in_0, in_1, in_2, in_3, in_4, in_5, 
    in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, 
    in_17, in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_375, n_373, n_371, n_369, n_367, n_365, n_363, n_361, n_359, n_357, 
    n_356, n_355, n_354, n_353, n_351, n_350, n_349, n_348, n_347, n_346, 
    n_345, n_344, n_343, n_342, n_341, n_340, n_339, n_338, n_337, n_336, 
    n_335, n_334, n_333, n_332, n_331, n_330, n_329, n_328, n_327, n_326, 
    n_325, n_324, n_323, n_322, n_321, n_320, n_319, n_317, n_316, n_315, 
    n_314, n_313, n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, 
    n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, 
    n_294, n_293, n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, 
    n_284, n_283, n_282, n_280, n_279, n_278, n_277, n_276, n_275, n_274, 
    n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, 
    n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
    n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_236, n_235, n_234, n_233, 
    n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
    n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, 
    n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, 
    n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, 
    n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
    n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, 
    n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
    n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_152, 
    n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, 
    n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, 
    n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, 
    n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
    n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, 
    n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, 
    n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
    n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  AOI21X2 g4698(.Y(out_0[18]), .A0(n_108), .A1(n_277), .B0(n_375));
  ADDFX1 g4699(.CO(n_375), .S(out_0[14]), .A(n_296), .B(n_325), .CI(n_373));
  ADDFX1 g4700(.CO(n_373), .S(out_0[13]), .A(n_326), .B(n_343), .CI(n_371));
  ADDFX1 g4701(.CO(n_371), .S(out_0[12]), .A(n_344), .B(n_355), .CI(n_369));
  ADDFX1 g4702(.CO(n_369), .S(out_0[11]), .A(n_347), .B(n_356), .CI(n_367));
  ADDFX1 g4703(.CO(n_367), .S(out_0[10]), .A(n_349), .B(n_365), .CI(n_348));
  ADDFX1 g4704(.CO(n_365), .S(out_0[9]), .A(n_353), .B(n_350), .CI(n_363));
  ADDFX1 g4705(.CO(n_363), .S(out_0[8]), .A(n_345), .B(n_354), .CI(n_361));
  ADDFX1 g4706(.CO(n_361), .S(out_0[7]), .A(n_341), .B(n_346), .CI(n_359));
  ADDFX1 g4707(.CO(n_359), .S(out_0[6]), .A(n_339), .B(n_342), .CI(n_357));
  ADDFX1 g4708(.CO(n_357), .S(out_0[5]), .A(n_327), .B(n_340), .CI(n_351));
  ADDFX1 g4709(.CO(n_355), .S(n_356), .A(n_312), .B(n_333), .CI(n_332));
  ADDFX1 g4710(.CO(n_353), .S(n_354), .A(n_335), .B(n_320), .CI(n_330));
  ADDFX1 g4711(.CO(n_351), .S(out_0[4]), .A(n_284), .B(n_317), .CI(n_328));
  ADDFX1 g4712(.CO(n_349), .S(n_350), .A(n_329), .B(n_310), .CI(n_338));
  ADDFX1 g4713(.CO(n_347), .S(n_348), .A(n_316), .B(n_337), .CI(n_334));
  ADDFX1 g4714(.CO(n_345), .S(n_346), .A(n_323), .B(n_308), .CI(n_336));
  ADDFX1 g4715(.CO(n_343), .S(n_344), .A(n_311), .B(n_306), .CI(n_331));
  ADDFX1 g4716(.CO(n_341), .S(n_342), .A(n_321), .B(n_314), .CI(n_324));
  ADDFX1 g4717(.CO(n_339), .S(n_340), .A(n_290), .B(n_295), .CI(n_322));
  ADDFX1 g4718(.CO(n_337), .S(n_338), .A(n_301), .B(n_304), .CI(n_319));
  ADDFX1 g4719(.CO(n_335), .S(n_336), .A(n_286), .B(n_313), .CI(n_289));
  ADDFX1 g4720(.CO(n_333), .S(n_334), .A(n_303), .B(n_309), .CI(n_300));
  ADDFX1 g4721(.CO(n_331), .S(n_332), .A(n_299), .B(n_271), .CI(n_315));
  ADDFX1 g4722(.CO(n_329), .S(n_330), .A(n_273), .B(n_302), .CI(n_307));
  ADDFX1 g4723(.CO(n_327), .S(n_328), .A(n_258), .B(n_293), .CI(n_291));
  ADDFX1 g4724(.CO(n_325), .S(n_326), .A(n_276), .B(n_278), .CI(n_305));
  ADDFX1 g4725(.CO(n_323), .S(n_324), .A(n_261), .B(n_294), .CI(n_287));
  ADDFX1 g4726(.CO(n_321), .S(n_322), .A(n_292), .B(n_249), .CI(n_298));
  ADDFX1 g4727(.CO(n_319), .S(n_320), .A(n_282), .B(n_288), .CI(n_267));
  ADDFX1 g4728(.CO(n_317), .S(out_0[3]), .A(n_280), .B(n_259), .CI(n_285));
  ADDFX1 g4729(.CO(n_315), .S(n_316), .A(n_263), .B(n_268), .CI(n_275));
  ADDFX1 g4730(.CO(n_313), .S(n_314), .A(n_221), .B(n_297), .CI(n_235));
  ADDFX1 g4731(.CO(n_311), .S(n_312), .A(n_262), .B(n_265), .CI(n_274));
  ADDFX1 g4732(.CO(n_309), .S(n_310), .A(n_272), .B(n_255), .CI(n_269));
  ADDFX1 g4733(.CO(n_307), .S(n_308), .A(n_260), .B(n_283), .CI(n_209));
  ADDFX1 g4734(.CO(n_305), .S(n_306), .A(n_264), .B(n_279), .CI(n_270));
  ADDFX1 g4735(.CO(n_303), .S(n_304), .A(n_201), .B(n_247), .CI(n_266));
  ADDFX1 g4736(.CO(n_301), .S(n_302), .A(n_250), .B(n_205), .CI(n_233));
  ADDFX1 g4737(.CO(n_299), .S(n_300), .A(n_246), .B(n_254), .CI(n_217));
  ADDFX1 g4738(.CO(n_297), .S(n_298), .A(n_244), .B(n_191), .CI(n_189));
  XOR2XL g4739(.Y(n_296), .A(n_108), .B(n_277));
  ADDFX1 g4740(.CO(n_294), .S(n_295), .A(n_212), .B(n_252), .CI(n_231));
  ADDFX1 g4741(.CO(n_292), .S(n_293), .A(n_242), .B(n_163), .CI(n_245));
  ADDFX1 g4742(.CO(n_290), .S(n_291), .A(n_240), .B(n_253), .CI(n_213));
  ADDFX1 g4743(.CO(n_288), .S(n_289), .A(n_234), .B(n_251), .CI(n_218));
  ADDFX1 g4744(.CO(n_286), .S(n_287), .A(n_230), .B(n_248), .CI(n_219));
  ADDFX1 g4745(.CO(n_284), .S(n_285), .A(n_243), .B(n_238), .CI(n_241));
  ADDFX1 g4746(.CO(n_282), .S(n_283), .A(n_220), .B(n_211), .CI(n_215));
  ADDFX1 g4747(.CO(n_280), .S(out_0[2]), .A(n_236), .B(n_227), .CI(n_239));
  ADDFX1 g4748(.CO(n_278), .S(n_279), .A(n_207), .B(n_222), .CI(n_257));
  ADDFX1 g4749(.CO(n_277), .S(n_276), .A(n_206), .B(n_109), .CI(n_256));
  ADDFX1 g4750(.CO(n_274), .S(n_275), .A(n_199), .B(n_200), .CI(n_225));
  ADDFX1 g4751(.CO(n_272), .S(n_273), .A(n_210), .B(n_193), .CI(n_208));
  ADDFX1 g4752(.CO(n_270), .S(n_271), .A(n_216), .B(n_229), .CI(n_223));
  ADDFX1 g4753(.CO(n_268), .S(n_269), .A(n_204), .B(n_197), .CI(n_232));
  ADDFX1 g4754(.CO(n_266), .S(n_267), .A(n_214), .B(n_195), .CI(n_131));
  ADDFX1 g4755(.CO(n_264), .S(n_265), .A(n_198), .B(n_70), .CI(n_224));
  ADDFX1 g4756(.CO(n_262), .S(n_263), .A(n_202), .B(n_71), .CI(n_196));
  ADDFX1 g4757(.CO(n_260), .S(n_261), .A(n_177), .B(n_190), .CI(n_188));
  ADDFX1 g4758(.CO(n_258), .S(n_259), .A(n_184), .B(n_226), .CI(n_183));
  ADDFX1 g4759(.CO(n_256), .S(n_257), .A(n_154), .B(in_2[12]), .CI(n_228));
  ADDFX1 g4760(.CO(n_254), .S(n_255), .A(n_192), .B(n_203), .CI(n_165));
  ADDFX1 g4761(.CO(n_252), .S(n_253), .A(n_186), .B(n_167), .CI(n_182));
  ADDFX1 g4762(.CO(n_250), .S(n_251), .A(n_176), .B(n_143), .CI(n_174));
  ADDFX1 g4763(.CO(n_248), .S(n_249), .A(n_157), .B(n_162), .CI(n_169));
  ADDFX1 g4764(.CO(n_246), .S(n_247), .A(n_57), .B(n_172), .CI(n_194));
  ADDFX1 g4765(.CO(n_244), .S(n_245), .A(n_160), .B(n_119), .CI(n_148));
  ADDFX1 g4766(.CO(n_242), .S(n_243), .A(n_161), .B(n_180), .CI(n_105));
  ADDFX1 g4767(.CO(n_240), .S(n_241), .A(n_178), .B(n_187), .CI(n_149));
  ADDFX1 g4768(.CO(n_238), .S(n_239), .A(n_179), .B(n_170), .CI(n_185));
  ADDFX1 g4769(.CO(n_236), .S(out_0[1]), .A(n_152), .B(n_129), .CI(n_171));
  ADDFX1 g4770(.CO(n_234), .S(n_235), .A(n_168), .B(n_175), .CI(n_85));
  ADDFX1 g4771(.CO(n_232), .S(n_233), .A(n_159), .B(n_110), .CI(n_173));
  ADDFX1 g4772(.CO(n_230), .S(n_231), .A(n_138), .B(n_166), .CI(n_151));
  ADDFX1 g4773(.CO(n_228), .S(n_229), .A(n_136), .B(n_16), .CI(n_135));
  ADDFX1 g4774(.CO(n_226), .S(n_227), .A(n_128), .B(n_103), .CI(n_181));
  ADDFX1 g4775(.CO(n_224), .S(n_225), .A(n_24), .B(n_137), .CI(in_2[10]));
  ADDFX1 g4776(.CO(n_222), .S(n_223), .A(n_155), .B(n_144), .CI(in_2[11]));
  ADDFX1 g4777(.CO(n_220), .S(n_221), .A(n_61), .B(n_150), .CI(n_120));
  ADDFX1 g4778(.CO(n_218), .S(n_219), .A(n_133), .B(n_156), .CI(n_49));
  ADDFX1 g4779(.CO(n_216), .S(n_217), .A(n_56), .B(n_164), .CI(n_145));
  ADDFX1 g4780(.CO(n_214), .S(n_215), .A(n_147), .B(n_107), .CI(n_84));
  ADDFX1 g4781(.CO(n_212), .S(n_213), .A(n_47), .B(n_117), .CI(n_139));
  ADDFX1 g4782(.CO(n_210), .S(n_211), .A(n_132), .B(n_60), .CI(n_48));
  ADDFX1 g4783(.CO(n_208), .S(n_209), .A(n_141), .B(n_113), .CI(n_111));
  ADDFX1 g4784(.CO(n_206), .S(n_207), .A(n_6), .B(n_27), .CI(n_134));
  ADDFX1 g4785(.CO(n_204), .S(n_205), .A(n_112), .B(n_83), .CI(n_140));
  ADDFX1 g4786(.CO(n_202), .S(n_203), .A(n_100), .B(n_158), .CI(in_0[9]));
  ADDFX1 g4787(.CO(n_200), .S(n_201), .A(n_79), .B(n_127), .CI(n_130));
  ADDFX1 g4788(.CO(n_198), .S(n_199), .A(n_78), .B(n_126), .CI(n_122));
  ADDFX1 g4789(.CO(n_196), .S(n_197), .A(n_82), .B(n_123), .CI(in_2[9]));
  ADDFX1 g4790(.CO(n_194), .S(n_195), .A(n_34), .B(n_146), .CI(in_2[8]));
  ADDFX1 g4791(.CO(n_192), .S(n_193), .A(n_101), .B(n_142), .CI(in_4[8]));
  ADDFX1 g4792(.CO(n_190), .S(n_191), .A(n_93), .B(n_46), .CI(n_116));
  ADDFX1 g4793(.CO(n_188), .S(n_189), .A(n_125), .B(n_75), .CI(n_121));
  ADDFX1 g4794(.CO(n_186), .S(n_187), .A(n_86), .B(n_94), .CI(n_102));
  ADDFX1 g4795(.CO(n_184), .S(n_185), .A(n_97), .B(n_87), .CI(n_95));
  ADDFX1 g4796(.CO(n_182), .S(n_183), .A(n_39), .B(n_33), .CI(n_99));
  ADDFX1 g4797(.CO(n_180), .S(n_181), .A(n_36), .B(in_5[2]), .CI(n_64));
  ADDFX1 g4798(.CO(n_178), .S(n_179), .A(n_43), .B(n_41), .CI(n_28));
  ADDFX1 g4799(.CO(n_176), .S(n_177), .A(n_53), .B(n_51), .CI(n_124));
  ADDFX1 g4800(.CO(n_174), .S(n_175), .A(n_92), .B(n_74), .CI(n_73));
  ADDFX1 g4801(.CO(n_172), .S(n_173), .A(n_115), .B(in_14[8]), .CI(in_7[8]));
  ADDFX1 g4802(.CO(n_170), .S(n_171), .A(n_37), .B(n_29), .CI(n_65));
  ADDFX1 g4803(.CO(n_168), .S(n_169), .A(n_66), .B(in_0[5]), .CI(n_118));
  ADDFX1 g4804(.CO(n_166), .S(n_167), .A(n_63), .B(n_30), .CI(n_104));
  ADDFX1 g4805(.CO(n_164), .S(n_165), .A(n_114), .B(in_4[9]), .CI(in_7[9]));
  ADDFX1 g4806(.CO(n_162), .S(n_163), .A(n_67), .B(n_55), .CI(n_98));
  ADDFX1 g4807(.CO(n_160), .S(n_161), .A(n_40), .B(n_42), .CI(n_96));
  ADDFX1 g4808(.CO(n_158), .S(n_159), .A(n_69), .B(in_1[8]), .CI(in_11[8]));
  ADDFX1 g4809(.CO(n_156), .S(n_157), .A(n_15), .B(n_91), .CI(in_4[5]));
  ADDFX1 g4810(.CO(n_154), .S(n_155), .A(n_5), .B(in_15[10]), .CI(n_44));
  ADDFX1 g4811(.CO(n_152), .S(out_0[0]), .A(in_7[0]), .B(n_18), .CI(n_89));
  ADDFX1 g4812(.CO(n_150), .S(n_151), .A(n_62), .B(in_16[5]), .CI(in_5[5]));
  ADDFX1 g4813(.CO(n_148), .S(n_149), .A(n_59), .B(n_31), .CI(in_7[3]));
  ADDFX1 g4814(.CO(n_146), .S(n_147), .A(n_52), .B(in_1[7]), .CI(in_11[7]));
  ADDFX1 g4815(.CO(n_144), .S(n_145), .A(n_9), .B(in_15[10]), .CI(n_45));
  ADDFX1 g4816(.CO(n_142), .S(n_143), .A(n_77), .B(in_15[7]), .CI(in_3[7]));
  ADDFX1 g4817(.CO(n_140), .S(n_141), .A(n_72), .B(in_7[7]), .CI(in_0[7]));
  ADDFX1 g4818(.CO(n_138), .S(n_139), .A(n_38), .B(in_4[4]), .CI(n_32));
  ADDFX1 g4819(.CO(n_136), .S(n_137), .A(n_80), .B(in_1[10]), .CI(in_14[10]));
  ADDFX1 g4820(.CO(n_134), .S(n_135), .A(in_18[10]), .B(n_1), .CI(n_25));
  ADDFX1 g4821(.CO(n_132), .S(n_133), .A(n_10), .B(n_90), .CI(in_11[6]));
  ADDFX1 g4822(.CO(n_130), .S(n_131), .A(n_106), .B(in_5[8]), .CI(in_0[8]));
  ADDFX1 g4823(.CO(n_128), .S(n_129), .A(n_17), .B(n_20), .CI(n_88));
  ADDFX1 g4824(.CO(n_126), .S(n_127), .A(n_81), .B(in_8[9]), .CI(in_3[9]));
  ADDFX1 g4825(.CO(n_124), .S(n_125), .A(n_21), .B(in_6[5]), .CI(in_15[5]));
  ADDFX1 g4826(.CO(n_122), .S(n_123), .A(n_68), .B(in_6[9]), .CI(in_16[8]));
  ADDFX1 g4827(.CO(n_120), .S(n_121), .A(n_54), .B(in_7[5]), .CI(in_2[5]));
  ADDFX1 g4828(.CO(n_118), .S(n_119), .A(n_22), .B(in_11[4]), .CI(in_3[4]));
  ADDFX1 g4829(.CO(n_116), .S(n_117), .A(n_58), .B(in_5[4]), .CI(in_0[4]));
  ADDFX1 g4830(.CO(n_114), .S(n_115), .A(in_9[8]), .B(in_18[8]), .CI(n_76));
  ADDFX1 g4831(.CO(n_112), .S(n_113), .A(n_50), .B(in_5[7]), .CI(in_16[7]));
  ADDFX1 g4832(.CO(n_110), .S(n_111), .A(n_35), .B(in_4[7]), .CI(in_2[7]));
  XNOR2X1 g4833(.Y(n_109), .A(n_26), .B(in_2[13]));
  NOR2BX1 g4834(.Y(n_108), .AN(n_26), .B(in_2[13]));
  ADDFX1 g4835(.CO(n_106), .S(n_107), .A(in_10[7]), .B(in_14[7]), .CI(in_8[7]));
  ADDFX1 g4836(.CO(n_104), .S(n_105), .A(in_10[3]), .B(in_4[3]), .CI(in_16[3]));
  ADDFX1 g4837(.CO(n_102), .S(n_103), .A(n_19), .B(in_3[2]), .CI(in_4[2]));
  ADDFX1 g4838(.CO(n_100), .S(n_101), .A(in_6[8]), .B(in_8[8]), .CI(in_10[8]));
  ADDFX1 g4839(.CO(n_98), .S(n_99), .A(in_2[3]), .B(in_5[3]), .CI(in_0[3]));
  ADDFX1 g4840(.CO(n_96), .S(n_97), .A(in_1[2]), .B(in_6[2]), .CI(in_19[2]));
  ADDFX1 g4841(.CO(n_94), .S(n_95), .A(in_7[2]), .B(in_0[2]), .CI(in_16[2]));
  ADDFX1 g4842(.CO(n_92), .S(n_93), .A(in_1[5]), .B(in_10[5]), .CI(in_11[5]));
  ADDFX1 g4843(.CO(n_90), .S(n_91), .A(in_18[5]), .B(in_19[5]), .CI(in_13[5]));
  ADDFX1 g4844(.CO(n_88), .S(n_89), .A(in_0[0]), .B(in_4[0]), .CI(in_17[0]));
  ADDFX1 g4845(.CO(n_86), .S(n_87), .A(in_8[2]), .B(in_2[2]), .CI(in_11[2]));
  ADDFX1 g4846(.CO(n_84), .S(n_85), .A(in_7[6]), .B(in_16[6]), .CI(in_4[6]));
  ADDFX1 g4847(.CO(n_82), .S(n_83), .A(in_15[8]), .B(in_16[8]), .CI(in_3[8]));
  ADDFX1 g4848(.CO(n_80), .S(n_81), .A(in_13[9]), .B(in_9[9]), .CI(in_18[9]));
  ADDFX1 g4849(.CO(n_78), .S(n_79), .A(in_1[9]), .B(in_10[9]), .CI(in_11[9]));
  ADDFX1 g4850(.CO(n_76), .S(n_77), .A(in_13[7]), .B(in_17[7]), .CI(in_19[7]));
  ADDFX1 g4851(.CO(n_74), .S(n_75), .A(in_8[5]), .B(in_14[5]), .CI(in_3[5]));
  ADDFX1 g4852(.CO(n_72), .S(n_73), .A(in_6[6]), .B(in_10[6]), .CI(in_14[6]));
  ADDFX1 g4853(.CO(n_70), .S(n_71), .A(in_10[10]), .B(in_4[10]), .CI(in_0[10]));
  ADDFX1 g4854(.CO(n_68), .S(n_69), .A(in_13[8]), .B(in_17[8]), .CI(in_19[8]));
  ADDFX1 g4855(.CO(n_66), .S(n_67), .A(in_1[4]), .B(in_6[4]), .CI(in_10[4]));
  ADDFX1 g4856(.CO(n_64), .S(n_65), .A(in_0[1]), .B(in_4[1]), .CI(in_5[1]));
  ADDFX1 g4857(.CO(n_62), .S(n_63), .A(in_9[4]), .B(in_13[4]), .CI(in_18[4]));
  ADDFX1 g4858(.CO(n_60), .S(n_61), .A(in_8[6]), .B(in_15[6]), .CI(in_3[6]));
  ADDFX1 g4859(.CO(n_58), .S(n_59), .A(in_13[3]), .B(in_17[3]), .CI(in_19[3]));
  ADDFX1 g4860(.CO(n_56), .S(n_57), .A(in_14[9]), .B(in_5[9]), .CI(in_15[9]));
  ADDFX1 g4861(.CO(n_54), .S(n_55), .A(in_14[4]), .B(in_15[4]), .CI(in_8[4]));
  ADDFX1 g4862(.CO(n_52), .S(n_53), .A(in_17[6]), .B(in_19[6]), .CI(in_13[6]));
  ADDFX1 g4863(.CO(n_50), .S(n_51), .A(in_9[6]), .B(in_18[6]), .CI(in_1[6]));
  ADDFX1 g4864(.CO(n_48), .S(n_49), .A(in_5[6]), .B(in_2[6]), .CI(in_0[6]));
  ADDFX1 g4865(.CO(n_46), .S(n_47), .A(in_7[4]), .B(in_2[4]), .CI(in_16[4]));
  ADDFX1 g4866(.CO(n_44), .S(n_45), .A(in_8[10]), .B(n_8), .CI(n_7));
  ADDFX1 g4867(.CO(n_42), .S(n_43), .A(in_9[2]), .B(in_15[2]), .CI(in_14[2]));
  ADDFX1 g4868(.CO(n_40), .S(n_41), .A(in_10[2]), .B(in_17[2]), .CI(in_13[2]));
  ADDFX1 g4869(.CO(n_38), .S(n_39), .A(in_6[3]), .B(in_8[3]), .CI(in_11[3]));
  ADDFX1 g4870(.CO(n_36), .S(n_37), .A(n_2), .B(in_17[1]), .CI(in_13[1]));
  ADDFX1 g4871(.CO(n_34), .S(n_35), .A(in_9[7]), .B(in_18[7]), .CI(in_6[7]));
  ADDFX1 g4872(.CO(n_32), .S(n_33), .A(in_1[3]), .B(in_14[3]), .CI(in_3[3]));
  ADDFX1 g4873(.CO(n_30), .S(n_31), .A(in_9[3]), .B(in_18[3]), .CI(in_15[3]));
  ADDFX1 g4874(.CO(n_28), .S(n_29), .A(in_7[1]), .B(in_19[1]), .CI(in_16[1]));
  XOR2XL g4875(.Y(n_27), .A(n_12), .B(n_23));
  NAND2BX1 g4876(.Y(n_26), .AN(n_12), .B(n_23));
  XNOR2X1 g4877(.Y(n_25), .A(in_7[10]), .B(n_14));
  XNOR2X1 g4878(.Y(n_24), .A(in_7[10]), .B(n_0));
  ADDHX1 g4879(.CO(n_21), .S(n_22), .A(in_17[4]), .B(in_19[4]));
  ADDHX1 g4880(.CO(n_19), .S(n_20), .A(in_3[1]), .B(in_11[1]));
  ADDHX1 g4881(.CO(n_17), .S(n_18), .A(in_5[0]), .B(in_16[0]));
  AOI21X1 g4882(.Y(n_23), .A0(n_4), .A1(n_13), .B0(n_11));
  OAI21X1 g4883(.Y(n_16), .A0(in_18[10]), .A1(n_11), .B0(n_13));
  OAI2BB1X1 g4884(.Y(n_15), .A0N(in_17[5]), .A1N(in_9[5]), .B0(n_10));
  MXI2XL g4886(.Y(n_14), .A(n_4), .B(in_14[10]), .S0(in_6[10]));
  NAND2X1 g4888(.Y(n_13), .A(in_6[10]), .B(in_7[10]));
  NOR2X1 g4889(.Y(n_12), .A(in_8[10]), .B(in_1[10]));
  NOR2X1 g4890(.Y(n_11), .A(in_6[10]), .B(in_7[10]));
  OR2X1 g4891(.Y(n_10), .A(in_17[5]), .B(in_9[5]));
  INVX1 g4892(.Y(n_9), .A(in_11[10]));
  INVX1 g4895(.Y(n_8), .A(in_3[9]));
  INVX1 g4896(.Y(n_7), .A(in_16[8]));
  INVX1 g4897(.Y(n_6), .A(in_15[10]));
  INVX1 g4898(.Y(n_5), .A(in_10[11]));
  INVX1 g4899(.Y(n_4), .A(in_14[10]));
  BUFX2 drc_bufs(.Y(n_2), .A(in_2[1]));
  CLKXOR2X1 g2(.Y(n_1), .A(in_8[10]), .B(in_1[10]));
  XOR2XL g4901(.Y(n_0), .A(in_18[10]), .B(in_6[10]));
endmodule

module csa_tree_ADD_TC_OP_19_group_8228(in_0, in_1, in_2, in_3, in_4, in_5, in_6
    , in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, 
    in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_351, n_350, n_347, n_345, n_343, n_341, n_339, n_337, n_335, n_333, 
    n_332, n_331, n_330, n_329, n_328, n_327, n_325, n_324, n_323, n_322, 
    n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, n_312, 
    n_311, n_310, n_309, n_308, n_307, n_305, n_304, n_303, n_302, n_301, 
    n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, n_291, 
    n_290, n_289, n_288, n_286, n_285, n_284, n_283, n_282, n_281, n_280, 
    n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, 
    n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, 
    n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, 
    n_249, n_248, n_247, n_246, n_244, n_243, n_242, n_241, n_240, n_239, 
    n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, 
    n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, 
    n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, 
    n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, 
    n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, 
    n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, 
    n_168, n_167, n_166, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  OA21X1 g4693(.Y(out_0[18]), .A0(in_7[11]), .A1(n_177), .B0(n_351));
  XNOR2X1 g4694(.Y(out_0[14]), .A(n_304), .B(n_350));
  NOR2X1 g4695(.Y(n_351), .A(n_299), .B(n_350));
  ADDFX1 g4696(.CO(n_350), .S(out_0[13]), .A(n_298), .B(n_323), .CI(n_347));
  ADDFX1 g4697(.CO(n_347), .S(out_0[12]), .A(n_324), .B(n_331), .CI(n_345));
  ADDFX1 g4698(.CO(n_345), .S(out_0[11]), .A(n_329), .B(n_332), .CI(n_343));
  ADDFX1 g4699(.CO(n_343), .S(out_0[10]), .A(n_327), .B(n_330), .CI(n_341));
  ADDFX1 g4700(.CO(n_341), .S(out_0[9]), .A(n_321), .B(n_328), .CI(n_339));
  ADDFX1 g4701(.CO(n_339), .S(out_0[8]), .A(n_319), .B(n_322), .CI(n_337));
  ADDFX1 g4702(.CO(n_337), .S(out_0[7]), .A(n_317), .B(n_320), .CI(n_335));
  ADDFX1 g4703(.CO(n_335), .S(out_0[6]), .A(n_313), .B(n_318), .CI(n_333));
  ADDFX1 g4704(.CO(n_333), .S(out_0[5]), .A(n_302), .B(n_314), .CI(n_325));
  ADDFX1 g4705(.CO(n_331), .S(n_332), .A(n_296), .B(n_307), .CI(n_316));
  ADDFX1 g4706(.CO(n_329), .S(n_330), .A(n_309), .B(n_297), .CI(n_308));
  ADDFX1 g4707(.CO(n_327), .S(n_328), .A(n_291), .B(n_311), .CI(n_310));
  ADDFX1 g4708(.CO(n_325), .S(out_0[4]), .A(n_272), .B(n_303), .CI(n_305));
  ADDFX1 g4709(.CO(n_323), .S(n_324), .A(n_284), .B(n_279), .CI(n_315));
  ADDFX1 g4710(.CO(n_321), .S(n_322), .A(n_289), .B(n_294), .CI(n_312));
  ADDFX1 g4711(.CO(n_319), .S(n_320), .A(n_292), .B(n_281), .CI(n_295));
  ADDFX1 g4712(.CO(n_317), .S(n_318), .A(n_300), .B(n_277), .CI(n_293));
  ADDFX1 g4713(.CO(n_315), .S(n_316), .A(n_274), .B(n_249), .CI(n_285));
  ADDFX1 g4714(.CO(n_313), .S(n_314), .A(n_268), .B(n_261), .CI(n_301));
  ADDFX1 g4715(.CO(n_311), .S(n_312), .A(n_263), .B(n_283), .CI(n_280));
  ADDFX1 g4716(.CO(n_309), .S(n_310), .A(n_282), .B(n_265), .CI(n_288));
  ADDFX1 g4717(.CO(n_307), .S(n_308), .A(n_264), .B(n_275), .CI(n_290));
  ADDFX1 g4718(.CO(n_305), .S(out_0[3]), .A(n_257), .B(n_286), .CI(n_273));
  XNOR2X1 g4719(.Y(n_304), .A(n_183), .B(n_299));
  ADDFX1 g4720(.CO(n_302), .S(n_303), .A(n_256), .B(n_271), .CI(n_269));
  ADDFX1 g4721(.CO(n_300), .S(n_301), .A(n_270), .B(n_235), .CI(n_231));
  ADDFX1 g4722(.CO(n_299), .S(n_298), .A(n_182), .B(n_212), .CI(n_278));
  ADDFX1 g4723(.CO(n_296), .S(n_297), .A(n_237), .B(n_255), .CI(n_266));
  ADDFX1 g4724(.CO(n_294), .S(n_295), .A(n_252), .B(n_259), .CI(n_276));
  ADDFX1 g4725(.CO(n_292), .S(n_293), .A(n_227), .B(n_260), .CI(n_253));
  ADDFX1 g4726(.CO(n_290), .S(n_291), .A(n_241), .B(n_262), .CI(n_267));
  ADDFX1 g4727(.CO(n_288), .S(n_289), .A(n_246), .B(n_239), .CI(n_258));
  ADDFX1 g4728(.CO(n_286), .S(out_0[2]), .A(n_233), .B(n_244), .CI(n_251));
  ADDFX1 g4729(.CO(n_284), .S(n_285), .A(n_187), .B(n_236), .CI(n_254));
  ADDFX1 g4730(.CO(n_282), .S(n_283), .A(n_242), .B(n_215), .CI(n_159));
  ADDFX1 g4731(.CO(n_280), .S(n_281), .A(n_226), .B(n_243), .CI(n_247));
  ADDFX1 g4732(.CO(n_278), .S(n_279), .A(n_186), .B(n_248), .CI(n_213));
  ADDFX1 g4733(.CO(n_276), .S(n_277), .A(n_230), .B(n_234), .CI(n_217));
  ADDFX1 g4734(.CO(n_274), .S(n_275), .A(n_202), .B(n_240), .CI(n_225));
  ADDFX1 g4735(.CO(n_272), .S(n_273), .A(n_221), .B(n_229), .CI(n_250));
  ADDFX1 g4736(.CO(n_270), .S(n_271), .A(n_220), .B(n_126), .CI(n_195));
  ADDFX1 g4737(.CO(n_268), .S(n_269), .A(n_205), .B(n_223), .CI(n_228));
  ADDFX1 g4738(.CO(n_266), .S(n_267), .A(n_116), .B(n_211), .CI(n_219));
  ADDFX1 g4739(.CO(n_264), .S(n_265), .A(n_158), .B(n_203), .CI(n_238));
  ADDFX1 g4740(.CO(n_262), .S(n_263), .A(n_206), .B(n_200), .CI(n_185));
  ADDFX1 g4741(.CO(n_260), .S(n_261), .A(n_209), .B(n_222), .CI(n_161));
  ADDFX1 g4742(.CO(n_258), .S(n_259), .A(n_207), .B(n_201), .CI(n_216));
  ADDFX1 g4743(.CO(n_256), .S(n_257), .A(n_232), .B(n_192), .CI(n_142));
  ADDFX1 g4744(.CO(n_254), .S(n_255), .A(n_118), .B(n_218), .CI(n_144));
  ADDFX1 g4745(.CO(n_252), .S(n_253), .A(n_197), .B(n_208), .CI(n_199));
  ADDFX1 g4746(.CO(n_250), .S(n_251), .A(n_122), .B(n_190), .CI(n_193));
  ADDFX1 g4747(.CO(n_248), .S(n_249), .A(n_93), .B(n_224), .CI(n_143));
  ADDFX1 g4748(.CO(n_246), .S(n_247), .A(n_189), .B(n_198), .CI(n_53));
  ADDFX1 g4749(.CO(n_244), .S(out_0[1]), .A(n_164), .B(n_179), .CI(n_191));
  ADDFX1 g4750(.CO(n_242), .S(n_243), .A(n_131), .B(n_196), .CI(n_171));
  ADDFX1 g4751(.CO(n_240), .S(n_241), .A(n_214), .B(n_97), .CI(n_184));
  ADDFX1 g4752(.CO(n_238), .S(n_239), .A(n_188), .B(n_140), .CI(n_69));
  ADDFX1 g4753(.CO(n_236), .S(n_237), .A(n_51), .B(n_115), .CI(n_210));
  ADDFX1 g4754(.CO(n_234), .S(n_235), .A(n_163), .B(n_125), .CI(n_204));
  ADDFX1 g4755(.CO(n_232), .S(n_233), .A(n_151), .B(n_178), .CI(n_175));
  ADDFX1 g4756(.CO(n_230), .S(n_231), .A(n_37), .B(n_181), .CI(n_194));
  ADDFX1 g4757(.CO(n_228), .S(n_229), .A(n_174), .B(n_173), .CI(n_138));
  ADDFX1 g4758(.CO(n_226), .S(n_227), .A(n_162), .B(n_132), .CI(n_160));
  ADDFX1 g4759(.CO(n_224), .S(n_225), .A(n_152), .B(n_96), .CI(in_13[10]));
  ADDFX1 g4760(.CO(n_222), .S(n_223), .A(n_167), .B(n_137), .CI(n_141));
  ADDFX1 g4761(.CO(n_220), .S(n_221), .A(n_150), .B(n_124), .CI(n_121));
  ADDFX1 g4762(.CO(n_218), .S(n_219), .A(n_19), .B(n_139), .CI(in_13[9]));
  ADDFX1 g4763(.CO(n_216), .S(n_217), .A(n_180), .B(n_157), .CI(n_105));
  ADDFX1 g4764(.CO(n_214), .S(n_215), .A(n_146), .B(n_133), .CI(n_170));
  ADDFX1 g4765(.CO(n_212), .S(n_213), .A(n_119), .B(n_92), .CI(n_147));
  ADDFX1 g4766(.CO(n_210), .S(n_211), .A(n_145), .B(in_8[9]), .CI(in_7[9]));
  ADDFX1 g4767(.CO(n_208), .S(n_209), .A(n_154), .B(n_166), .CI(n_130));
  ADDFX1 g4768(.CO(n_206), .S(n_207), .A(n_127), .B(n_156), .CI(n_104));
  ADDFX1 g4769(.CO(n_204), .S(n_205), .A(n_155), .B(n_172), .CI(n_71));
  ADDFX1 g4770(.CO(n_202), .S(n_203), .A(n_153), .B(n_26), .CI(n_68));
  ADDFX1 g4771(.CO(n_200), .S(n_201), .A(n_33), .B(n_136), .CI(n_134));
  ADDFX1 g4772(.CO(n_198), .S(n_199), .A(n_149), .B(n_113), .CI(n_128));
  ADDFX1 g4773(.CO(n_196), .S(n_197), .A(n_59), .B(n_129), .CI(n_36));
  ADDFX1 g4774(.CO(n_194), .S(n_195), .A(n_123), .B(n_84), .CI(n_61));
  ADDFX1 g4775(.CO(n_192), .S(n_193), .A(n_168), .B(n_87), .CI(n_79));
  ADDFX1 g4776(.CO(n_190), .S(n_191), .A(n_63), .B(n_65), .CI(n_169));
  ADDFX1 g4777(.CO(n_188), .S(n_189), .A(n_58), .B(in_13[7]), .CI(n_148));
  ADDFX1 g4778(.CO(n_186), .S(n_187), .A(n_50), .B(n_117), .CI(n_120));
  ADDFX1 g4779(.CO(n_184), .S(n_185), .A(n_32), .B(n_135), .CI(in_16[8]));
  OR2XL g4780(.Y(n_183), .A(in_7[11]), .B(n_177));
  XOR2XL g4781(.Y(n_182), .A(n_112), .B(n_176));
  ADDFX1 g4782(.CO(n_180), .S(n_181), .A(n_89), .B(in_7[5]), .CI(n_60));
  ADDFX1 g4783(.CO(n_178), .S(n_179), .A(n_111), .B(n_101), .CI(n_91));
  NAND2BX1 g4784(.Y(n_177), .AN(n_18), .B(n_176));
  ADDFX1 g4785(.CO(n_174), .S(n_175), .A(n_62), .B(n_41), .CI(n_109));
  ADDFX1 g4786(.CO(n_172), .S(n_173), .A(n_31), .B(n_108), .CI(n_86));
  ADDFX1 g4787(.CO(n_170), .S(n_171), .A(n_95), .B(in_12[7]), .CI(in_8[7]));
  ADDFX1 g4788(.CO(n_168), .S(n_169), .A(n_12), .B(n_82), .CI(n_80));
  ADDFX1 g4789(.CO(n_166), .S(n_167), .A(n_55), .B(n_56), .CI(n_24));
  ADDFX1 g4790(.CO(n_164), .S(out_0[0]), .A(n_13), .B(n_81), .CI(n_83));
  ADDFX1 g4791(.CO(n_162), .S(n_163), .A(n_42), .B(n_72), .CI(n_70));
  ADDFX1 g4792(.CO(n_160), .S(n_161), .A(n_39), .B(n_29), .CI(n_114));
  ADDFX1 g4793(.CO(n_158), .S(n_159), .A(n_75), .B(n_52), .CI(n_27));
  ADDFX1 g4794(.CO(n_156), .S(n_157), .A(n_23), .B(n_99), .CI(in_3[6]));
  ADDFX1 g4795(.CO(n_154), .S(n_155), .A(n_30), .B(n_102), .CI(n_47));
  ADDFX1 g4796(.CO(n_152), .S(n_153), .A(n_106), .B(n_4), .CI(in_1[9]));
  ADDFX1 g4797(.CO(n_150), .S(n_151), .A(n_90), .B(n_100), .CI(n_110));
  ADDFX1 g4798(.CO(n_148), .S(n_149), .A(n_88), .B(in_10[6]), .CI(in_2[6]));
  ADDFX1 g4799(.CO(n_176), .S(n_147), .A(in_17[12]), .B(n_16), .CI(n_20));
  ADDFX1 g4800(.CO(n_145), .S(n_146), .A(n_76), .B(n_94), .CI(in_5[8]));
  ADDFX1 g4801(.CO(n_143), .S(n_144), .A(n_15), .B(n_17), .CI(in_7[10]));
  ADDFX1 g4802(.CO(n_141), .S(n_142), .A(n_78), .B(n_49), .CI(n_85));
  ADDFX1 g4803(.CO(n_139), .S(n_140), .A(n_9), .B(n_107), .CI(in_17[8]));
  ADDFX1 g4804(.CO(n_137), .S(n_138), .A(n_103), .B(n_57), .CI(n_25));
  ADDFX1 g4805(.CO(n_135), .S(n_136), .A(n_98), .B(n_22), .CI(in_10[7]));
  ADDFX1 g4806(.CO(n_133), .S(n_134), .A(n_77), .B(in_5[7]), .CI(in_2[7]));
  ADDFX1 g4807(.CO(n_131), .S(n_132), .A(n_38), .B(in_8[6]), .CI(n_28));
  ADDFX1 g4808(.CO(n_129), .S(n_130), .A(n_46), .B(n_54), .CI(in_3[5]));
  ADDFX1 g4809(.CO(n_127), .S(n_128), .A(n_34), .B(in_17[6]), .CI(in_5[6]));
  ADDFX1 g4810(.CO(n_125), .S(n_126), .A(n_43), .B(n_48), .CI(n_73));
  ADDFX1 g4811(.CO(n_123), .S(n_124), .A(n_40), .B(n_44), .CI(n_66));
  ADDFX1 g4812(.CO(n_121), .S(n_122), .A(n_67), .B(n_45), .CI(n_64));
  ADDHX1 g4813(.CO(n_119), .S(n_120), .A(in_7[11]), .B(n_21));
  ADDFX1 g4814(.CO(n_117), .S(n_118), .A(n_7), .B(in_8[10]), .CI(in_17[10]));
  ADDFX1 g4815(.CO(n_115), .S(n_116), .A(n_74), .B(in_10[9]), .CI(in_16[9]));
  ADDFX1 g4816(.CO(n_113), .S(n_114), .A(n_35), .B(in_16[5]), .CI(in_2[5]));
  NOR2X1 g4817(.Y(n_112), .A(in_7[11]), .B(n_18));
  ADDFX1 g4818(.CO(n_110), .S(n_111), .A(in_10[1]), .B(in_8[1]), .CI(in_14[1]));
  ADDFX1 g4819(.CO(n_108), .S(n_109), .A(in_0[2]), .B(in_7[2]), .CI(in_8[2]));
  ADDFX1 g4820(.CO(n_106), .S(n_107), .A(in_0[8]), .B(in_11[8]), .CI(in_15[8]));
  ADDFX1 g4821(.CO(n_104), .S(n_105), .A(in_13[6]), .B(in_7[6]), .CI(in_16[6]));
  ADDFX1 g4822(.CO(n_102), .S(n_103), .A(in_0[3]), .B(in_6[3]), .CI(in_15[3]));
  ADDFX1 g4823(.CO(n_100), .S(n_101), .A(in_13[1]), .B(in_16[1]), .CI(in_17[1]));
  ADDFX1 g4824(.CO(n_98), .S(n_99), .A(in_0[6]), .B(in_6[6]), .CI(in_15[6]));
  ADDFX1 g4825(.CO(n_96), .S(n_97), .A(n_11), .B(in_3[9]), .CI(in_17[9]));
  ADDFX1 g4826(.CO(n_94), .S(n_95), .A(in_0[7]), .B(in_6[7]), .CI(in_15[7]));
  ADDFX1 g4827(.CO(n_92), .S(n_93), .A(n_14), .B(in_17[11]), .CI(in_13[11]));
  ADDFX1 g4828(.CO(n_90), .S(n_91), .A(in_11[1]), .B(in_0[1]), .CI(in_3[1]));
  ADDFX1 g4829(.CO(n_88), .S(n_89), .A(in_0[5]), .B(in_6[5]), .CI(in_15[5]));
  ADDFX1 g4830(.CO(n_86), .S(n_87), .A(in_16[2]), .B(in_13[2]), .CI(in_10[2]));
  ADDFX1 g4831(.CO(n_84), .S(n_85), .A(in_5[3]), .B(in_2[3]), .CI(in_16[3]));
  ADDFX1 g4832(.CO(n_82), .S(n_83), .A(in_6[0]), .B(in_8[0]), .CI(in_16[0]));
  ADDFX1 g4833(.CO(n_80), .S(n_81), .A(in_5[0]), .B(in_13[0]), .CI(in_11[0]));
  ADDFX1 g4834(.CO(n_78), .S(n_79), .A(in_3[2]), .B(in_2[2]), .CI(in_5[2]));
  ADDFX1 g4835(.CO(n_76), .S(n_77), .A(in_4[7]), .B(in_11[7]), .CI(in_19[7]));
  ADDFX1 g4836(.CO(n_74), .S(n_75), .A(in_14[8]), .B(in_12[8]), .CI(in_1[8]));
  ADDFX1 g4837(.CO(n_72), .S(n_73), .A(in_5[4]), .B(in_3[4]), .CI(in_8[4]));
  ADDFX1 g4838(.CO(n_70), .S(n_71), .A(in_7[4]), .B(in_2[4]), .CI(in_16[4]));
  ADDFX1 g4839(.CO(n_68), .S(n_69), .A(in_8[8]), .B(in_13[8]), .CI(in_7[8]));
  ADDFX1 g4840(.CO(n_66), .S(n_67), .A(in_1[2]), .B(in_6[2]), .CI(in_15[2]));
  ADDFX1 g4841(.CO(n_64), .S(n_65), .A(in_7[1]), .B(in_2[1]), .CI(in_5[1]));
  ADDFX1 g4842(.CO(n_62), .S(n_63), .A(in_4[1]), .B(in_6[1]), .CI(in_19[1]));
  ADDFX1 g4843(.CO(n_60), .S(n_61), .A(in_17[4]), .B(in_13[4]), .CI(in_10[4]));
  ADDFX1 g4844(.CO(n_58), .S(n_59), .A(in_14[6]), .B(in_1[6]), .CI(in_12[6]));
  ADDFX1 g4845(.CO(n_56), .S(n_57), .A(in_14[3]), .B(in_17[3]), .CI(in_12[3]));
  ADDFX1 g4846(.CO(n_54), .S(n_55), .A(in_0[4]), .B(in_11[4]), .CI(in_19[4]));
  ADDFX1 g4847(.CO(n_52), .S(n_53), .A(in_3[7]), .B(in_7[7]), .CI(in_16[7]));
  ADDFX1 g4848(.CO(n_50), .S(n_51), .A(n_3), .B(in_16[10]), .CI(n_5));
  ADDFX1 g4849(.CO(n_48), .S(n_49), .A(in_3[3]), .B(in_13[3]), .CI(in_8[3]));
  ADDFX1 g4850(.CO(n_46), .S(n_47), .A(in_6[4]), .B(in_14[4]), .CI(in_15[4]));
  ADDFX1 g4851(.CO(n_44), .S(n_45), .A(in_14[2]), .B(in_17[2]), .CI(in_19[2]));
  ADDFX1 g4852(.CO(n_42), .S(n_43), .A(n_2), .B(in_1[4]), .CI(in_12[4]));
  ADDFX1 g4853(.CO(n_40), .S(n_41), .A(in_4[2]), .B(in_11[2]), .CI(in_12[2]));
  ADDFX1 g4854(.CO(n_38), .S(n_39), .A(in_4[4]), .B(in_1[5]), .CI(in_10[5]));
  ADDFX1 g4855(.CO(n_36), .S(n_37), .A(in_5[5]), .B(in_8[5]), .CI(in_13[5]));
  ADDFX1 g4856(.CO(n_34), .S(n_35), .A(in_4[5]), .B(in_11[5]), .CI(in_19[5]));
  ADDFX1 g4857(.CO(n_32), .S(n_33), .A(in_14[7]), .B(in_1[7]), .CI(in_17[7]));
  ADDFX1 g4858(.CO(n_30), .S(n_31), .A(in_4[3]), .B(in_11[3]), .CI(in_19[3]));
  ADDFX1 g4859(.CO(n_28), .S(n_29), .A(in_14[5]), .B(in_12[5]), .CI(in_17[5]));
  ADDFX1 g4860(.CO(n_26), .S(n_27), .A(in_2[8]), .B(in_10[8]), .CI(in_3[8]));
  ADDFX1 g4861(.CO(n_24), .S(n_25), .A(in_7[3]), .B(in_1[3]), .CI(in_10[3]));
  ADDFX1 g4862(.CO(n_22), .S(n_23), .A(in_11[6]), .B(in_4[6]), .CI(in_19[6]));
  OAI21X1 g4863(.Y(n_21), .A0(in_12[10]), .A1(n_10), .B0(n_16));
  AO21XL g4864(.Y(n_20), .A0(in_7[11]), .A1(n_8), .B0(n_18));
  OAI2BB1X1 g4865(.Y(n_19), .A0N(n_6), .A1N(in_12[9]), .B0(n_17));
  NOR2XL g4866(.Y(n_18), .A(in_7[11]), .B(n_8));
  OR2X1 g4867(.Y(n_17), .A(n_6), .B(in_12[9]));
  NAND2X1 g4868(.Y(n_16), .A(in_12[10]), .B(n_10));
  ADDHX1 g4869(.CO(n_14), .S(n_15), .A(in_12[10]), .B(in_1[10]));
  ADDHX1 g4870(.CO(n_12), .S(n_13), .A(n_0), .B(in_7[0]));
  XNOR2X1 g4871(.Y(n_11), .A(in_15[9]), .B(in_5[8]));
  XNOR2X1 g4872(.Y(n_10), .A(in_1[10]), .B(in_16[10]));
  XNOR2X1 g4873(.Y(n_9), .A(in_4[8]), .B(in_19[8]));
  NOR2X1 g4874(.Y(n_8), .A(in_1[10]), .B(in_16[10]));
  NOR2BX1 g4875(.Y(n_7), .AN(in_15[9]), .B(in_5[8]));
  OR2XL g4876(.Y(n_6), .A(in_19[8]), .B(in_4[8]));
  INVX1 g4877(.Y(n_5), .A(in_10[10]));
  INVX1 g4878(.Y(n_4), .A(in_2[9]));
  INVX1 g4879(.Y(n_3), .A(in_3[9]));
  INVX1 g4880(.Y(n_2), .A(in_4[4]));
  BUFX2 drc_bufs(.Y(n_0), .A(in_2[0]));
endmodule

module csa_tree_ADD_TC_OP_19_group_6301(in_0, in_1, in_2, in_3, in_4, in_5, in_6
    , in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, 
    in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_332, n_330, n_328, n_326, n_324, n_322, n_320, n_318, n_316, n_314, 
    n_313, n_312, n_311, n_310, n_309, n_308, n_306, n_305, n_304, n_303, 
    n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_292, 
    n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, n_282, 
    n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, 
    n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, 
    n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, 
    n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, 
    n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, 
    n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, 
    n_220, n_219, n_218, n_216, n_215, n_214, n_213, n_212, n_211, n_210, 
    n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, 
    n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, 
    n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, 
    n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, 
    n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, 
    n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, 
    n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  AOI21X2 g4206(.Y(out_0[18]), .A0(n_13), .A1(n_180), .B0(n_332));
  ADDFX1 g4207(.CO(n_332), .S(out_0[14]), .A(n_189), .B(n_274), .CI(n_330));
  ADDFX1 g4208(.CO(n_330), .S(out_0[13]), .A(n_275), .B(n_298), .CI(n_328));
  ADDFX1 g4209(.CO(n_328), .S(out_0[12]), .A(n_312), .B(n_299), .CI(n_326));
  ADDFX1 g4210(.CO(n_326), .S(out_0[11]), .A(n_310), .B(n_313), .CI(n_324));
  ADDFX1 g4211(.CO(n_324), .S(out_0[10]), .A(n_302), .B(n_311), .CI(n_322));
  ADDFX1 g4212(.CO(n_322), .S(out_0[9]), .A(n_300), .B(n_303), .CI(n_320));
  ADDFX1 g4213(.CO(n_320), .S(out_0[8]), .A(n_308), .B(n_301), .CI(n_318));
  ADDFX1 g4214(.CO(n_318), .S(out_0[7]), .A(n_304), .B(n_309), .CI(n_316));
  ADDFX1 g4215(.CO(n_316), .S(out_0[6]), .A(n_290), .B(n_305), .CI(n_314));
  ADDFX1 g4216(.CO(n_314), .S(out_0[5]), .A(n_280), .B(n_291), .CI(n_306));
  ADDFX1 g4217(.CO(n_312), .S(n_313), .A(n_267), .B(n_295), .CI(n_296));
  ADDFX1 g4218(.CO(n_310), .S(n_311), .A(n_276), .B(n_286), .CI(n_297));
  ADDFX1 g4219(.CO(n_308), .S(n_309), .A(n_259), .B(n_288), .CI(n_283));
  ADDFX1 g4220(.CO(n_306), .S(out_0[4]), .A(n_268), .B(n_292), .CI(n_281));
  ADDFX1 g4221(.CO(n_304), .S(n_305), .A(n_272), .B(n_251), .CI(n_289));
  ADDFX1 g4222(.CO(n_302), .S(n_303), .A(n_277), .B(n_284), .CI(n_287));
  ADDFX1 g4223(.CO(n_300), .S(n_301), .A(n_282), .B(n_271), .CI(n_285));
  ADDFX1 g4224(.CO(n_298), .S(n_299), .A(n_266), .B(n_294), .CI(n_257));
  ADDFX1 g4225(.CO(n_296), .S(n_297), .A(n_248), .B(n_231), .CI(n_279));
  ADDFX1 g4226(.CO(n_294), .S(n_295), .A(n_230), .B(n_225), .CI(n_278));
  ADDFX1 g4227(.CO(n_292), .S(out_0[3]), .A(n_233), .B(n_260), .CI(n_269));
  ADDFX1 g4228(.CO(n_290), .S(n_291), .A(n_262), .B(n_265), .CI(n_273));
  ADDFX1 g4229(.CO(n_288), .S(n_289), .A(n_203), .B(n_264), .CI(n_255));
  ADDFX1 g4230(.CO(n_286), .S(n_287), .A(n_239), .B(n_270), .CI(n_249));
  ADDFX1 g4231(.CO(n_284), .S(n_285), .A(n_245), .B(n_258), .CI(n_247));
  ADDFX1 g4232(.CO(n_282), .S(n_283), .A(n_254), .B(n_253), .CI(n_250));
  ADDFX1 g4233(.CO(n_280), .S(n_281), .A(n_232), .B(n_237), .CI(n_263));
  ADDFX1 g4234(.CO(n_278), .S(n_279), .A(n_240), .B(n_243), .CI(n_238));
  ADDFX1 g4235(.CO(n_276), .S(n_277), .A(n_241), .B(n_244), .CI(n_246));
  ADDFX1 g4236(.CO(n_274), .S(n_275), .A(n_179), .B(n_196), .CI(n_256));
  ADDFX1 g4237(.CO(n_272), .S(n_273), .A(n_236), .B(n_213), .CI(n_211));
  ADDFX1 g4238(.CO(n_270), .S(n_271), .A(n_234), .B(n_221), .CI(n_252));
  ADDFX1 g4239(.CO(n_268), .S(n_269), .A(n_204), .B(n_219), .CI(n_226));
  ADDFX1 g4240(.CO(n_266), .S(n_267), .A(n_182), .B(n_137), .CI(n_242));
  ADDFX1 g4241(.CO(n_264), .S(n_265), .A(n_194), .B(n_228), .CI(n_223));
  ADDFX1 g4242(.CO(n_262), .S(n_263), .A(n_218), .B(n_195), .CI(n_229));
  ADDFX1 g4243(.CO(n_260), .S(out_0[2]), .A(n_205), .B(n_216), .CI(n_227));
  ADDFX1 g4244(.CO(n_258), .S(n_259), .A(n_214), .B(n_209), .CI(n_235));
  ADDFX1 g4245(.CO(n_256), .S(n_257), .A(n_181), .B(n_197), .CI(n_224));
  ADDFX1 g4246(.CO(n_254), .S(n_255), .A(n_153), .B(n_188), .CI(n_222));
  ADDFX1 g4247(.CO(n_252), .S(n_253), .A(n_207), .B(n_202), .CI(n_193));
  ADDFX1 g4248(.CO(n_250), .S(n_251), .A(n_212), .B(n_210), .CI(n_215));
  ADDFX1 g4249(.CO(n_248), .S(n_249), .A(n_191), .B(n_220), .CI(n_201));
  ADDFX1 g4250(.CO(n_246), .S(n_247), .A(n_206), .B(n_199), .CI(n_208));
  ADDFX1 g4251(.CO(n_244), .S(n_245), .A(n_192), .B(n_186), .CI(n_124));
  ADDFX1 g4252(.CO(n_242), .S(n_243), .A(n_200), .B(n_177), .CI(n_190));
  ADDFX1 g4253(.CO(n_240), .S(n_241), .A(n_125), .B(n_185), .CI(n_45));
  ADDFX1 g4254(.CO(n_238), .S(n_239), .A(n_123), .B(n_198), .CI(n_178));
  ADDFX1 g4255(.CO(n_236), .S(n_237), .A(n_150), .B(n_148), .CI(n_183));
  ADDFX1 g4256(.CO(n_234), .S(n_235), .A(n_175), .B(n_187), .CI(n_136));
  ADDFX1 g4257(.CO(n_232), .S(n_233), .A(n_165), .B(n_174), .CI(n_184));
  ADDFX1 g4258(.CO(n_230), .S(n_231), .A(n_168), .B(n_144), .CI(n_138));
  ADDFX1 g4259(.CO(n_228), .S(n_229), .A(n_122), .B(n_173), .CI(n_170));
  ADDFX1 g4260(.CO(n_226), .S(n_227), .A(n_172), .B(n_166), .CI(n_161));
  ADDFX1 g4261(.CO(n_224), .S(n_225), .A(n_167), .B(n_143), .CI(n_120));
  ADDFX1 g4262(.CO(n_222), .S(n_223), .A(n_121), .B(n_169), .CI(n_51));
  ADDFX1 g4263(.CO(n_220), .S(n_221), .A(n_151), .B(n_126), .CI(n_134));
  ADDFX1 g4264(.CO(n_218), .S(n_219), .A(n_171), .B(n_118), .CI(n_146));
  ADDFX1 g4265(.CO(n_216), .S(out_0[1]), .A(n_141), .B(n_164), .CI(n_162));
  ADDFX1 g4266(.CO(n_214), .S(n_215), .A(n_155), .B(n_108), .CI(n_176));
  ADDFX1 g4267(.CO(n_212), .S(n_213), .A(n_149), .B(n_156), .CI(n_114));
  ADDFX1 g4268(.CO(n_210), .S(n_211), .A(n_147), .B(n_154), .CI(n_140));
  ADDFX1 g4269(.CO(n_208), .S(n_209), .A(n_152), .B(n_89), .CI(n_91));
  ADDFX1 g4270(.CO(n_206), .S(n_207), .A(n_157), .B(in_1[7]), .CI(n_96));
  ADDFX1 g4271(.CO(n_204), .S(n_205), .A(n_163), .B(n_79), .CI(n_116));
  ADDFX1 g4272(.CO(n_202), .S(n_203), .A(n_139), .B(n_97), .CI(n_128));
  ADDFX1 g4273(.CO(n_200), .S(n_201), .A(n_85), .B(n_101), .CI(n_133));
  ADDFX1 g4274(.CO(n_198), .S(n_199), .A(n_132), .B(n_90), .CI(n_135));
  ADDFX1 g4275(.CO(n_196), .S(n_197), .A(n_111), .B(n_119), .CI(n_130));
  ADDFX1 g4276(.CO(n_194), .S(n_195), .A(n_117), .B(n_145), .CI(n_43));
  ADDFX1 g4277(.CO(n_192), .S(n_193), .A(n_160), .B(n_107), .CI(n_127));
  ADDFX1 g4278(.CO(n_190), .S(n_191), .A(n_80), .B(n_131), .CI(in_11[9]));
  XOR2XL g4279(.Y(n_189), .A(n_13), .B(n_180));
  ADDFX1 g4280(.CO(n_187), .S(n_188), .A(n_53), .B(n_158), .CI(n_50));
  ADDFX1 g4281(.CO(n_185), .S(n_186), .A(n_159), .B(n_88), .CI(in_2[8]));
  ADDFX1 g4282(.CO(n_183), .S(n_184), .A(n_115), .B(n_71), .CI(n_110));
  ADDFX1 g4283(.CO(n_181), .S(n_182), .A(n_93), .B(n_112), .CI(n_98));
  ADDFX1 g4284(.CO(n_180), .S(n_179), .A(n_24), .B(n_23), .CI(n_129));
  ADDFX1 g4285(.CO(n_177), .S(n_178), .A(n_106), .B(in_2[9]), .CI(in_10[9]));
  ADDFX1 g4286(.CO(n_175), .S(n_176), .A(n_102), .B(n_62), .CI(n_113));
  ADDFX1 g4287(.CO(n_173), .S(n_174), .A(n_83), .B(n_78), .CI(n_26));
  ADDFX1 g4288(.CO(n_171), .S(n_172), .A(n_74), .B(n_77), .CI(n_37));
  ADDFX1 g4289(.CO(n_169), .S(n_170), .A(n_82), .B(n_65), .CI(in_11[4]));
  ADDFX1 g4290(.CO(n_167), .S(n_168), .A(n_69), .B(n_84), .CI(in_2[10]));
  ADDFX1 g4291(.CO(n_165), .S(n_166), .A(n_30), .B(n_94), .CI(n_87));
  ADDFX1 g4292(.CO(n_163), .S(n_164), .A(n_31), .B(n_27), .CI(n_75));
  ADDFX1 g4293(.CO(n_161), .S(n_162), .A(n_47), .B(n_38), .CI(n_95));
  ADDFX1 g4294(.CO(n_159), .S(n_160), .A(n_58), .B(n_60), .CI(in_13[7]));
  ADDFX1 g4295(.CO(n_157), .S(n_158), .A(n_56), .B(n_33), .CI(in_19[6]));
  ADDFX1 g4296(.CO(n_155), .S(n_156), .A(n_34), .B(n_57), .CI(n_42));
  ADDFX1 g4297(.CO(n_153), .S(n_154), .A(n_104), .B(n_103), .CI(n_63));
  ADDFX1 g4298(.CO(n_151), .S(n_152), .A(n_36), .B(n_40), .CI(in_16[7]));
  ADDFX1 g4299(.CO(n_149), .S(n_150), .A(n_55), .B(n_25), .CI(n_109));
  ADDFX1 g4300(.CO(n_147), .S(n_148), .A(n_49), .B(n_70), .CI(n_105));
  ADDFX1 g4301(.CO(n_145), .S(n_146), .A(n_29), .B(n_73), .CI(n_86));
  ADDFX1 g4302(.CO(n_143), .S(n_144), .A(n_15), .B(n_100), .CI(in_11[10]));
  ADDFX1 g4303(.CO(n_141), .S(out_0[0]), .A(n_17), .B(n_32), .CI(n_28));
  ADDFX1 g4304(.CO(n_139), .S(n_140), .A(n_48), .B(n_64), .CI(in_11[5]));
  ADDFX1 g4305(.CO(n_137), .S(n_138), .A(n_44), .B(n_67), .CI(n_99));
  ADDFX1 g4306(.CO(n_135), .S(n_136), .A(n_52), .B(in_5[7]), .CI(in_11[7]));
  ADDFX1 g4307(.CO(n_133), .S(n_134), .A(n_41), .B(in_1[8]), .CI(in_5[8]));
  ADDFX1 g4308(.CO(n_131), .S(n_132), .A(n_35), .B(in_19[8]), .CI(in_13[8]));
  ADDFX1 g4309(.CO(n_129), .S(n_130), .A(n_92), .B(n_1), .CI(in_11[12]));
  ADDFX1 g4310(.CO(n_127), .S(n_128), .A(n_61), .B(in_10[6]), .CI(in_2[6]));
  ADDFX1 g4311(.CO(n_125), .S(n_126), .A(n_39), .B(in_12[8]), .CI(in_10[8]));
  ADDFX1 g4312(.CO(n_123), .S(n_124), .A(n_12), .B(n_81), .CI(in_11[8]));
  ADDFX1 g4313(.CO(n_121), .S(n_122), .A(n_72), .B(in_10[4]), .CI(in_2[4]));
  ADDFX1 g4314(.CO(n_119), .S(n_120), .A(n_14), .B(n_66), .CI(in_11[11]));
  ADDFX1 g4315(.CO(n_117), .S(n_118), .A(n_18), .B(n_76), .CI(in_12[3]));
  ADDFX1 g4316(.CO(n_115), .S(n_116), .A(n_19), .B(n_46), .CI(in_10[2]));
  ADDFX1 g4317(.CO(n_113), .S(n_114), .A(n_54), .B(in_1[5]), .CI(in_12[5]));
  ADDFX1 g4318(.CO(n_111), .S(n_112), .A(in_19[10]), .B(n_11), .CI(in_2[11]));
  ADDFX1 g4319(.CO(n_109), .S(n_110), .A(n_21), .B(in_5[3]), .CI(in_1[3]));
  ADDFX1 g4320(.CO(n_107), .S(n_108), .A(n_59), .B(in_12[6]), .CI(in_1[6]));
  OAI2BB1X1 g4321(.Y(n_106), .A0N(n_68), .A1N(in_19[9]), .B0(n_69));
  ADDFX1 g4322(.CO(n_104), .S(n_105), .A(n_5), .B(n_20), .CI(in_19[4]));
  ADDFX1 g4323(.CO(n_102), .S(n_103), .A(in_16[5]), .B(in_17[5]), .CI(in_19[5]));
  ADDFX1 g4324(.CO(n_100), .S(n_101), .A(in_0[9]), .B(n_9), .CI(in_13[9]));
  ADDFX1 g4325(.CO(n_98), .S(n_99), .A(n_4), .B(in_1[10]), .CI(in_10[10]));
  ADDFX1 g4326(.CO(n_96), .S(n_97), .A(in_7[6]), .B(in_5[6]), .CI(in_11[6]));
  ADDFX1 g4327(.CO(n_94), .S(n_95), .A(n_16), .B(in_11[1]), .CI(in_1[1]));
  ADDFX1 g4328(.CO(n_92), .S(n_93), .A(in_16[11]), .B(in_17[11]), .CI(n_7));
  ADDFX1 g4329(.CO(n_90), .S(n_91), .A(in_12[7]), .B(in_2[7]), .CI(in_10[7]));
  ADDFX1 g4330(.CO(n_88), .S(n_89), .A(in_17[7]), .B(in_19[7]), .CI(in_7[7]));
  ADDFX1 g4331(.CO(n_86), .S(n_87), .A(in_8[2]), .B(in_5[2]), .CI(in_11[2]));
  ADDFX1 g4332(.CO(n_84), .S(n_85), .A(in_17[9]), .B(in_7[9]), .CI(in_16[9]));
  ADDFX1 g4333(.CO(n_82), .S(n_83), .A(in_8[3]), .B(in_18[3]), .CI(in_15[3]));
  ADDFX1 g4334(.CO(n_80), .S(n_81), .A(in_16[8]), .B(in_17[8]), .CI(in_7[8]));
  ADDFX1 g4335(.CO(n_78), .S(n_79), .A(in_2[2]), .B(in_1[2]), .CI(in_12[2]));
  ADDFX1 g4336(.CO(n_76), .S(n_77), .A(in_3[2]), .B(in_0[2]), .CI(in_13[2]));
  ADDFX1 g4337(.CO(n_74), .S(n_75), .A(in_3[1]), .B(in_18[1]), .CI(in_8[1]));
  ADDFX1 g4338(.CO(n_72), .S(n_73), .A(in_0[3]), .B(in_14[3]), .CI(in_16[3]));
  ADDFX1 g4339(.CO(n_70), .S(n_71), .A(in_2[3]), .B(in_10[3]), .CI(in_11[3]));
  OR2X1 g4340(.Y(n_69), .A(n_68), .B(in_19[9]));
  ADDFX1 g4341(.CO(n_66), .S(n_67), .A(in_16[10]), .B(in_13[10]), .CI(in_5[10]));
  ADDFX1 g4342(.CO(n_64), .S(n_65), .A(in_0[4]), .B(in_8[4]), .CI(in_7[4]));
  ADDFX1 g4343(.CO(n_62), .S(n_63), .A(in_18[4]), .B(in_13[5]), .CI(in_7[5]));
  ADDFX1 g4344(.CO(n_60), .S(n_61), .A(in_8[6]), .B(in_0[6]), .CI(in_14[6]));
  ADDFX1 g4345(.CO(n_58), .S(n_59), .A(in_3[6]), .B(in_15[6]), .CI(in_18[6]));
  ADDFX1 g4346(.CO(n_56), .S(n_57), .A(in_3[5]), .B(in_15[5]), .CI(in_18[5]));
  ADDFX1 g4347(.CO(n_54), .S(n_55), .A(in_3[4]), .B(in_14[4]), .CI(in_15[4]));
  ADDFX1 g4348(.CO(n_52), .S(n_53), .A(in_16[6]), .B(in_17[6]), .CI(in_13[6]));
  ADDFX1 g4349(.CO(n_50), .S(n_51), .A(in_5[5]), .B(in_2[5]), .CI(in_10[5]));
  ADDFX1 g4350(.CO(n_48), .S(n_49), .A(in_16[4]), .B(in_17[4]), .CI(in_13[4]));
  ADDFX1 g4351(.CO(n_46), .S(n_47), .A(in_5[1]), .B(in_2[1]), .CI(in_15[1]));
  ADDFX1 g4352(.CO(n_44), .S(n_45), .A(in_12[9]), .B(in_1[9]), .CI(in_5[9]));
  ADDFX1 g4353(.CO(n_42), .S(n_43), .A(in_5[4]), .B(in_1[4]), .CI(in_12[4]));
  ADDFX1 g4354(.CO(n_68), .S(n_41), .A(in_8[8]), .B(in_0[8]), .CI(in_15[8]));
  ADDFX1 g4355(.CO(n_39), .S(n_40), .A(in_0[7]), .B(in_8[7]), .CI(n_6));
  ADDFX1 g4356(.CO(n_37), .S(n_38), .A(in_14[1]), .B(in_10[1]), .CI(in_12[1]));
  ADDFX1 g4357(.CO(n_35), .S(n_36), .A(in_14[7]), .B(in_15[7]), .CI(in_18[7]));
  ADDFX1 g4358(.CO(n_33), .S(n_34), .A(in_8[5]), .B(in_0[5]), .CI(in_14[5]));
  ADDFX1 g4359(.CO(n_31), .S(n_32), .A(n_2), .B(in_3[0]), .CI(in_11[0]));
  ADDFX1 g4360(.CO(n_29), .S(n_30), .A(in_7[2]), .B(in_18[2]), .CI(in_15[2]));
  ADDFX1 g4361(.CO(n_27), .S(n_28), .A(in_1[0]), .B(in_10[0]), .CI(in_18[0]));
  ADDFX1 g4362(.CO(n_25), .S(n_26), .A(in_13[3]), .B(in_7[3]), .CI(in_19[3]));
  OAI2BB1X1 g4363(.Y(n_24), .A0N(in_16[11]), .A1N(in_17[12]), .B0(n_22));
  XNOR2X1 g4365(.Y(n_23), .A(n_0), .B(in_11[13]));
  OAI21XL g4366(.Y(n_22), .A0(in_16[11]), .A1(in_17[12]), .B0(n_8));
  ADDHX1 g4368(.CO(n_20), .S(n_21), .A(in_3[3]), .B(in_17[3]));
  ADDHX1 g4369(.CO(n_18), .S(n_19), .A(in_14[2]), .B(in_19[2]));
  ADDHX1 g4370(.CO(n_16), .S(n_17), .A(in_5[0]), .B(in_12[0]));
  ADDHX1 g4371(.CO(n_14), .S(n_15), .A(in_7[10]), .B(in_17[10]));
  OAI22X1 g4372(.Y(n_13), .A0(in_17[12]), .A1(n_10), .B0(in_16[11]), .B1(
    in_11[13]));
  OAI2BB1X1 g4373(.Y(n_12), .A0N(in_14[8]), .A1N(in_3[7]), .B0(n_9));
  MXI2XL g4374(.Y(n_11), .A(n_4), .B(in_19[10]), .S0(in_7[10]));
  AND2XL g4376(.Y(n_10), .A(in_16[11]), .B(in_11[13]));
  OR2X1 g4377(.Y(n_9), .A(in_14[8]), .B(in_3[7]));
  NOR2X1 g4378(.Y(n_8), .A(in_19[10]), .B(in_7[10]));
  INVX1 g4379(.Y(n_7), .A(in_13[11]));
  INVX1 g4380(.Y(n_6), .A(in_3[7]));
  INVX1 g4381(.Y(n_5), .A(in_18[4]));
  INVX1 g4383(.Y(n_4), .A(in_19[10]));
  BUFX2 drc_bufs(.Y(n_2), .A(in_2[0]));
  CLKXOR2X1 g2(.Y(n_1), .A(n_8), .B(n_0));
  XOR2XL g4384(.Y(n_0), .A(in_16[11]), .B(in_17[12]));
endmodule

module csa_tree_ADD_TC_OP_19_group_4361(in_0, in_1, in_2, in_3, in_4, in_5, in_6
    , in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, 
    in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_357, n_355, n_353, n_351, n_349, n_347, n_345, n_343, n_341, n_339, 
    n_337, n_336, n_335, n_334, n_333, n_332, n_331, n_330, n_329, n_328, 
    n_327, n_325, n_324, n_323, n_322, n_321, n_320, n_319, n_318, n_317, 
    n_316, n_315, n_313, n_312, n_311, n_310, n_309, n_308, n_307, n_306, 
    n_305, n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, 
    n_295, n_294, n_293, n_292, n_290, n_289, n_288, n_287, n_286, n_285, 
    n_284, n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, 
    n_274, n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, 
    n_264, n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, 
    n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, 
    n_223, n_222, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, 
    n_213, n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, 
    n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 
    n_193, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, 
    n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, 
    n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, 
    n_162, n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, 
    n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
    n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
    n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, 
    n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, 
    n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
    n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, 
    n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
    n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  OR2X1 g4518(.Y(out_0[18]), .A(n_292), .B(n_357));
  AOI21X1 g4519(.Y(n_357), .A0(n_102), .A1(n_287), .B0(n_355));
  ADDFX1 g4520(.CO(n_355), .S(out_0[14]), .A(n_286), .B(n_319), .CI(n_353));
  ADDFX1 g4521(.CO(n_353), .S(out_0[13]), .A(n_320), .B(n_331), .CI(n_351));
  ADDFX1 g4522(.CO(n_351), .S(out_0[12]), .A(n_329), .B(n_332), .CI(n_349));
  ADDFX1 g4523(.CO(n_349), .S(out_0[11]), .A(n_335), .B(n_330), .CI(n_347));
  ADDFX1 g4524(.CO(n_347), .S(out_0[10]), .A(n_333), .B(n_336), .CI(n_345));
  ADDFX1 g4525(.CO(n_345), .S(out_0[9]), .A(n_327), .B(n_334), .CI(n_343));
  ADDFX1 g4526(.CO(n_343), .S(out_0[8]), .A(n_321), .B(n_328), .CI(n_341));
  ADDFX1 g4527(.CO(n_341), .S(out_0[7]), .A(n_323), .B(n_322), .CI(n_339));
  ADDFX1 g4528(.CO(n_339), .S(out_0[6]), .A(n_311), .B(n_337), .CI(n_324));
  ADDFX1 g4529(.CO(n_337), .S(out_0[5]), .A(n_299), .B(n_312), .CI(n_325));
  ADDFX1 g4530(.CO(n_335), .S(n_336), .A(n_294), .B(n_317), .CI(n_316));
  ADDFX1 g4531(.CO(n_333), .S(n_334), .A(n_288), .B(n_309), .CI(n_318));
  ADDFX1 g4532(.CO(n_331), .S(n_332), .A(n_282), .B(n_307), .CI(n_306));
  ADDFX1 g4533(.CO(n_329), .S(n_330), .A(n_283), .B(n_315), .CI(n_308));
  ADDFX1 g4534(.CO(n_327), .S(n_328), .A(n_301), .B(n_289), .CI(n_310));
  ADDFX1 g4535(.CO(n_325), .S(out_0[4]), .A(n_278), .B(n_313), .CI(n_300));
  ADDFX1 g4536(.CO(n_323), .S(n_324), .A(n_297), .B(n_265), .CI(n_296));
  ADDFX1 g4537(.CO(n_321), .S(n_322), .A(n_295), .B(n_285), .CI(n_302));
  ADDFX1 g4538(.CO(n_319), .S(n_320), .A(n_276), .B(n_267), .CI(n_305));
  ADDFX1 g4539(.CO(n_317), .S(n_318), .A(n_253), .B(n_255), .CI(n_304));
  ADDFX1 g4540(.CO(n_315), .S(n_316), .A(n_254), .B(n_275), .CI(n_303));
  ADDFX1 g4541(.CO(n_313), .S(out_0[3]), .A(n_249), .B(n_279), .CI(n_290));
  ADDFX1 g4542(.CO(n_311), .S(n_312), .A(n_262), .B(n_273), .CI(n_298));
  ADDFX1 g4543(.CO(n_309), .S(n_310), .A(n_281), .B(n_201), .CI(n_284));
  ADDFX1 g4544(.CO(n_307), .S(n_308), .A(n_269), .B(n_274), .CI(n_293));
  ADDFX1 g4545(.CO(n_305), .S(n_306), .A(n_196), .B(n_268), .CI(n_277));
  ADDFX1 g4546(.CO(n_303), .S(n_304), .A(n_280), .B(n_229), .CI(n_200));
  ADDFX1 g4547(.CO(n_301), .S(n_302), .A(n_260), .B(n_264), .CI(n_271));
  ADDFX1 g4548(.CO(n_299), .S(n_300), .A(n_248), .B(n_259), .CI(n_263));
  ADDFX1 g4549(.CO(n_297), .S(n_298), .A(n_226), .B(n_258), .CI(n_241));
  ADDFX1 g4550(.CO(n_295), .S(n_296), .A(n_272), .B(n_261), .CI(n_245));
  ADDFX1 g4551(.CO(n_293), .S(n_294), .A(n_187), .B(n_251), .CI(n_252));
  NOR2XL g4552(.Y(n_292), .A(n_102), .B(n_287));
  ADDFX1 g4553(.CO(n_290), .S(out_0[2]), .A(n_231), .B(n_246), .CI(n_257));
  ADDFX1 g4554(.CO(n_288), .S(n_289), .A(n_221), .B(n_270), .CI(n_236));
  ADDFX1 g4555(.CO(n_287), .S(n_286), .A(n_103), .B(n_130), .CI(n_266));
  ADDFX1 g4556(.CO(n_284), .S(n_285), .A(n_239), .B(n_244), .CI(n_237));
  ADDFX1 g4557(.CO(n_282), .S(n_283), .A(n_186), .B(n_197), .CI(n_250));
  ADDFX1 g4558(.CO(n_280), .S(n_281), .A(n_195), .B(n_238), .CI(n_205));
  ADDFX1 g4559(.CO(n_278), .S(n_279), .A(n_230), .B(n_217), .CI(n_256));
  ADDFX1 g4560(.CO(n_276), .S(n_277), .A(n_234), .B(n_112), .CI(n_243));
  ADDFX1 g4561(.CO(n_274), .S(n_275), .A(n_164), .B(n_228), .CI(n_233));
  ADDFX1 g4562(.CO(n_272), .S(n_273), .A(n_151), .B(n_223), .CI(n_209));
  ADDFX1 g4563(.CO(n_270), .S(n_271), .A(n_183), .B(n_224), .CI(n_181));
  ADDFX1 g4564(.CO(n_268), .S(n_269), .A(n_232), .B(n_235), .CI(n_113));
  ADDFX1 g4565(.CO(n_266), .S(n_267), .A(n_218), .B(n_131), .CI(n_242));
  ADDFX1 g4566(.CO(n_264), .S(n_265), .A(n_208), .B(n_225), .CI(n_240));
  ADDFX1 g4567(.CO(n_262), .S(n_263), .A(n_216), .B(n_207), .CI(n_227));
  ADDFX1 g4568(.CO(n_260), .S(n_261), .A(n_215), .B(n_150), .CI(n_213));
  ADDFX1 g4569(.CO(n_258), .S(n_259), .A(n_184), .B(n_202), .CI(n_189));
  ADDFX1 g4570(.CO(n_256), .S(n_257), .A(n_198), .B(n_175), .CI(n_193));
  ADDFX1 g4571(.CO(n_254), .S(n_255), .A(n_204), .B(n_220), .CI(n_211));
  ADDFX1 g4572(.CO(n_252), .S(n_253), .A(n_194), .B(n_108), .CI(n_165));
  ADDFX1 g4573(.CO(n_250), .S(n_251), .A(n_210), .B(n_119), .CI(n_123));
  ADDFX1 g4574(.CO(n_248), .S(n_249), .A(n_192), .B(n_185), .CI(n_203));
  ADDFX1 g4575(.CO(n_246), .S(out_0[1]), .A(n_162), .B(n_179), .CI(n_199));
  ADDFX1 g4576(.CO(n_244), .S(n_245), .A(n_133), .B(n_222), .CI(n_115));
  ADDFX1 g4577(.CO(n_242), .S(n_243), .A(n_219), .B(n_86), .CI(n_22));
  ADDFX1 g4578(.CO(n_240), .S(n_241), .A(n_188), .B(n_206), .CI(n_173));
  ADDFX1 g4579(.CO(n_238), .S(n_239), .A(n_135), .B(n_214), .CI(n_141));
  ADDFX1 g4580(.CO(n_236), .S(n_237), .A(n_125), .B(n_212), .CI(n_147));
  ADDFX1 g4581(.CO(n_234), .S(n_235), .A(n_170), .B(in_3[11]), .CI(n_191));
  ADDFX1 g4582(.CO(n_232), .S(n_233), .A(n_176), .B(n_171), .CI(in_18[10]));
  ADDFX1 g4583(.CO(n_230), .S(n_231), .A(n_121), .B(n_178), .CI(n_139));
  ADDFX1 g4584(.CO(n_228), .S(n_229), .A(n_81), .B(n_177), .CI(n_153));
  ADDFX1 g4585(.CO(n_226), .S(n_227), .A(n_166), .B(n_129), .CI(n_157));
  ADDFX1 g4586(.CO(n_224), .S(n_225), .A(n_63), .B(n_41), .CI(n_172));
  ADDFX1 g4587(.CO(n_222), .S(n_223), .A(n_154), .B(n_143), .CI(n_156));
  ADDFX1 g4588(.CO(n_220), .S(n_221), .A(n_145), .B(n_182), .CI(n_146));
  ADDFX1 g4589(.CO(n_218), .S(n_219), .A(in_17[12]), .B(in_13[12]), .CI(n_190));
  ADDFX1 g4590(.CO(n_216), .S(n_217), .A(n_174), .B(n_167), .CI(n_159));
  ADDFX1 g4591(.CO(n_214), .S(n_215), .A(n_33), .B(n_142), .CI(n_28));
  ADDFX1 g4592(.CO(n_212), .S(n_213), .A(n_107), .B(n_136), .CI(n_160));
  ADDFX1 g4593(.CO(n_210), .S(n_211), .A(n_126), .B(n_144), .CI(in_3[9]));
  ADDFX1 g4594(.CO(n_208), .S(n_209), .A(n_128), .B(n_161), .CI(n_137));
  ADDFX1 g4595(.CO(n_206), .S(n_207), .A(n_158), .B(n_45), .CI(n_155));
  ADDFX1 g4596(.CO(n_204), .S(n_205), .A(n_140), .B(n_124), .CI(n_127));
  ADDFX1 g4597(.CO(n_202), .S(n_203), .A(n_138), .B(n_31), .CI(n_149));
  ADDFX1 g4598(.CO(n_200), .S(n_201), .A(n_111), .B(n_180), .CI(n_109));
  ADDFX1 g4599(.CO(n_198), .S(n_199), .A(n_76), .B(n_101), .CI(n_169));
  ADDFX1 g4600(.CO(n_196), .S(n_197), .A(n_87), .B(n_118), .CI(n_122));
  ADDFX1 g4601(.CO(n_194), .S(n_195), .A(n_16), .B(n_105), .CI(n_134));
  ADDFX1 g4602(.CO(n_192), .S(n_193), .A(n_168), .B(n_75), .CI(n_91));
  ADDFX1 g4603(.CO(n_190), .S(n_191), .A(n_11), .B(n_5), .CI(n_116));
  ADDFX1 g4604(.CO(n_188), .S(n_189), .A(n_73), .B(n_65), .CI(n_148));
  ADDFX1 g4605(.CO(n_186), .S(n_187), .A(n_97), .B(n_80), .CI(n_152));
  ADDFX1 g4606(.CO(n_184), .S(n_185), .A(n_120), .B(n_90), .CI(n_57));
  ADDFX1 g4607(.CO(n_182), .S(n_183), .A(n_132), .B(n_62), .CI(n_40));
  ADDFX1 g4608(.CO(n_180), .S(n_181), .A(n_59), .B(n_55), .CI(n_114));
  ADDFX1 g4609(.CO(n_178), .S(n_179), .A(n_67), .B(n_83), .CI(n_39));
  ADDFX1 g4610(.CO(n_176), .S(n_177), .A(n_98), .B(in_13[9]), .CI(n_23));
  ADDFX1 g4611(.CO(n_174), .S(n_175), .A(n_35), .B(n_100), .CI(n_85));
  ADDFX1 g4612(.CO(n_172), .S(n_173), .A(n_64), .B(n_72), .CI(in_18[5]));
  ADDHX1 g4613(.CO(n_170), .S(n_171), .A(in_17[10]), .B(n_117));
  ADDFX1 g4614(.CO(n_168), .S(n_169), .A(n_92), .B(n_48), .CI(n_69));
  ADDFX1 g4615(.CO(n_166), .S(n_167), .A(n_43), .B(n_37), .CI(n_47));
  ADDFX1 g4616(.CO(n_164), .S(n_165), .A(n_61), .B(n_110), .CI(in_18[9]));
  ADDFX1 g4617(.CO(n_162), .S(out_0[0]), .A(n_49), .B(n_93), .CI(n_77));
  ADDFX1 g4618(.CO(n_160), .S(n_161), .A(n_17), .B(n_79), .CI(in_3[5]));
  ADDFX1 g4619(.CO(n_158), .S(n_159), .A(n_34), .B(n_84), .CI(n_74));
  ADDFX1 g4620(.CO(n_156), .S(n_157), .A(n_36), .B(n_46), .CI(in_3[4]));
  ADDFX1 g4621(.CO(n_154), .S(n_155), .A(n_42), .B(n_95), .CI(in_18[4]));
  ADDFX1 g4622(.CO(n_152), .S(n_153), .A(in_9[9]), .B(n_104), .CI(in_8[9]));
  ADDFX1 g4623(.CO(n_150), .S(n_151), .A(n_71), .B(n_44), .CI(n_29));
  ADDFX1 g4624(.CO(n_148), .S(n_149), .A(n_88), .B(in_3[3]), .CI(in_18[3]));
  ADDFX1 g4625(.CO(n_146), .S(n_147), .A(n_106), .B(in_3[7]), .CI(in_18[7]));
  ADDFX1 g4626(.CO(n_144), .S(n_145), .A(n_99), .B(in_14[8]), .CI(in_13[8]));
  ADDFX1 g4627(.CO(n_142), .S(n_143), .A(n_94), .B(in_9[5]), .CI(in_19[5]));
  ADDFX1 g4628(.CO(n_140), .S(n_141), .A(n_32), .B(in_13[7]), .CI(in_16[7]));
  ADDFX1 g4629(.CO(n_138), .S(n_139), .A(n_68), .B(n_89), .CI(n_38));
  ADDFX1 g4630(.CO(n_136), .S(n_137), .A(n_26), .B(in_13[5]), .CI(in_8[5]));
  ADDFX1 g4631(.CO(n_134), .S(n_135), .A(n_18), .B(n_52), .CI(in_14[7]));
  ADDFX1 g4632(.CO(n_132), .S(n_133), .A(n_53), .B(n_78), .CI(in_11[6]));
  ADDFX1 g4633(.CO(n_130), .S(n_131), .A(n_4), .B(n_25), .CI(n_1));
  ADDFX1 g4634(.CO(n_128), .S(n_129), .A(n_27), .B(n_56), .CI(n_30));
  ADDFX1 g4635(.CO(n_126), .S(n_127), .A(n_50), .B(in_9[8]), .CI(in_11[8]));
  ADDFX1 g4636(.CO(n_124), .S(n_125), .A(n_51), .B(in_6[7]), .CI(in_8[7]));
  ADDFX1 g4637(.CO(n_122), .S(n_123), .A(n_60), .B(in_8[10]), .CI(in_3[10]));
  ADDFX1 g4638(.CO(n_120), .S(n_121), .A(n_82), .B(n_66), .CI(in_19[2]));
  ADDFX1 g4639(.CO(n_118), .S(n_119), .A(in_11[10]), .B(n_24), .CI(in_13[10]));
  ADDFX1 g4640(.CO(n_116), .S(n_117), .A(in_2[10]), .B(n_14), .CI(n_7));
  ADDFX1 g4641(.CO(n_114), .S(n_115), .A(n_70), .B(in_3[6]), .CI(in_18[6]));
  ADDFX1 g4642(.CO(n_112), .S(n_113), .A(n_96), .B(in_13[11]), .CI(in_8[11]));
  ADDFX1 g4643(.CO(n_110), .S(n_111), .A(n_58), .B(in_6[8]), .CI(in_8[8]));
  ADDFX1 g4644(.CO(n_108), .S(n_109), .A(n_54), .B(in_3[8]), .CI(in_18[8]));
  ADDFX1 g4645(.CO(n_106), .S(n_107), .A(n_9), .B(in_19[6]), .CI(in_12[6]));
  ADDFX1 g4646(.CO(n_104), .S(n_105), .A(n_13), .B(in_10[8]), .CI(in_16[8]));
  OAI2BB1X1 g4647(.Y(n_103), .A0N(n_8), .A1N(n_21), .B0(n_102));
  OR2X1 g4648(.Y(n_102), .A(n_8), .B(n_21));
  ADDFX1 g4649(.CO(n_100), .S(n_101), .A(n_19), .B(in_19[1]), .CI(in_3[1]));
  ADDFX1 g4650(.CO(n_98), .S(n_99), .A(in_2[8]), .B(in_15[8]), .CI(in_19[8]));
  ADDFX1 g4651(.CO(n_96), .S(n_97), .A(in_10[10]), .B(in_6[10]), .CI(in_9[10]));
  ADDFX1 g4652(.CO(n_94), .S(n_95), .A(in_2[4]), .B(in_5[4]), .CI(in_15[4]));
  ADDFX1 g4653(.CO(n_92), .S(n_93), .A(in_3[0]), .B(in_18[0]), .CI(in_5[0]));
  ADDFX1 g4654(.CO(n_90), .S(n_91), .A(in_8[2]), .B(in_3[2]), .CI(in_18[2]));
  ADDFX1 g4655(.CO(n_88), .S(n_89), .A(n_2), .B(in_10[2]), .CI(in_15[2]));
  ADDFX1 g4656(.CO(n_86), .S(n_87), .A(in_17[11]), .B(in_11[11]), .CI(in_18[11]));
  ADDFX1 g4657(.CO(n_84), .S(n_85), .A(in_9[2]), .B(in_11[2]), .CI(in_14[2]));
  ADDFX1 g4658(.CO(n_82), .S(n_83), .A(in_0[1]), .B(in_9[1]), .CI(in_5[1]));
  ADDFX1 g4659(.CO(n_80), .S(n_81), .A(n_12), .B(in_6[9]), .CI(in_11[9]));
  ADDFX1 g4660(.CO(n_78), .S(n_79), .A(in_0[5]), .B(in_15[5]), .CI(in_17[5]));
  ADDFX1 g4661(.CO(n_76), .S(n_77), .A(in_0[0]), .B(in_8[0]), .CI(n_20));
  ADDFX1 g4662(.CO(n_74), .S(n_75), .A(in_12[2]), .B(in_16[2]), .CI(in_6[2]));
  ADDFX1 g4663(.CO(n_72), .S(n_73), .A(in_11[4]), .B(in_14[4]), .CI(in_6[4]));
  ADDFX1 g4664(.CO(n_70), .S(n_71), .A(in_10[5]), .B(in_12[5]), .CI(in_14[5]));
  ADDFX1 g4665(.CO(n_68), .S(n_69), .A(in_11[1]), .B(in_13[1]), .CI(in_14[1]));
  ADDFX1 g4666(.CO(n_66), .S(n_67), .A(in_12[1]), .B(in_8[1]), .CI(in_15[1]));
  ADDFX1 g4667(.CO(n_64), .S(n_65), .A(in_9[4]), .B(in_12[4]), .CI(in_19[4]));
  ADDFX1 g4668(.CO(n_62), .S(n_63), .A(in_6[6]), .B(in_13[6]), .CI(in_16[6]));
  ADDFX1 g4669(.CO(n_60), .S(n_61), .A(in_2[9]), .B(in_17[9]), .CI(in_10[9]));
  ADDFX1 g4670(.CO(n_58), .S(n_59), .A(in_17[7]), .B(in_10[7]), .CI(in_12[7]));
  ADDFX1 g4671(.CO(n_56), .S(n_57), .A(in_11[3]), .B(in_16[3]), .CI(in_19[3]));
  ADDFX1 g4672(.CO(n_54), .S(n_55), .A(in_19[7]), .B(in_9[7]), .CI(in_11[7]));
  ADDFX1 g4673(.CO(n_52), .S(n_53), .A(in_0[6]), .B(in_2[6]), .CI(in_15[6]));
  ADDFX1 g4674(.CO(n_50), .S(n_51), .A(in_5[6]), .B(in_0[7]), .CI(in_15[7]));
  ADDFX1 g4675(.CO(n_48), .S(n_49), .A(in_9[0]), .B(in_11[0]), .CI(in_19[0]));
  ADDFX1 g4676(.CO(n_46), .S(n_47), .A(in_13[3]), .B(in_12[3]), .CI(in_14[3]));
  ADDFX1 g4677(.CO(n_44), .S(n_45), .A(in_13[4]), .B(in_8[4]), .CI(in_16[4]));
  ADDFX1 g4678(.CO(n_42), .S(n_43), .A(in_2[3]), .B(in_5[3]), .CI(in_17[3]));
  ADDFX1 g4679(.CO(n_40), .S(n_41), .A(in_14[6]), .B(in_9[6]), .CI(in_8[6]));
  ADDFX1 g4680(.CO(n_38), .S(n_39), .A(in_16[1]), .B(in_18[1]), .CI(in_6[1]));
  ADDFX1 g4681(.CO(n_36), .S(n_37), .A(in_0[3]), .B(in_15[3]), .CI(in_10[3]));
  ADDFX1 g4682(.CO(n_34), .S(n_35), .A(in_5[2]), .B(in_0[2]), .CI(in_13[2]));
  ADDFX1 g4683(.CO(n_32), .S(n_33), .A(n_6), .B(in_10[6]), .CI(in_17[6]));
  ADDFX1 g4684(.CO(n_30), .S(n_31), .A(in_9[3]), .B(in_6[3]), .CI(in_8[3]));
  ADDFX1 g4685(.CO(n_28), .S(n_29), .A(in_11[5]), .B(in_6[5]), .CI(in_16[5]));
  ADDFX1 g4686(.CO(n_26), .S(n_27), .A(in_0[4]), .B(in_17[4]), .CI(in_10[4]));
  OAI21X1 g4687(.Y(n_25), .A0(n_11), .A1(n_10), .B0(n_8));
  AO22XL g4688(.Y(n_24), .A0(n_11), .A1(n_15), .B0(in_12[9]), .B1(in_14[9]));
  XOR2XL g4689(.Y(n_23), .A(n_14), .B(n_15));
  XNOR2X1 g4691(.Y(n_22), .A(n_11), .B(n_0));
  NOR2XL g4692(.Y(n_21), .A(in_17[12]), .B(n_0));
  ADDHX1 g4694(.CO(n_19), .S(n_20), .A(in_6[0]), .B(in_16[0]));
  OAI2BB1X1 g4695(.Y(n_18), .A0N(in_5[7]), .A1N(in_2[7]), .B0(n_13));
  OAI2BB1X1 g4696(.Y(n_17), .A0N(in_5[5]), .A1N(in_2[5]), .B0(n_9));
  OAI2BB1X1 g4697(.Y(n_16), .A0N(in_17[8]), .A1N(in_12[8]), .B0(n_12));
  XNOR2X1 g4699(.Y(n_15), .A(in_19[8]), .B(in_16[8]));
  XOR2XL g4700(.Y(n_14), .A(in_12[9]), .B(in_14[9]));
  OR2X1 g4701(.Y(n_13), .A(in_5[7]), .B(in_2[7]));
  OR2X1 g4702(.Y(n_12), .A(in_17[8]), .B(in_12[8]));
  OR2X1 g4703(.Y(n_11), .A(in_12[9]), .B(in_14[9]));
  NOR2X1 g4704(.Y(n_10), .A(in_8[12]), .B(in_18[11]));
  OR2X1 g4705(.Y(n_9), .A(in_5[5]), .B(in_2[5]));
  NAND2X1 g4706(.Y(n_8), .A(in_8[12]), .B(in_18[11]));
  NAND2XL g4707(.Y(n_7), .A(in_19[8]), .B(in_16[8]));
  INVX1 g4708(.Y(n_6), .A(in_5[6]));
  INVX1 g4709(.Y(n_5), .A(in_10[11]));
  INVX1 g4711(.Y(n_4), .A(in_13[12]));
  BUFX2 drc_bufs(.Y(n_2), .A(in_2[2]));
  XOR2XL g2(.Y(n_1), .A(in_17[12]), .B(n_0));
  CLKXOR2X1 g4712(.Y(n_0), .A(in_18[11]), .B(in_8[12]));
endmodule

module csa_tree_ADD_TC_OP_19_group_2425(in_0, in_1, in_2, in_3, in_4, in_5, in_6
    , in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, 
    in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_445, n_443, n_441, n_439, n_437, n_435, n_433, n_431, n_429, n_427, 
    n_426, n_425, n_424, n_423, n_421, n_420, n_419, n_418, n_417, n_416, 
    n_415, n_414, n_413, n_412, n_411, n_409, n_408, n_407, n_406, n_405, 
    n_404, n_403, n_402, n_401, n_400, n_399, n_398, n_397, n_396, n_395, 
    n_394, n_393, n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, 
    n_383, n_382, n_381, n_380, n_379, n_378, n_377, n_376, n_375, n_374, 
    n_373, n_372, n_371, n_370, n_369, n_368, n_367, n_365, n_364, n_363, 
    n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, 
    n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, 
    n_342, n_341, n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, 
    n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, 
    n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, n_312, 
    n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, 
    n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, 
    n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, n_282, 
    n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, 
    n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, 
    n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, n_252, 
    n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_243, n_242, n_241, 
    n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, 
    n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, 
    n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, 
    n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, 
    n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, 
    n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, 
    n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, 
    n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, 
    n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, 
    n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, 
    n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
    n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
    n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, 
    n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
    n_3, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  AOI21X2 g6018(.Y(out_0[18]), .A0(n_131), .A1(n_285), .B0(n_445));
  ADDFX1 g6019(.CO(n_445), .S(out_0[15]), .A(n_310), .B(n_389), .CI(n_443));
  ADDFX1 g6020(.CO(n_443), .S(out_0[14]), .A(n_390), .B(n_417), .CI(n_441));
  ADDFX1 g6021(.CO(n_441), .S(out_0[13]), .A(n_423), .B(n_418), .CI(n_439));
  ADDFX1 g6022(.CO(n_439), .S(out_0[12]), .A(n_425), .B(n_424), .CI(n_437));
  ADDFX1 g6023(.CO(n_437), .S(out_0[11]), .A(n_419), .B(n_426), .CI(n_435));
  ADDFX1 g6024(.CO(n_435), .S(out_0[10]), .A(n_411), .B(n_420), .CI(n_433));
  ADDFX1 g6025(.CO(n_433), .S(out_0[9]), .A(n_415), .B(n_412), .CI(n_431));
  ADDFX1 g6026(.CO(n_431), .S(out_0[8]), .A(n_413), .B(n_416), .CI(n_429));
  ADDFX1 g6027(.CO(n_429), .S(out_0[7]), .A(n_407), .B(n_414), .CI(n_427));
  ADDFX1 g6028(.CO(n_427), .S(out_0[6]), .A(n_399), .B(n_421), .CI(n_408));
  ADDFX1 g6029(.CO(n_425), .S(n_426), .A(n_384), .B(n_406), .CI(n_403));
  ADDFX1 g6030(.CO(n_423), .S(n_424), .A(n_383), .B(n_405), .CI(n_402));
  ADDFX1 g6031(.CO(n_421), .S(out_0[5]), .A(n_379), .B(n_400), .CI(n_409));
  ADDFX1 g6032(.CO(n_419), .S(n_420), .A(n_382), .B(n_397), .CI(n_404));
  ADDFX1 g6033(.CO(n_417), .S(n_418), .A(n_385), .B(n_401), .CI(n_372));
  ADDFX1 g6034(.CO(n_415), .S(n_416), .A(n_387), .B(n_370), .CI(n_396));
  ADDFX1 g6035(.CO(n_413), .S(n_414), .A(n_393), .B(n_368), .CI(n_388));
  ADDFX1 g6036(.CO(n_411), .S(n_412), .A(n_374), .B(n_395), .CI(n_398));
  ADDFX1 g6037(.CO(n_409), .S(out_0[4]), .A(n_355), .B(n_380), .CI(n_391));
  ADDFX1 g6038(.CO(n_407), .S(n_408), .A(n_375), .B(n_394), .CI(n_362));
  ADDFX1 g6039(.CO(n_405), .S(n_406), .A(n_364), .B(n_377), .CI(n_381));
  ADDFX1 g6040(.CO(n_403), .S(n_404), .A(n_351), .B(n_373), .CI(n_378));
  ADDFX1 g6041(.CO(n_401), .S(n_402), .A(n_363), .B(n_346), .CI(n_386));
  ADDFX1 g6042(.CO(n_399), .S(n_400), .A(n_357), .B(n_360), .CI(n_376));
  ADDFX1 g6043(.CO(n_397), .S(n_398), .A(n_348), .B(n_369), .CI(n_352));
  ADDFX1 g6044(.CO(n_395), .S(n_396), .A(n_324), .B(n_367), .CI(n_354));
  ADDFX1 g6045(.CO(n_393), .S(n_394), .A(n_316), .B(n_359), .CI(n_338));
  ADDFX1 g6046(.CO(n_391), .S(out_0[3]), .A(n_365), .B(n_334), .CI(n_356));
  ADDFX1 g6047(.CO(n_389), .S(n_390), .A(n_272), .B(n_329), .CI(n_371));
  ADDFX1 g6048(.CO(n_387), .S(n_388), .A(n_314), .B(n_340), .CI(n_361));
  ADDFX1 g6049(.CO(n_385), .S(n_386), .A(n_343), .B(n_276), .CI(n_349));
  ADDFX1 g6050(.CO(n_383), .S(n_384), .A(n_344), .B(n_341), .CI(n_350));
  ADDFX1 g6051(.CO(n_381), .S(n_382), .A(n_347), .B(n_303), .CI(n_342));
  ADDFX1 g6052(.CO(n_379), .S(n_380), .A(n_333), .B(n_336), .CI(n_358));
  ADDFX1 g6053(.CO(n_377), .S(n_378), .A(n_273), .B(n_320), .CI(n_317));
  ADDFX1 g6054(.CO(n_375), .S(n_376), .A(n_335), .B(n_309), .CI(n_332));
  ADDFX1 g6055(.CO(n_373), .S(n_374), .A(n_323), .B(n_318), .CI(n_353));
  ADDFX1 g6056(.CO(n_371), .S(n_372), .A(n_275), .B(n_345), .CI(n_330));
  ADDFX1 g6057(.CO(n_369), .S(n_370), .A(n_313), .B(n_339), .CI(n_328));
  ADDFX1 g6058(.CO(n_367), .S(n_368), .A(n_315), .B(n_337), .CI(n_293));
  ADDFX1 g6059(.CO(n_365), .S(out_0[2]), .A(n_280), .B(n_321), .CI(n_326));
  ADDFX1 g6060(.CO(n_363), .S(n_364), .A(n_263), .B(n_319), .CI(n_302));
  ADDFX1 g6061(.CO(n_361), .S(n_362), .A(n_308), .B(n_331), .CI(n_287));
  ADDFX1 g6062(.CO(n_359), .S(n_360), .A(n_301), .B(n_311), .CI(n_232));
  ADDFX1 g6063(.CO(n_357), .S(n_358), .A(n_298), .B(n_307), .CI(n_312));
  ADDFX1 g6064(.CO(n_355), .S(n_356), .A(n_325), .B(n_282), .CI(n_299));
  ADDFX1 g6065(.CO(n_353), .S(n_354), .A(n_238), .B(n_292), .CI(n_305));
  ADDFX1 g6066(.CO(n_351), .S(n_352), .A(n_289), .B(n_274), .CI(n_327));
  ADDFX1 g6067(.CO(n_349), .S(n_350), .A(n_221), .B(n_225), .CI(n_284));
  ADDFX1 g6068(.CO(n_347), .S(n_348), .A(n_237), .B(n_297), .CI(n_304));
  ADDFX1 g6069(.CO(n_345), .S(n_346), .A(n_283), .B(n_265), .CI(n_262));
  ADDFX1 g6070(.CO(n_343), .S(n_344), .A(n_290), .B(n_187), .CI(n_194));
  ADDFX1 g6071(.CO(n_341), .S(n_342), .A(n_291), .B(n_288), .CI(n_226));
  ADDFX1 g6072(.CO(n_339), .S(n_340), .A(n_295), .B(n_286), .CI(n_254));
  ADDFX1 g6073(.CO(n_337), .S(n_338), .A(n_300), .B(n_278), .CI(n_242));
  ADDFX1 g6074(.CO(n_335), .S(n_336), .A(n_281), .B(n_258), .CI(n_240));
  ADDFX1 g6075(.CO(n_333), .S(n_334), .A(n_266), .B(n_279), .CI(n_271));
  ADDFX1 g6076(.CO(n_331), .S(n_332), .A(n_239), .B(n_306), .CI(n_250));
  ADDFX1 g6077(.CO(n_329), .S(n_330), .A(n_202), .B(n_264), .CI(n_251));
  ADDFX1 g6078(.CO(n_327), .S(n_328), .A(n_247), .B(n_294), .CI(n_181));
  ADDFX1 g6079(.CO(n_325), .S(n_326), .A(n_268), .B(n_197), .CI(n_267));
  ADDFX1 g6080(.CO(n_323), .S(n_324), .A(n_224), .B(n_253), .CI(n_260));
  ADDFX1 g6081(.CO(n_321), .S(out_0[1]), .A(n_243), .B(n_269), .CI(n_189));
  ADDFX1 g6082(.CO(n_319), .S(n_320), .A(n_235), .B(n_296), .CI(n_85));
  ADDFX1 g6083(.CO(n_317), .S(n_318), .A(n_236), .B(n_259), .CI(n_219));
  ADDFX1 g6084(.CO(n_315), .S(n_316), .A(n_246), .B(n_230), .CI(n_231));
  ADDFX1 g6085(.CO(n_313), .S(n_314), .A(n_248), .B(n_241), .CI(n_277));
  ADDFX1 g6086(.CO(n_311), .S(n_312), .A(n_217), .B(n_215), .CI(n_270));
  XOR2XL g6087(.Y(n_310), .A(n_131), .B(n_285));
  ADDFX1 g6088(.CO(n_308), .S(n_309), .A(n_173), .B(n_183), .CI(n_257));
  ADDFX1 g6089(.CO(n_306), .S(n_307), .A(n_213), .B(n_204), .CI(n_255));
  ADDFX1 g6090(.CO(n_304), .S(n_305), .A(n_160), .B(n_234), .CI(n_167));
  ADDFX1 g6091(.CO(n_302), .S(n_303), .A(n_222), .B(n_218), .CI(n_195));
  ADDFX1 g6092(.CO(n_300), .S(n_301), .A(n_216), .B(n_179), .CI(n_214));
  ADDFX1 g6093(.CO(n_298), .S(n_299), .A(n_196), .B(n_205), .CI(n_256));
  ADDFX1 g6094(.CO(n_296), .S(n_297), .A(n_52), .B(n_233), .CI(n_166));
  ADDFX1 g6095(.CO(n_294), .S(n_295), .A(n_245), .B(n_190), .CI(n_135));
  ADDFX1 g6096(.CO(n_292), .S(n_293), .A(n_229), .B(n_161), .CI(n_207));
  ADDFX1 g6097(.CO(n_290), .S(n_291), .A(n_227), .B(n_177), .CI(n_184));
  ADDFX1 g6098(.CO(n_288), .S(n_289), .A(n_228), .B(n_121), .CI(n_180));
  ADDFX1 g6099(.CO(n_286), .S(n_287), .A(n_172), .B(n_249), .CI(n_191));
  ADDFX1 g6100(.CO(n_283), .S(n_284), .A(n_176), .B(n_132), .CI(in_8[11]));
  ADDFX1 g6101(.CO(n_281), .S(n_282), .A(n_175), .B(n_171), .CI(n_210));
  ADDFX1 g6102(.CO(n_279), .S(n_280), .A(n_201), .B(n_188), .CI(n_211));
  ADDFX1 g6103(.CO(n_277), .S(n_278), .A(n_178), .B(n_182), .CI(n_95));
  ADDFX1 g6104(.CO(n_275), .S(n_276), .A(n_203), .B(n_148), .CI(n_186));
  ADDFX1 g6105(.CO(n_273), .S(n_274), .A(n_185), .B(n_223), .CI(n_45));
  OAI2BB1X1 g6106(.Y(n_285), .A0N(n_130), .A1N(n_209), .B0(n_261));
  CLKXOR2X1 g6107(.Y(n_272), .A(n_220), .B(n_252));
  ADDFX1 g6108(.CO(n_270), .S(n_271), .A(n_200), .B(n_87), .CI(n_147));
  ADDFX1 g6109(.CO(n_268), .S(n_269), .A(n_156), .B(n_165), .CI(n_193));
  ADDFX1 g6110(.CO(n_266), .S(n_267), .A(n_164), .B(n_169), .CI(n_192));
  ADDFX1 g6111(.CO(n_264), .S(n_265), .A(in_13[12]), .B(n_198), .CI(n_159));
  ADDFX1 g6112(.CO(n_262), .S(n_263), .A(n_199), .B(n_84), .CI(n_149));
  OAI21X1 g6113(.Y(n_261), .A0(n_130), .A1(n_209), .B0(n_252));
  ADDFX1 g6114(.CO(n_259), .S(n_260), .A(n_104), .B(n_152), .CI(n_206));
  ADDFX1 g6115(.CO(n_257), .S(n_258), .A(n_174), .B(n_25), .CI(n_139));
  ADDFX1 g6116(.CO(n_255), .S(n_256), .A(n_168), .B(n_65), .CI(n_115));
  ADDFX1 g6117(.CO(n_253), .S(n_254), .A(n_105), .B(n_153), .CI(n_123));
  ADDFX1 g6118(.CO(n_252), .S(n_251), .A(n_5), .B(n_158), .CI(n_208));
  ADDFX1 g6119(.CO(n_249), .S(n_250), .A(n_212), .B(n_138), .CI(n_59));
  ADDFX1 g6120(.CO(n_247), .S(n_248), .A(n_154), .B(n_141), .CI(n_94));
  ADDFX1 g6121(.CO(n_245), .S(n_246), .A(n_151), .B(n_56), .CI(n_58));
  ADDFX1 g6122(.CO(n_243), .S(out_0[0]), .A(n_127), .B(n_63), .CI(n_157));
  ADDFX1 g6123(.CO(n_241), .S(n_242), .A(n_79), .B(n_155), .CI(n_31));
  ADDFX1 g6124(.CO(n_239), .S(n_240), .A(n_170), .B(n_97), .CI(n_33));
  ADDFX1 g6125(.CO(n_237), .S(n_238), .A(n_134), .B(n_67), .CI(n_53));
  ADDFX1 g6126(.CO(n_235), .S(n_236), .A(n_144), .B(n_137), .CI(n_66));
  ADDFX1 g6127(.CO(n_233), .S(n_234), .A(n_48), .B(n_143), .CI(in_8[8]));
  ADDFX1 g6128(.CO(n_231), .S(n_232), .A(n_57), .B(n_47), .CI(n_163));
  ADDFX1 g6129(.CO(n_229), .S(n_230), .A(n_27), .B(n_162), .CI(n_46));
  ADDFX1 g6130(.CO(n_227), .S(n_228), .A(in_14[9]), .B(n_142), .CI(in_9[9]));
  ADDFX1 g6131(.CO(n_225), .S(n_226), .A(n_89), .B(n_120), .CI(n_133));
  ADDFX1 g6132(.CO(n_223), .S(n_224), .A(n_145), .B(n_125), .CI(n_122));
  ADDFX1 g6133(.CO(n_221), .S(n_222), .A(n_136), .B(n_50), .CI(n_44));
  NOR2X1 g6134(.Y(n_220), .A(n_131), .B(n_209));
  ADDFX1 g6135(.CO(n_218), .S(n_219), .A(n_124), .B(n_51), .CI(in_6[9]));
  ADDFX1 g6136(.CO(n_216), .S(n_217), .A(n_64), .B(n_114), .CI(n_113));
  ADDFX1 g6137(.CO(n_214), .S(n_215), .A(n_86), .B(n_99), .CI(n_146));
  ADDFX1 g6138(.CO(n_212), .S(n_213), .A(n_35), .B(n_92), .CI(n_38));
  ADDFX1 g6139(.CO(n_210), .S(n_211), .A(n_110), .B(n_83), .CI(n_55));
  ADDFX1 g6140(.CO(n_209), .S(n_208), .A(n_128), .B(in_6[11]), .CI(n_0));
  ADDFX1 g6141(.CO(n_206), .S(n_207), .A(n_150), .B(n_26), .CI(in_6[7]));
  ADDFX1 g6142(.CO(n_204), .S(n_205), .A(n_39), .B(n_93), .CI(n_118));
  ADDFX1 g6143(.CO(n_202), .S(n_203), .A(n_10), .B(in_17[12]), .CI(n_129));
  ADDFX1 g6144(.CO(n_200), .S(n_201), .A(n_69), .B(n_41), .CI(n_100));
  ADDFX1 g6145(.CO(n_198), .S(n_199), .A(n_20), .B(n_23), .CI(in_17[11]));
  ADDFX1 g6146(.CO(n_196), .S(n_197), .A(n_29), .B(n_77), .CI(n_119));
  ADDFX1 g6147(.CO(n_194), .S(n_195), .A(n_117), .B(in_5[10]), .CI(in_6[10]));
  ADDFX1 g6148(.CO(n_192), .S(n_193), .A(n_108), .B(n_103), .CI(n_61));
  ADDFX1 g6149(.CO(n_190), .S(n_191), .A(n_36), .B(n_72), .CI(in_6[6]));
  ADDFX1 g6150(.CO(n_188), .S(n_189), .A(n_75), .B(n_101), .CI(n_111));
  ADDFX1 g6151(.CO(n_186), .S(n_187), .A(n_116), .B(n_88), .CI(in_13[11]));
  ADDFX1 g6152(.CO(n_184), .S(n_185), .A(n_107), .B(in_16[9]), .CI(in_4[9]));
  ADDFX1 g6153(.CO(n_182), .S(n_183), .A(n_34), .B(n_98), .CI(in_6[5]));
  ADDFX1 g6154(.CO(n_180), .S(n_181), .A(in_4[8]), .B(n_140), .CI(in_6[8]));
  ADDFX1 g6155(.CO(n_178), .S(n_179), .A(n_112), .B(n_96), .CI(n_37));
  ADDFX1 g6156(.CO(n_176), .S(n_177), .A(n_106), .B(in_14[10]), .CI(in_3[10]));
  ADDFX1 g6157(.CO(n_174), .S(n_175), .A(n_28), .B(n_76), .CI(n_82));
  ADDFX1 g6158(.CO(n_172), .S(n_173), .A(n_24), .B(n_73), .CI(n_32));
  ADDFX1 g6159(.CO(n_170), .S(n_171), .A(n_40), .B(n_81), .CI(n_54));
  ADDFX1 g6160(.CO(n_168), .S(n_169), .A(n_102), .B(n_60), .CI(n_74));
  ADDFX1 g6161(.CO(n_166), .S(n_167), .A(n_42), .B(in_19[8]), .CI(in_13[8]));
  ADDFX1 g6162(.CO(n_164), .S(n_165), .A(n_19), .B(n_126), .CI(n_62));
  ADDFX1 g6163(.CO(n_162), .S(n_163), .A(n_71), .B(in_4[5]), .CI(in_3[5]));
  ADDFX1 g6164(.CO(n_160), .S(n_161), .A(n_43), .B(n_78), .CI(n_30));
  ADDFX1 g6165(.CO(n_158), .S(n_159), .A(n_22), .B(in_8[12]), .CI(n_3));
  ADDFX1 g6166(.CO(n_156), .S(n_157), .A(in_13[0]), .B(in_16[0]), .CI(n_109));
  ADDFX1 g6167(.CO(n_154), .S(n_155), .A(n_91), .B(in_19[6]), .CI(in_2[6]));
  ADDFX1 g6168(.CO(n_152), .S(n_153), .A(in_14[7]), .B(n_90), .CI(in_3[7]));
  ADDFX1 g6169(.CO(n_150), .S(n_151), .A(n_4), .B(n_70), .CI(in_0[6]));
  ADDFX1 g6170(.CO(n_148), .S(n_149), .A(n_14), .B(in_5[11]), .CI(in_6[11]));
  ADDFX1 g6171(.CO(n_146), .S(n_147), .A(n_68), .B(in_19[3]), .CI(in_3[3]));
  ADDFX1 g6172(.CO(n_144), .S(n_145), .A(n_11), .B(in_11[8]), .CI(in_10[8]));
  ADDFX1 g6173(.CO(n_142), .S(n_143), .A(in_7[8]), .B(n_17), .CI(in_12[8]));
  ADDFX1 g6174(.CO(n_140), .S(n_141), .A(n_15), .B(in_17[7]), .CI(in_9[7]));
  ADDFX1 g6175(.CO(n_138), .S(n_139), .A(n_80), .B(in_8[4]), .CI(in_6[4]));
  ADDFX1 g6176(.CO(n_136), .S(n_137), .A(n_16), .B(in_11[9]), .CI(in_19[9]));
  ADDFX1 g6177(.CO(n_134), .S(n_135), .A(n_49), .B(in_2[7]), .CI(in_8[7]));
  ADDFX1 g6178(.CO(n_132), .S(n_133), .A(n_21), .B(in_2[10]), .CI(in_17[10]));
  INVX1 g6179(.Y(n_130), .A(n_131));
  OAI22X1 g6180(.Y(n_131), .A0(in_8[12]), .A1(n_13), .B0(in_5[12]), .B1(in_6[11]));
  ADDHX1 g6181(.CO(n_128), .S(n_129), .A(in_5[12]), .B(n_9));
  ADDFX1 g6182(.CO(n_126), .S(n_127), .A(in_3[0]), .B(in_5[0]), .CI(in_6[0]));
  ADDFX1 g6183(.CO(n_124), .S(n_125), .A(in_0[8]), .B(in_14[8]), .CI(in_17[8]));
  ADDFX1 g6184(.CO(n_122), .S(n_123), .A(in_15[7]), .B(in_19[7]), .CI(in_13[7]));
  ADDFX1 g6185(.CO(n_120), .S(n_121), .A(in_3[9]), .B(in_2[9]), .CI(in_13[9]));
  ADDFX1 g6186(.CO(n_118), .S(n_119), .A(n_18), .B(in_6[2]), .CI(in_5[2]));
  ADDFX1 g6187(.CO(n_116), .S(n_117), .A(in_0[10]), .B(n_8), .CI(n_7));
  ADDFX1 g6188(.CO(n_114), .S(n_115), .A(in_8[3]), .B(in_5[3]), .CI(in_4[3]));
  ADDFX1 g6189(.CO(n_112), .S(n_113), .A(in_11[4]), .B(in_17[4]), .CI(in_9[4]));
  ADDFX1 g6190(.CO(n_110), .S(n_111), .A(in_6[1]), .B(in_4[1]), .CI(in_5[1]));
  ADDFX1 g6191(.CO(n_108), .S(n_109), .A(in_4[0]), .B(in_15[0]), .CI(in_9[0]));
  ADDFX1 g6192(.CO(n_106), .S(n_107), .A(in_7[9]), .B(in_18[9]), .CI(in_12[9]));
  ADDFX1 g6193(.CO(n_104), .S(n_105), .A(in_16[7]), .B(in_5[7]), .CI(in_4[7]));
  ADDFX1 g6194(.CO(n_102), .S(n_103), .A(in_2[1]), .B(in_16[1]), .CI(in_8[1]));
  ADDFX1 g6195(.CO(n_100), .S(n_101), .A(in_12[1]), .B(in_13[1]), .CI(in_3[1]));
  ADDFX1 g6196(.CO(n_98), .S(n_99), .A(n_6), .B(in_14[4]), .CI(in_12[4]));
  ADDFX1 g6197(.CO(n_96), .S(n_97), .A(in_15[4]), .B(in_16[4]), .CI(in_10[4]));
  ADDFX1 g6198(.CO(n_94), .S(n_95), .A(in_15[6]), .B(in_4[6]), .CI(in_13[6]));
  ADDFX1 g6199(.CO(n_92), .S(n_93), .A(in_17[3]), .B(in_14[3]), .CI(in_12[3]));
  ADDFX1 g6200(.CO(n_90), .S(n_91), .A(in_1[6]), .B(in_7[6]), .CI(in_11[6]));
  ADDFX1 g6201(.CO(n_88), .S(n_89), .A(in_9[10]), .B(in_15[10]), .CI(in_16[10]));
  ADDFX1 g6202(.CO(n_86), .S(n_87), .A(in_13[3]), .B(in_2[3]), .CI(in_6[3]));
  ADDFX1 g6203(.CO(n_84), .S(n_85), .A(in_4[10]), .B(in_8[10]), .CI(in_13[10]));
  ADDFX1 g6204(.CO(n_82), .S(n_83), .A(in_8[2]), .B(in_16[2]), .CI(in_4[2]));
  ADDFX1 g6205(.CO(n_80), .S(n_81), .A(in_1[3]), .B(in_7[3]), .CI(in_18[3]));
  ADDFX1 g6206(.CO(n_78), .S(n_79), .A(in_17[6]), .B(in_9[6]), .CI(in_5[6]));
  ADDFX1 g6207(.CO(n_76), .S(n_77), .A(in_2[2]), .B(in_19[2]), .CI(in_13[2]));
  ADDFX1 g6208(.CO(n_74), .S(n_75), .A(in_1[1]), .B(in_10[1]), .CI(in_11[1]));
  ADDFX1 g6209(.CO(n_72), .S(n_73), .A(in_11[5]), .B(in_17[5]), .CI(in_10[5]));
  ADDFX1 g6210(.CO(n_70), .S(n_71), .A(in_1[5]), .B(in_7[5]), .CI(in_18[5]));
  ADDFX1 g6211(.CO(n_68), .S(n_69), .A(in_1[2]), .B(in_17[2]), .CI(in_0[2]));
  ADDFX1 g6212(.CO(n_66), .S(n_67), .A(in_15[8]), .B(in_2[8]), .CI(in_16[8]));
  ADDFX1 g6213(.CO(n_64), .S(n_65), .A(in_9[3]), .B(in_15[3]), .CI(in_16[3]));
  ADDFX1 g6214(.CO(n_62), .S(n_63), .A(n_1), .B(in_17[0]), .CI(in_19[0]));
  ADDFX1 g6215(.CO(n_60), .S(n_61), .A(in_9[1]), .B(in_14[1]), .CI(in_15[1]));
  ADDFX1 g6216(.CO(n_58), .S(n_59), .A(in_9[5]), .B(in_16[5]), .CI(in_8[5]));
  ADDFX1 g6217(.CO(n_56), .S(n_57), .A(in_0[5]), .B(in_15[5]), .CI(in_2[5]));
  ADDFX1 g6218(.CO(n_54), .S(n_55), .A(in_9[2]), .B(in_12[2]), .CI(in_3[2]));
  ADDFX1 g6219(.CO(n_52), .S(n_53), .A(in_9[8]), .B(in_5[8]), .CI(in_3[8]));
  ADDFX1 g6220(.CO(n_50), .S(n_51), .A(in_0[9]), .B(in_10[9]), .CI(in_17[9]));
  ADDFX1 g6221(.CO(n_48), .S(n_49), .A(in_7[7]), .B(in_18[6]), .CI(in_0[7]));
  ADDFX1 g6222(.CO(n_46), .S(n_47), .A(in_19[5]), .B(in_13[5]), .CI(in_5[5]));
  ADDFX1 g6223(.CO(n_44), .S(n_45), .A(in_15[9]), .B(in_5[9]), .CI(in_8[9]));
  ADDFX1 g6224(.CO(n_42), .S(n_43), .A(in_11[7]), .B(in_12[7]), .CI(in_10[7]));
  ADDFX1 g6225(.CO(n_40), .S(n_41), .A(in_7[2]), .B(in_14[2]), .CI(in_18[2]));
  ADDFX1 g6226(.CO(n_38), .S(n_39), .A(in_0[3]), .B(in_11[3]), .CI(in_10[3]));
  ADDFX1 g6227(.CO(n_36), .S(n_37), .A(in_18[4]), .B(in_14[5]), .CI(in_12[5]));
  ADDFX1 g6228(.CO(n_34), .S(n_35), .A(in_1[4]), .B(in_7[4]), .CI(in_0[4]));
  ADDFX1 g6229(.CO(n_32), .S(n_33), .A(in_4[4]), .B(in_3[4]), .CI(in_19[4]));
  ADDFX1 g6230(.CO(n_30), .S(n_31), .A(in_16[6]), .B(in_8[6]), .CI(in_3[6]));
  ADDFX1 g6231(.CO(n_28), .S(n_29), .A(in_15[2]), .B(in_11[2]), .CI(in_10[2]));
  ADDFX1 g6232(.CO(n_26), .S(n_27), .A(in_14[6]), .B(in_10[6]), .CI(in_12[6]));
  ADDFX1 g6233(.CO(n_24), .S(n_25), .A(in_5[4]), .B(in_2[4]), .CI(in_13[4]));
  OAI21X1 g6234(.Y(n_23), .A0(in_2[11]), .A1(n_12), .B0(n_22));
  NAND2X1 g6236(.Y(n_22), .A(in_2[11]), .B(n_12));
  ADDHX1 g6237(.CO(n_20), .S(n_21), .A(in_12[9]), .B(in_19[10]));
  ADDHX1 g6238(.CO(n_18), .S(n_19), .A(in_17[1]), .B(in_19[1]));
  ADDHX1 g6239(.CO(n_16), .S(n_17), .A(in_1[8]), .B(in_18[8]));
  OAI2BB1X1 g6240(.Y(n_15), .A0N(in_18[7]), .A1N(in_1[7]), .B0(n_11));
  XNOR2X1 g6241(.Y(n_14), .A(in_12[9]), .B(in_14[11]));
  XNOR2X1 g6242(.Y(n_13), .A(in_5[12]), .B(in_6[11]));
  XNOR2X1 g6243(.Y(n_12), .A(in_19[10]), .B(in_0[10]));
  OR2X1 g6244(.Y(n_11), .A(in_18[7]), .B(in_1[7]));
  NOR2BX1 g6245(.Y(n_10), .AN(in_14[11]), .B(in_12[9]));
  NOR2X1 g6246(.Y(n_9), .A(in_19[10]), .B(in_0[10]));
  INVX1 g6247(.Y(n_8), .A(in_11[10]));
  INVX1 g6248(.Y(n_7), .A(in_10[10]));
  INVX1 g6249(.Y(n_6), .A(in_18[4]));
  INVX1 g6250(.Y(n_5), .A(in_13[13]));
  INVX1 g6252(.Y(n_4), .A(in_18[6]));
  INVX1 g6253(.Y(n_3), .A(in_6[11]));
  BUFX2 drc_bufs(.Y(n_1), .A(in_2[0]));
  XOR2XL g2(.Y(n_0), .A(in_8[12]), .B(n_13));
endmodule

module csa_tree_ADD_TC_OP_19_group_2(in_0, in_1, in_2, in_3, in_4, in_5, in_6, 
    in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, 
    in_18, in_19, out_0);
input   [13:0] in_0;
input   [13:0] in_1;
input   [13:0] in_2;
input   [13:0] in_3;
input   [13:0] in_4;
input   [13:0] in_5;
input   [13:0] in_6;
input   [13:0] in_7;
input   [13:0] in_8;
input   [13:0] in_9;
input   [13:0] in_10;
input   [13:0] in_11;
input   [13:0] in_12;
input   [13:0] in_13;
input   [13:0] in_14;
input   [13:0] in_15;
input   [13:0] in_16;
input   [13:0] in_17;
input   [13:0] in_18;
input   [13:0] in_19;
output  [18:0] out_0;
wire  n_402, n_400, n_398, n_396, n_394, n_392, n_390, n_388, n_386, n_384, 
    n_383, n_382, n_380, n_379, n_378, n_377, n_376, n_375, n_374, n_373, 
    n_372, n_370, n_369, n_368, n_367, n_366, n_365, n_364, n_363, n_362, 
    n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, n_352, n_351, 
    n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, n_342, n_341, 
    n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, n_332, n_331, 
    n_330, n_328, n_327, n_326, n_325, n_324, n_323, n_322, n_321, n_320, 
    n_319, n_318, n_317, n_316, n_315, n_314, n_313, n_312, n_311, n_310, 
    n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, n_301, n_300, 
    n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, n_291, n_290, 
    n_289, n_288, n_287, n_286, n_284, n_283, n_282, n_281, n_280, n_279, 
    n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, 
    n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, 
    n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, n_249, 
    n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
    n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_219, n_218, 
    n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
    n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, 
    n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, n_188, 
    n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, 
    n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, 
    n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, 
    n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
    n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
    n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, 
    n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, 
    n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, 
    n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, 
    n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_3, n_2, n_1, n_0;
wire   [18:0] out_0;
wire   [13:0] in_19;
wire   [13:0] in_18;
wire   [13:0] in_17;
wire   [13:0] in_16;
wire   [13:0] in_15;
wire   [13:0] in_14;
wire   [13:0] in_13;
wire   [13:0] in_12;
wire   [13:0] in_11;
wire   [13:0] in_10;
wire   [13:0] in_9;
wire   [13:0] in_8;
wire   [13:0] in_7;
wire   [13:0] in_6;
wire   [13:0] in_5;
wire   [13:0] in_4;
wire   [13:0] in_3;
wire   [13:0] in_2;
wire   [13:0] in_1;
wire   [13:0] in_0;
  assign out_0[17] = 1'b0;
  assign out_0[16] = 1'b0;
  assign out_0[15] = 1'b0;
  OR2X1 g5320(.Y(out_0[18]), .A(n_281), .B(n_402));
  AOI21X1 g5321(.Y(n_402), .A0(n_9), .A1(n_278), .B0(n_400));
  ADDFX1 g5322(.CO(n_400), .S(out_0[14]), .A(n_277), .B(n_346), .CI(n_398));
  ADDFX1 g5323(.CO(n_398), .S(out_0[13]), .A(n_368), .B(n_347), .CI(n_396));
  ADDFX1 g5324(.CO(n_396), .S(out_0[12]), .A(n_372), .B(n_369), .CI(n_394));
  ADDFX1 g5325(.CO(n_394), .S(out_0[11]), .A(n_382), .B(n_373), .CI(n_392));
  ADDFX1 g5326(.CO(n_392), .S(out_0[10]), .A(n_383), .B(n_378), .CI(n_390));
  ADDFX1 g5327(.CO(n_390), .S(out_0[9]), .A(n_376), .B(n_388), .CI(n_379));
  ADDFX1 g5328(.CO(n_388), .S(out_0[8]), .A(n_374), .B(n_377), .CI(n_386));
  ADDFX1 g5329(.CO(n_386), .S(out_0[7]), .A(n_362), .B(n_375), .CI(n_384));
  ADDFX1 g5330(.CO(n_384), .S(out_0[6]), .A(n_366), .B(n_363), .CI(n_380));
  ADDFX1 g5331(.CO(n_382), .S(n_383), .A(n_337), .B(n_364), .CI(n_353));
  ADDFX1 g5332(.CO(n_380), .S(out_0[5]), .A(n_350), .B(n_367), .CI(n_370));
  ADDFX1 g5333(.CO(n_378), .S(n_379), .A(n_343), .B(n_358), .CI(n_365));
  ADDFX1 g5334(.CO(n_376), .S(n_377), .A(n_356), .B(n_345), .CI(n_359));
  ADDFX1 g5335(.CO(n_374), .S(n_375), .A(n_321), .B(n_348), .CI(n_357));
  ADDFX1 g5336(.CO(n_372), .S(n_373), .A(n_336), .B(n_352), .CI(n_355));
  ADDFX1 g5337(.CO(n_370), .S(out_0[4]), .A(n_338), .B(n_360), .CI(n_351));
  ADDFX1 g5338(.CO(n_368), .S(n_369), .A(n_334), .B(n_354), .CI(n_333));
  ADDFX1 g5339(.CO(n_366), .S(n_367), .A(n_340), .B(n_317), .CI(n_331));
  ADDFX1 g5340(.CO(n_364), .S(n_365), .A(n_307), .B(n_344), .CI(n_315));
  ADDFX1 g5341(.CO(n_362), .S(n_363), .A(n_330), .B(n_325), .CI(n_349));
  ADDFX1 g5342(.CO(n_360), .S(out_0[3]), .A(n_297), .B(n_328), .CI(n_339));
  ADDFX1 g5343(.CO(n_358), .S(n_359), .A(n_326), .B(n_320), .CI(n_319));
  ADDFX1 g5344(.CO(n_356), .S(n_357), .A(n_324), .B(n_313), .CI(n_327));
  ADDFX1 g5345(.CO(n_354), .S(n_355), .A(n_322), .B(n_301), .CI(n_335));
  ADDFX1 g5346(.CO(n_352), .S(n_353), .A(n_314), .B(n_323), .CI(n_342));
  ADDFX1 g5347(.CO(n_350), .S(n_351), .A(n_296), .B(n_309), .CI(n_341));
  ADDFX1 g5348(.CO(n_348), .S(n_349), .A(n_293), .B(n_316), .CI(n_305));
  ADDFX1 g5349(.CO(n_346), .S(n_347), .A(n_242), .B(n_275), .CI(n_332));
  ADDFX1 g5350(.CO(n_344), .S(n_345), .A(n_312), .B(n_266), .CI(n_289));
  ADDFX1 g5351(.CO(n_342), .S(n_343), .A(n_288), .B(n_318), .CI(n_311));
  ADDFX1 g5352(.CO(n_340), .S(n_341), .A(n_294), .B(n_260), .CI(n_287));
  ADDFX1 g5353(.CO(n_338), .S(n_339), .A(n_255), .B(n_298), .CI(n_295));
  ADDFX1 g5354(.CO(n_336), .S(n_337), .A(n_306), .B(n_303), .CI(n_272));
  ADDFX1 g5355(.CO(n_334), .S(n_335), .A(n_302), .B(n_271), .CI(n_262));
  ADDFX1 g5356(.CO(n_332), .S(n_333), .A(n_261), .B(n_300), .CI(n_276));
  ADDFX1 g5357(.CO(n_330), .S(n_331), .A(n_308), .B(n_291), .CI(n_274));
  ADDFX1 g5358(.CO(n_328), .S(out_0[2]), .A(n_284), .B(n_256), .CI(n_299));
  ADDFX1 g5359(.CO(n_326), .S(n_327), .A(n_282), .B(n_292), .CI(n_218));
  ADDFX1 g5360(.CO(n_324), .S(n_325), .A(n_290), .B(n_283), .CI(n_273));
  ADDFX1 g5361(.CO(n_322), .S(n_323), .A(n_251), .B(n_230), .CI(n_310));
  ADDFX1 g5362(.CO(n_320), .S(n_321), .A(n_280), .B(n_268), .CI(n_304));
  ADDFX1 g5363(.CO(n_318), .S(n_319), .A(n_279), .B(n_267), .CI(n_270));
  ADDFX1 g5364(.CO(n_316), .S(n_317), .A(n_259), .B(n_286), .CI(n_264));
  ADDFX1 g5365(.CO(n_314), .S(n_315), .A(n_269), .B(n_265), .CI(n_236));
  ADDFX1 g5366(.CO(n_312), .S(n_313), .A(n_234), .B(n_253), .CI(n_204));
  ADDFX1 g5367(.CO(n_310), .S(n_311), .A(n_240), .B(n_249), .CI(n_160));
  ADDFX1 g5368(.CO(n_308), .S(n_309), .A(n_206), .B(n_257), .CI(n_232));
  ADDFX1 g5369(.CO(n_306), .S(n_307), .A(n_243), .B(n_179), .CI(n_252));
  ADDFX1 g5370(.CO(n_304), .S(n_305), .A(n_226), .B(n_263), .CI(n_254));
  ADDFX1 g5371(.CO(n_302), .S(n_303), .A(n_113), .B(n_239), .CI(n_159));
  ADDFX1 g5372(.CO(n_300), .S(n_301), .A(n_139), .B(n_208), .CI(n_229));
  ADDFX1 g5373(.CO(n_298), .S(n_299), .A(n_228), .B(n_221), .CI(n_246));
  ADDFX1 g5374(.CO(n_296), .S(n_297), .A(n_224), .B(n_258), .CI(n_216));
  ADDFX1 g5375(.CO(n_294), .S(n_295), .A(n_227), .B(n_245), .CI(n_176));
  ADDFX1 g5376(.CO(n_292), .S(n_293), .A(n_214), .B(n_237), .CI(n_198));
  ADDFX1 g5377(.CO(n_290), .S(n_291), .A(n_182), .B(n_231), .CI(n_238));
  ADDFX1 g5378(.CO(n_288), .S(n_289), .A(n_250), .B(n_244), .CI(n_180));
  ADDFX1 g5379(.CO(n_286), .S(n_287), .A(n_223), .B(n_215), .CI(n_212));
  ADDFX1 g5380(.CO(n_284), .S(out_0[1]), .A(n_219), .B(n_200), .CI(n_222));
  ADDFX1 g5381(.CO(n_282), .S(n_283), .A(n_209), .B(n_90), .CI(n_247));
  NOR2X1 g5382(.Y(n_281), .A(n_9), .B(n_278));
  ADDFX1 g5383(.CO(n_279), .S(n_280), .A(n_213), .B(n_197), .CI(n_134));
  ADDFX1 g5384(.CO(n_278), .S(n_277), .A(n_26), .B(n_88), .CI(n_241));
  ADDFX1 g5385(.CO(n_275), .S(n_276), .A(n_155), .B(n_207), .CI(n_202));
  ADDFX1 g5386(.CO(n_273), .S(n_274), .A(n_205), .B(n_210), .CI(n_248));
  ADDFX1 g5387(.CO(n_271), .S(n_272), .A(n_140), .B(n_162), .CI(n_235));
  ADDFX1 g5388(.CO(n_269), .S(n_270), .A(n_133), .B(n_233), .CI(n_203));
  ADDFX1 g5389(.CO(n_267), .S(n_268), .A(n_225), .B(n_62), .CI(n_50));
  ADDFX1 g5390(.CO(n_265), .S(n_266), .A(n_148), .B(n_194), .CI(n_217));
  ADDFX1 g5391(.CO(n_263), .S(n_264), .A(n_195), .B(n_144), .CI(n_211));
  ADDFX1 g5392(.CO(n_261), .S(n_262), .A(n_189), .B(n_156), .CI(n_161));
  ADDFX1 g5393(.CO(n_259), .S(n_260), .A(n_178), .B(n_175), .CI(n_196));
  ADDFX1 g5394(.CO(n_257), .S(n_258), .A(n_183), .B(n_172), .CI(n_170));
  ADDFX1 g5395(.CO(n_255), .S(n_256), .A(n_188), .B(n_199), .CI(n_184));
  ADDFX1 g5396(.CO(n_253), .S(n_254), .A(n_181), .B(n_154), .CI(n_40));
  ADDFX1 g5397(.CO(n_251), .S(n_252), .A(n_104), .B(n_193), .CI(n_114));
  ADDFX1 g5398(.CO(n_249), .S(n_250), .A(in_5[8]), .B(n_174), .CI(in_0[8]));
  ADDFX1 g5399(.CO(n_247), .S(n_248), .A(n_177), .B(n_124), .CI(n_102));
  ADDFX1 g5400(.CO(n_245), .S(n_246), .A(n_145), .B(n_164), .CI(n_142));
  ADDFX1 g5401(.CO(n_243), .S(n_244), .A(n_167), .B(n_59), .CI(n_61));
  ADDFX1 g5402(.CO(n_241), .S(n_242), .A(n_97), .B(n_87), .CI(n_201));
  ADDFX1 g5403(.CO(n_239), .S(n_240), .A(n_173), .B(n_55), .CI(in_15[9]));
  ADDFX1 g5404(.CO(n_237), .S(n_238), .A(n_95), .B(n_151), .CI(n_186));
  ADDFX1 g5405(.CO(n_235), .S(n_236), .A(n_71), .B(n_147), .CI(n_192));
  ADDFX1 g5406(.CO(n_233), .S(n_234), .A(n_168), .B(n_35), .CI(n_89));
  ADDFX1 g5407(.CO(n_231), .S(n_232), .A(n_169), .B(n_46), .CI(n_152));
  ADDFX1 g5408(.CO(n_229), .S(n_230), .A(in_0[10]), .B(n_191), .CI(n_190));
  ADDFX1 g5409(.CO(n_227), .S(n_228), .A(n_137), .B(n_165), .CI(n_122));
  ADDFX1 g5410(.CO(n_225), .S(n_226), .A(n_36), .B(n_150), .CI(n_143));
  ADDFX1 g5411(.CO(n_223), .S(n_224), .A(n_163), .B(n_141), .CI(n_126));
  ADDFX1 g5412(.CO(n_221), .S(n_222), .A(n_166), .B(n_157), .CI(n_146));
  ADDFX1 g5413(.CO(n_219), .S(out_0[0]), .A(n_92), .B(n_42), .CI(n_158));
  ADDFX1 g5414(.CO(n_217), .S(n_218), .A(n_153), .B(n_60), .CI(n_39));
  ADDFX1 g5415(.CO(n_215), .S(n_216), .A(n_187), .B(n_68), .CI(n_132));
  ADDFX1 g5416(.CO(n_213), .S(n_214), .A(n_119), .B(n_94), .CI(n_185));
  ADDFX1 g5417(.CO(n_211), .S(n_212), .A(n_112), .B(n_171), .CI(n_67));
  ADDFX1 g5418(.CO(n_209), .S(n_210), .A(n_127), .B(n_45), .CI(n_74));
  ADDFX1 g5419(.CO(n_207), .S(n_208), .A(n_136), .B(in_0[11]), .CI(in_10[11]));
  ADDFX1 g5420(.CO(n_205), .S(n_206), .A(n_128), .B(n_131), .CI(n_96));
  ADDFX1 g5421(.CO(n_203), .S(n_204), .A(n_93), .B(n_149), .CI(in_0[7]));
  ADDFX1 g5422(.CO(n_201), .S(n_202), .A(n_135), .B(in_10[12]), .CI(n_98));
  ADDFX1 g5423(.CO(n_199), .S(n_200), .A(n_86), .B(n_84), .CI(n_138));
  ADDFX1 g5424(.CO(n_197), .S(n_198), .A(n_123), .B(n_73), .CI(n_101));
  ADDFX1 g5425(.CO(n_195), .S(n_196), .A(n_53), .B(n_99), .CI(n_125));
  ADDFX1 g5426(.CO(n_193), .S(n_194), .A(n_110), .B(in_17[8]), .CI(in_10[8]));
  ADDFX1 g5427(.CO(n_191), .S(n_192), .A(n_109), .B(in_16[9]), .CI(n_34));
  ADDFX1 g5428(.CO(n_189), .S(n_190), .A(in_2[10]), .B(n_28), .CI(n_2));
  ADDFX1 g5429(.CO(n_187), .S(n_188), .A(n_66), .B(n_83), .CI(n_85));
  ADDFX1 g5430(.CO(n_185), .S(n_186), .A(n_115), .B(in_3[5]), .CI(in_8[5]));
  ADDFX1 g5431(.CO(n_183), .S(n_184), .A(n_82), .B(n_38), .CI(n_118));
  ADDFX1 g5432(.CO(n_181), .S(n_182), .A(n_111), .B(n_120), .CI(in_0[5]));
  ADDFX1 g5433(.CO(n_179), .S(n_180), .A(n_56), .B(n_49), .CI(n_72));
  ADDFX1 g5434(.CO(n_177), .S(n_178), .A(n_19), .B(n_116), .CI(in_0[4]));
  ADDFX1 g5435(.CO(n_175), .S(n_176), .A(n_54), .B(n_121), .CI(n_100));
  ADDFX1 g5436(.CO(n_173), .S(n_174), .A(n_15), .B(n_107), .CI(in_12[8]));
  ADDFX1 g5437(.CO(n_171), .S(n_172), .A(n_79), .B(n_65), .CI(in_16[3]));
  ADDFX1 g5438(.CO(n_169), .S(n_170), .A(n_37), .B(n_81), .CI(n_117));
  ADDFX1 g5439(.CO(n_167), .S(n_168), .A(n_57), .B(n_108), .CI(in_12[7]));
  ADDFX1 g5440(.CO(n_165), .S(n_166), .A(n_91), .B(n_69), .CI(n_41));
  ADDFX1 g5441(.CO(n_163), .S(n_164), .A(n_77), .B(n_47), .CI(n_80));
  ADDFX1 g5442(.CO(n_161), .S(n_162), .A(n_33), .B(n_31), .CI(in_15[10]));
  ADDFX1 g5443(.CO(n_159), .S(n_160), .A(n_32), .B(in_10[9]), .CI(in_0[9]));
  ADDFX1 g5444(.CO(n_157), .S(n_158), .A(in_0[0]), .B(n_70), .CI(n_52));
  ADDFX1 g5445(.CO(n_155), .S(n_156), .A(in_15[11]), .B(n_21), .CI(n_1));
  ADDFX1 g5446(.CO(n_153), .S(n_154), .A(n_58), .B(in_15[6]), .CI(in_14[6]));
  ADDFX1 g5447(.CO(n_151), .S(n_152), .A(n_63), .B(in_14[4]), .CI(in_10[4]));
  ADDFX1 g5448(.CO(n_149), .S(n_150), .A(n_75), .B(in_9[6]), .CI(in_8[6]));
  ADDFX1 g5449(.CO(n_147), .S(n_148), .A(n_43), .B(in_14[8]), .CI(in_16[8]));
  ADDFX1 g5450(.CO(n_145), .S(n_146), .A(n_106), .B(n_48), .CI(n_78));
  ADDFX1 g5451(.CO(n_143), .S(n_144), .A(n_76), .B(in_15[5]), .CI(in_10[5]));
  ADDFX1 g5452(.CO(n_141), .S(n_142), .A(n_24), .B(n_105), .CI(in_0[2]));
  ADDFX1 g5453(.CO(n_139), .S(n_140), .A(n_103), .B(in_17[10]), .CI(in_10[10]));
  ADDFX1 g5454(.CO(n_137), .S(n_138), .A(in_10[1]), .B(n_25), .CI(n_51));
  INVX1 g5455(.Y(n_136), .A(n_130));
  INVX1 g5456(.Y(n_135), .A(n_129));
  ADDFX1 g5457(.CO(n_133), .S(n_134), .A(n_44), .B(in_14[7]), .CI(in_16[7]));
  ADDFX1 g5458(.CO(n_131), .S(n_132), .A(n_64), .B(in_2[3]), .CI(in_0[3]));
  ADDFX1 g5459(.CO(n_129), .S(n_130), .A(in_2[11]), .B(in_17[11]), .CI(n_17));
  ADDFX1 g5460(.CO(n_127), .S(n_128), .A(n_22), .B(in_12[4]), .CI(in_3[4]));
  ADDFX1 g5461(.CO(n_125), .S(n_126), .A(n_23), .B(in_18[3]), .CI(in_3[3]));
  ADDFX1 g5462(.CO(n_123), .S(n_124), .A(n_10), .B(in_19[5]), .CI(in_2[5]));
  ADDFX1 g5463(.CO(n_121), .S(n_122), .A(in_16[2]), .B(in_19[2]), .CI(in_5[2]));
  ADDFX1 g5464(.CO(n_119), .S(n_120), .A(in_6[5]), .B(in_7[5]), .CI(in_12[5]));
  ADDFX1 g5465(.CO(n_117), .S(n_118), .A(in_14[2]), .B(in_10[2]), .CI(in_3[2]));
  ADDFX1 g5466(.CO(n_115), .S(n_116), .A(in_1[4]), .B(in_7[4]), .CI(in_13[4]));
  ADDFX1 g5467(.CO(n_113), .S(n_114), .A(in_2[9]), .B(in_14[9]), .CI(in_17[9]));
  ADDFX1 g5468(.CO(n_111), .S(n_112), .A(in_9[4]), .B(in_18[4]), .CI(in_19[4]));
  ADDFX1 g5469(.CO(n_109), .S(n_110), .A(in_1[8]), .B(in_4[7]), .CI(in_8[8]));
  ADDFX1 g5470(.CO(n_107), .S(n_108), .A(in_7[7]), .B(in_1[7]), .CI(in_6[7]));
  ADDFX1 g5471(.CO(n_105), .S(n_106), .A(in_9[1]), .B(in_6[1]), .CI(in_12[1]));
  ADDFX1 g5472(.CO(n_103), .S(n_104), .A(in_9[9]), .B(in_19[9]), .CI(in_5[9]));
  ADDFX1 g5473(.CO(n_101), .S(n_102), .A(in_14[5]), .B(in_17[5]), .CI(in_5[5]));
  ADDFX1 g5474(.CO(n_99), .S(n_100), .A(in_5[3]), .B(in_10[3]), .CI(in_8[3]));
  ADDHX1 g5475(.CO(n_97), .S(n_98), .A(n_12), .B(n_27));
  ADDFX1 g5476(.CO(n_95), .S(n_96), .A(in_5[4]), .B(in_15[4]), .CI(in_16[4]));
  ADDFX1 g5477(.CO(n_93), .S(n_94), .A(in_6[6]), .B(in_7[6]), .CI(in_19[6]));
  ADDFX1 g5478(.CO(n_91), .S(n_92), .A(in_5[0]), .B(in_10[0]), .CI(in_14[0]));
  ADDFX1 g5479(.CO(n_89), .S(n_90), .A(in_5[6]), .B(in_16[6]), .CI(in_17[6]));
  OAI22X1 g5480(.Y(n_88), .A0(n_14), .A1(n_30), .B0(in_10[13]), .B1(n_0));
  XOR2XL g5481(.Y(n_87), .A(in_10[13]), .B(n_29));
  ADDFX1 g5482(.CO(n_85), .S(n_86), .A(in_13[1]), .B(in_3[1]), .CI(in_8[1]));
  ADDFX1 g5483(.CO(n_83), .S(n_84), .A(in_0[1]), .B(in_5[1]), .CI(in_19[1]));
  ADDFX1 g5484(.CO(n_81), .S(n_82), .A(in_9[2]), .B(in_12[2]), .CI(in_8[2]));
  ADDFX1 g5485(.CO(n_79), .S(n_80), .A(in_13[2]), .B(in_4[2]), .CI(in_15[2]));
  ADDFX1 g5486(.CO(n_77), .S(n_78), .A(in_15[1]), .B(in_17[1]), .CI(in_18[1]));
  ADDFX1 g5487(.CO(n_75), .S(n_76), .A(in_1[5]), .B(in_4[5]), .CI(in_13[5]));
  ADDFX1 g5488(.CO(n_73), .S(n_74), .A(in_9[5]), .B(in_18[5]), .CI(in_16[5]));
  ADDFX1 g5489(.CO(n_71), .S(n_72), .A(in_19[8]), .B(in_2[8]), .CI(in_15[8]));
  ADDFX1 g5490(.CO(n_69), .S(n_70), .A(in_3[0]), .B(in_8[0]), .CI(in_16[0]));
  ADDFX1 g5491(.CO(n_67), .S(n_68), .A(in_19[3]), .B(in_17[3]), .CI(in_14[3]));
  ADDFX1 g5492(.CO(n_65), .S(n_66), .A(in_6[2]), .B(in_7[2]), .CI(in_1[2]));
  ADDFX1 g5493(.CO(n_63), .S(n_64), .A(in_6[3]), .B(in_7[3]), .CI(in_1[3]));
  ADDFX1 g5494(.CO(n_61), .S(n_62), .A(in_19[7]), .B(in_5[7]), .CI(in_17[7]));
  ADDFX1 g5495(.CO(n_59), .S(n_60), .A(in_9[7]), .B(in_18[7]), .CI(in_3[7]));
  ADDFX1 g5496(.CO(n_57), .S(n_58), .A(in_1[6]), .B(in_4[6]), .CI(in_13[6]));
  ADDFX1 g5497(.CO(n_55), .S(n_56), .A(in_9[8]), .B(in_18[8]), .CI(in_3[8]));
  ADDFX1 g5498(.CO(n_53), .S(n_54), .A(in_15[3]), .B(in_9[3]), .CI(in_12[3]));
  ADDFX1 g5499(.CO(n_51), .S(n_52), .A(n_3), .B(in_17[0]), .CI(in_19[0]));
  ADDFX1 g5500(.CO(n_49), .S(n_50), .A(in_2[7]), .B(in_15[7]), .CI(in_10[7]));
  ADDFX1 g5501(.CO(n_47), .S(n_48), .A(in_4[1]), .B(in_7[1]), .CI(in_14[1]));
  ADDFX1 g5502(.CO(n_45), .S(n_46), .A(in_2[4]), .B(in_8[4]), .CI(in_17[4]));
  ADDFX1 g5503(.CO(n_43), .S(n_44), .A(n_5), .B(in_13[7]), .CI(in_8[7]));
  ADDFX1 g5504(.CO(n_41), .S(n_42), .A(in_6[0]), .B(in_7[0]), .CI(in_13[0]));
  ADDFX1 g5505(.CO(n_39), .S(n_40), .A(in_2[6]), .B(in_10[6]), .CI(in_0[6]));
  ADDFX1 g5506(.CO(n_37), .S(n_38), .A(in_17[2]), .B(in_2[2]), .CI(in_18[2]));
  ADDFX1 g5507(.CO(n_35), .S(n_36), .A(in_12[6]), .B(in_18[6]), .CI(in_3[6]));
  XNOR2X1 g5509(.Y(n_34), .A(in_1[9]), .B(n_18));
  OAI21X1 g5510(.Y(n_33), .A0(n_8), .A1(n_11), .B0(n_7));
  XNOR2X1 g5511(.Y(n_32), .A(n_8), .B(n_16));
  MX2XL g5513(.Y(n_31), .A(in_9[9]), .B(n_6), .S0(n_17));
  NOR2BX1 g5514(.Y(n_30), .AN(in_10[13]), .B(n_27));
  NOR2X1 g5515(.Y(n_29), .A(n_14), .B(n_0));
  NOR2BX1 g5516(.Y(n_28), .AN(in_1[9]), .B(n_18));
  INVX1 g5519(.Y(n_27), .A(n_0));
  INVX1 g5520(.Y(n_26), .A(n_9));
  ADDHX1 g5521(.CO(n_24), .S(n_25), .A(in_2[1]), .B(in_16[1]));
  ADDHX1 g5522(.CO(n_22), .S(n_23), .A(in_4[3]), .B(in_13[3]));
  OAI2BB1X1 g5523(.Y(n_21), .A0N(in_14[10]), .A1N(n_6), .B0(n_20));
  OAI21X1 g5524(.Y(n_20), .A0(in_14[10]), .A1(n_6), .B0(in_16[10]));
  OAI2BB1X1 g5525(.Y(n_19), .A0N(in_4[4]), .A1N(in_6[4]), .B0(n_10));
  XNOR2X1 g5526(.Y(n_18), .A(in_8[8]), .B(in_3[8]));
  XNOR2X1 g5527(.Y(n_17), .A(in_14[10]), .B(in_16[10]));
  XOR2XL g5529(.Y(n_16), .A(in_12[9]), .B(in_18[9]));
  XOR2XL g5530(.Y(n_15), .A(in_4[8]), .B(in_13[8]));
  NOR2X1 g5531(.Y(n_14), .A(in_15[11]), .B(in_0[11]));
  NOR2X1 g5532(.Y(n_13), .A(in_8[8]), .B(in_3[8]));
  NOR2X1 g5533(.Y(n_12), .A(in_14[10]), .B(in_16[10]));
  NOR2X1 g5534(.Y(n_11), .A(in_12[9]), .B(in_18[9]));
  OR2X1 g5535(.Y(n_10), .A(in_4[4]), .B(in_6[4]));
  NAND2X1 g5536(.Y(n_9), .A(in_15[11]), .B(in_0[11]));
  NAND2X1 g5537(.Y(n_8), .A(in_13[8]), .B(in_4[8]));
  NAND2X1 g5538(.Y(n_7), .A(in_12[9]), .B(in_18[9]));
  INVX1 g5539(.Y(n_6), .A(in_9[9]));
  INVX1 g5540(.Y(n_5), .A(in_4[7]));
  BUFX2 drc_bufs(.Y(n_3), .A(in_2[0]));
  XOR2XL g2(.Y(n_2), .A(n_13), .B(n_16));
  AO21XL g5543(.Y(n_1), .A0(n_7), .A1(n_13), .B0(n_11));
  CLKXOR2X1 g5544(.Y(n_0), .A(in_15[11]), .B(in_0[11]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_34, n_32, n_30, 
    n_28, n_26, n_24, n_22, n_20, n_18, n_17, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_44), .S(n_40), .A(n_7), .B(in_3[2]), .CI(n_6));
  ADDFX1 cdnfadd_006_0(.CO(n_45), .S(n_41), .A(n_5), .B(in_3[3]), .CI(n_3));
  ADDFX1 cdnfadd_007_0(.CO(n_46), .S(n_42), .A(n_2), .B(in_3[4]), .CI(n_1));
  ADDFX1 cdnfadd_008_0(.CO(n_47), .S(n_43), .A(n_0), .B(in_3[5]), .CI(n_4));
  NAND3BXL g510(.Y(out_0[13]), .AN(in_3[8]), .B(n_1), .C(n_37));
  XOR2XL g511(.Y(out_0[12]), .A(n_11), .B(n_37));
  ADDFX1 g512(.CO(n_37), .S(out_0[11]), .A(n_9), .B(n_17), .CI(n_34));
  ADDFX1 g513(.CO(n_34), .S(out_0[10]), .A(n_12), .B(n_13), .CI(n_32));
  ADDFX1 g514(.CO(n_32), .S(out_0[9]), .A(n_15), .B(n_47), .CI(n_30));
  ADDFX1 g515(.CO(n_30), .S(out_0[8]), .A(n_46), .B(n_43), .CI(n_28));
  ADDFX1 g516(.CO(n_28), .S(out_0[7]), .A(n_45), .B(n_42), .CI(n_26));
  ADDFX1 g517(.CO(n_26), .S(out_0[6]), .A(n_44), .B(n_41), .CI(n_24));
  ADDFX1 g518(.CO(n_24), .S(out_0[5]), .A(n_10), .B(n_40), .CI(n_22));
  ADDFX1 g519(.CO(n_22), .S(out_0[4]), .A(in_3[1]), .B(n_14), .CI(n_20));
  ADDFX1 g520(.CO(n_20), .S(out_0[3]), .A(n_2), .B(in_3[0]), .CI(n_18));
  AOI2BB1X1 g521(.Y(out_0[2]), .A0N(n_5), .A1N(n_8), .B0(n_18));
  AND2XL g522(.Y(n_18), .A(n_5), .B(n_8));
  AOI21X1 g523(.Y(n_17), .A0(in_3[7]), .A1(in_3[8]), .B0(n_11));
  AOI21X1 g524(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_8));
  OAI2BB1X1 g525(.Y(n_15), .A0N(in_3[6]), .A1N(n_6), .B0(n_12));
  OAI21X1 g526(.Y(n_14), .A0(in_3[4]), .A1(in_3[0]), .B0(n_10));
  OAI2BB1X1 g527(.Y(n_13), .A0N(in_3[7]), .A1N(n_3), .B0(n_9));
  NAND2X1 g528(.Y(n_12), .A(in_3[5]), .B(n_3));
  NOR2X1 g529(.Y(n_11), .A(in_3[7]), .B(in_3[8]));
  NAND2X1 g530(.Y(n_10), .A(in_3[4]), .B(in_3[0]));
  NAND2X1 g531(.Y(n_9), .A(in_3[6]), .B(n_1));
  NOR2XL g532(.Y(n_8), .A(in_3[1]), .B(in_3[0]));
  INVX1 g533(.Y(n_7), .A(in_3[1]));
  INVX1 g534(.Y(n_6), .A(in_3[5]));
  INVX1 g535(.Y(n_5), .A(in_3[2]));
  INVX1 g536(.Y(n_4), .A(in_3[8]));
  INVX1 g537(.Y(n_3), .A(in_3[6]));
  INVX1 g538(.Y(n_2), .A(in_3[3]));
  INVX1 g539(.Y(n_1), .A(in_3[7]));
  INVX1 g540(.Y(n_0), .A(in_3[4]));
endmodule

module csa_tree_SUB_TC_OP_4_group_1752(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [12:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
    n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_35, n_33, n_31, n_29, n_27, 
    n_25, n_23, n_21, n_20, n_19, n_18, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [12:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[11] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_004_1(.CO(n_53), .S(n_46), .A(in_3[3]), .B(n_3), .CI(n_13));
  ADDFX1 cdnfadd_005_0(.CO(n_45), .S(n_44), .A(n_7), .B(in_3[5]), .CI(in_3[4]));
  ADDFX1 cdnfadd_005_1(.CO(n_54), .S(n_47), .A(in_3[2]), .B(n_14), .CI(n_44));
  ADDFX1 cdnfadd_006_0(.CO(n_43), .S(n_42), .A(n_2), .B(in_3[6]), .CI(in_3[5]));
  ADDFX1 cdnfadd_006_1(.CO(n_55), .S(n_48), .A(in_3[3]), .B(n_45), .CI(n_42));
  ADDFX1 cdnfadd_007_0(.CO(n_41), .S(n_40), .A(n_1), .B(in_3[7]), .CI(in_3[6]));
  ADDFX1 cdnfadd_007_1(.CO(n_56), .S(n_49), .A(in_3[4]), .B(n_43), .CI(n_40));
  ADDFX1 cdnfadd_008_1(.CO(n_51), .S(n_50), .A(n_6), .B(n_41), .CI(n_18));
  ADDFX1 cdnfadd_009_0(.CO(n_52), .S(n_57), .A(n_5), .B(in_3[6]), .CI(n_12));
  OAI2BB1X1 g525(.Y(out_0[13]), .A0N(in_3[7]), .A1N(n_10), .B0(n_37));
  ADDFX1 g526(.CO(n_37), .S(out_0[10]), .A(n_15), .B(n_52), .CI(n_35));
  ADDFX1 g527(.CO(n_35), .S(out_0[9]), .A(n_57), .B(n_51), .CI(n_33));
  ADDFX1 g528(.CO(n_33), .S(out_0[8]), .A(n_56), .B(n_50), .CI(n_31));
  ADDFX1 g529(.CO(n_31), .S(out_0[7]), .A(n_55), .B(n_49), .CI(n_29));
  ADDFX1 g530(.CO(n_29), .S(out_0[6]), .A(n_54), .B(n_48), .CI(n_27));
  ADDFX1 g531(.CO(n_27), .S(out_0[5]), .A(n_53), .B(n_25), .CI(n_47));
  ADDFX1 g532(.CO(n_25), .S(out_0[4]), .A(n_16), .B(n_23), .CI(n_46));
  ADDFX1 g533(.CO(n_23), .S(out_0[3]), .A(in_3[2]), .B(n_19), .CI(n_21));
  CLKXOR2X1 g534(.Y(out_0[2]), .A(n_11), .B(n_20));
  NAND2XL g535(.Y(n_21), .A(n_8), .B(n_11));
  OAI2BB1X1 g536(.Y(n_20), .A0N(n_7), .A1N(n_2), .B0(n_8));
  AOI21X1 g537(.Y(n_19), .A0(n_1), .A1(n_3), .B0(n_13));
  AOI21X1 g538(.Y(n_18), .A0(n_5), .A1(n_4), .B0(n_12));
  OA21X1 g539(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_11));
  OAI2BB1X1 g540(.Y(n_16), .A0N(in_3[1]), .A1N(in_3[4]), .B0(n_14));
  AOI21X1 g541(.Y(n_15), .A0(in_3[6]), .A1(n_4), .B0(n_9));
  NAND2X1 g542(.Y(n_14), .A(n_7), .B(n_6));
  NOR2X1 g543(.Y(n_13), .A(n_1), .B(n_3));
  NOR2X1 g544(.Y(n_12), .A(n_5), .B(n_4));
  NAND2X1 g545(.Y(n_11), .A(in_3[0]), .B(in_3[1]));
  INVXL g546(.Y(n_10), .A(n_9));
  NOR2X1 g547(.Y(n_9), .A(in_3[6]), .B(n_4));
  NAND2X1 g548(.Y(n_8), .A(in_3[1]), .B(in_3[2]));
  INVX1 g549(.Y(n_7), .A(in_3[1]));
  INVX1 g550(.Y(n_6), .A(in_3[4]));
  INVX1 g551(.Y(n_5), .A(in_3[5]));
  INVX1 g552(.Y(n_4), .A(in_3[7]));
  INVX1 g553(.Y(n_3), .A(in_3[0]));
  INVX1 g554(.Y(n_2), .A(in_3[2]));
  INVX1 g555(.Y(n_1), .A(in_3[3]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_1(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_34, n_32, n_30, 
    n_28, n_26, n_24, n_22, n_20, n_18, n_17, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_44), .S(n_40), .A(n_7), .B(in_3[2]), .CI(n_6));
  ADDFX1 cdnfadd_006_0(.CO(n_45), .S(n_41), .A(n_5), .B(in_3[3]), .CI(n_3));
  ADDFX1 cdnfadd_007_0(.CO(n_46), .S(n_42), .A(n_2), .B(in_3[4]), .CI(n_1));
  ADDFX1 cdnfadd_008_0(.CO(n_47), .S(n_43), .A(n_0), .B(in_3[5]), .CI(n_4));
  NAND3BXL g510(.Y(out_0[13]), .AN(in_3[8]), .B(n_1), .C(n_37));
  XOR2XL g511(.Y(out_0[12]), .A(n_11), .B(n_37));
  ADDFX1 g512(.CO(n_37), .S(out_0[11]), .A(n_9), .B(n_17), .CI(n_34));
  ADDFX1 g513(.CO(n_34), .S(out_0[10]), .A(n_12), .B(n_13), .CI(n_32));
  ADDFX1 g514(.CO(n_32), .S(out_0[9]), .A(n_15), .B(n_47), .CI(n_30));
  ADDFX1 g515(.CO(n_30), .S(out_0[8]), .A(n_46), .B(n_43), .CI(n_28));
  ADDFX1 g516(.CO(n_28), .S(out_0[7]), .A(n_45), .B(n_42), .CI(n_26));
  ADDFX1 g517(.CO(n_26), .S(out_0[6]), .A(n_44), .B(n_41), .CI(n_24));
  ADDFX1 g518(.CO(n_24), .S(out_0[5]), .A(n_10), .B(n_40), .CI(n_22));
  ADDFX1 g519(.CO(n_22), .S(out_0[4]), .A(in_3[1]), .B(n_14), .CI(n_20));
  ADDFX1 g520(.CO(n_20), .S(out_0[3]), .A(n_2), .B(in_3[0]), .CI(n_18));
  AOI2BB1X1 g521(.Y(out_0[2]), .A0N(n_5), .A1N(n_8), .B0(n_18));
  AND2XL g522(.Y(n_18), .A(n_5), .B(n_8));
  AOI21X1 g523(.Y(n_17), .A0(in_3[7]), .A1(in_3[8]), .B0(n_11));
  AOI21X1 g524(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_8));
  OAI2BB1X1 g525(.Y(n_15), .A0N(in_3[6]), .A1N(n_6), .B0(n_12));
  OAI21X1 g526(.Y(n_14), .A0(in_3[4]), .A1(in_3[0]), .B0(n_10));
  OAI2BB1X1 g527(.Y(n_13), .A0N(in_3[7]), .A1N(n_3), .B0(n_9));
  NAND2X1 g528(.Y(n_12), .A(in_3[5]), .B(n_3));
  NOR2X1 g529(.Y(n_11), .A(in_3[7]), .B(in_3[8]));
  NAND2X1 g530(.Y(n_10), .A(in_3[0]), .B(in_3[4]));
  NAND2X1 g531(.Y(n_9), .A(in_3[6]), .B(n_1));
  NOR2X1 g532(.Y(n_8), .A(in_3[0]), .B(in_3[1]));
  INVX1 g533(.Y(n_7), .A(in_3[1]));
  INVX1 g534(.Y(n_6), .A(in_3[5]));
  INVX1 g535(.Y(n_5), .A(in_3[2]));
  INVX1 g536(.Y(n_4), .A(in_3[8]));
  INVX1 g537(.Y(n_3), .A(in_3[6]));
  INVX1 g538(.Y(n_2), .A(in_3[3]));
  INVX1 g539(.Y(n_1), .A(in_3[7]));
  INVX1 g540(.Y(n_0), .A(in_3[4]));
endmodule

module csa_tree_SUB_TC_OP_3_group_11408(in_0, in_1, in_2, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
output  [13:0] out_0;
wire  n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, 
    n_20, n_19, n_18, n_17, n_14, n_13, n_12, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[1] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd3(.CO(n_22), .S(out_0[3]), .A(in_2[2]), .B(in_2[3]), .CI(n_9));
  ADDFX1 cdnfadd4(.CO(n_21), .S(out_0[4]), .A(in_2[4]), .B(n_12), .CI(n_22));
  ADDFX1 cdnfadd5(.CO(n_20), .S(out_0[5]), .A(n_8), .B(n_23), .CI(n_21));
  ADDFX1 cdnfadd6(.CO(n_19), .S(out_0[6]), .A(n_29), .B(n_24), .CI(n_20));
  ADDFX1 cdnfadd7(.CO(n_18), .S(out_0[7]), .A(n_30), .B(n_25), .CI(n_19));
  ADDFX1 cdnfadd8(.CO(n_17), .S(out_0[8]), .A(n_31), .B(n_26), .CI(n_18));
  ADDFX1 cdnfadd9(.CO(n_28), .S(out_0[9]), .A(n_32), .B(n_10), .CI(n_17));
  ADDFX1 cdnfadd10(.CO(n_27), .S(out_0[10]), .A(n_2), .B(n_7), .CI(n_28));
  ADDFX1 cdnfadd_005_0(.CO(n_29), .S(n_23), .A(n_4), .B(in_2[5]), .CI(in_2[4]));
  ADDFX1 cdnfadd_006_0(.CO(n_30), .S(n_24), .A(n_5), .B(in_2[6]), .CI(in_2[5]));
  ADDFX1 cdnfadd_007_0(.CO(n_31), .S(n_25), .A(n_6), .B(in_2[7]), .CI(in_2[6]));
  ADDFX1 cdnfadd_008_0(.CO(n_32), .S(n_26), .A(n_1), .B(in_2[8]), .CI(in_2[7]));
  AOI21X1 g294(.Y(out_0[11]), .A0(in_2[8]), .A1(n_13), .B0(n_14));
  INVX1 g295(.Y(out_0[13]), .A(n_14));
  NOR2X1 g296(.Y(n_14), .A(in_2[8]), .B(n_13));
  INVX1 g297(.Y(n_13), .A(n_27));
  OAI21X1 g298(.Y(n_12), .A0(in_2[1]), .A1(n_5), .B0(n_8));
  AOI2BB1X1 g299(.Y(out_0[2]), .A0N(in_2[2]), .A1N(in_2[1]), .B0(n_9));
  AOI21X1 g300(.Y(n_10), .A0(in_2[6]), .A1(n_3), .B0(n_7));
  AND2XL g301(.Y(n_9), .A(in_2[2]), .B(in_2[1]));
  NAND2X1 g302(.Y(n_8), .A(n_5), .B(in_2[1]));
  NOR2X1 g303(.Y(n_7), .A(in_2[6]), .B(n_3));
  INVX1 g304(.Y(n_6), .A(in_2[4]));
  INVX1 g305(.Y(n_5), .A(in_2[3]));
  INVX1 g306(.Y(n_4), .A(in_2[2]));
  INVX1 g307(.Y(n_3), .A(in_2[8]));
  INVX1 g308(.Y(n_2), .A(in_2[7]));
  INVX1 g309(.Y(n_1), .A(in_2[5]));
endmodule

module csa_tree_SUB_TC_OP_4_group_1752_1(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [12:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
    n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_35, n_33, n_31, n_29, n_27, 
    n_25, n_23, n_21, n_20, n_19, n_18, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [12:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[11] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_004_1(.CO(n_53), .S(n_46), .A(in_3[3]), .B(n_3), .CI(n_13));
  ADDFX1 cdnfadd_005_0(.CO(n_45), .S(n_44), .A(n_7), .B(in_3[5]), .CI(in_3[4]));
  ADDFX1 cdnfadd_005_1(.CO(n_54), .S(n_47), .A(in_3[2]), .B(n_14), .CI(n_44));
  ADDFX1 cdnfadd_006_0(.CO(n_43), .S(n_42), .A(n_2), .B(in_3[6]), .CI(in_3[5]));
  ADDFX1 cdnfadd_006_1(.CO(n_55), .S(n_48), .A(in_3[3]), .B(n_45), .CI(n_42));
  ADDFX1 cdnfadd_007_0(.CO(n_41), .S(n_40), .A(n_1), .B(in_3[7]), .CI(in_3[6]));
  ADDFX1 cdnfadd_007_1(.CO(n_56), .S(n_49), .A(in_3[4]), .B(n_43), .CI(n_40));
  ADDFX1 cdnfadd_008_1(.CO(n_51), .S(n_50), .A(n_6), .B(n_41), .CI(n_18));
  ADDFX1 cdnfadd_009_0(.CO(n_52), .S(n_57), .A(n_5), .B(in_3[6]), .CI(n_12));
  OAI2BB1X1 g525(.Y(out_0[13]), .A0N(in_3[7]), .A1N(n_10), .B0(n_37));
  ADDFX1 g526(.CO(n_37), .S(out_0[10]), .A(n_15), .B(n_52), .CI(n_35));
  ADDFX1 g527(.CO(n_35), .S(out_0[9]), .A(n_57), .B(n_51), .CI(n_33));
  ADDFX1 g528(.CO(n_33), .S(out_0[8]), .A(n_56), .B(n_50), .CI(n_31));
  ADDFX1 g529(.CO(n_31), .S(out_0[7]), .A(n_55), .B(n_49), .CI(n_29));
  ADDFX1 g530(.CO(n_29), .S(out_0[6]), .A(n_54), .B(n_48), .CI(n_27));
  ADDFX1 g531(.CO(n_27), .S(out_0[5]), .A(n_53), .B(n_25), .CI(n_47));
  ADDFX1 g532(.CO(n_25), .S(out_0[4]), .A(n_16), .B(n_23), .CI(n_46));
  ADDFX1 g533(.CO(n_23), .S(out_0[3]), .A(in_3[2]), .B(n_19), .CI(n_21));
  XOR2XL g534(.Y(out_0[2]), .A(n_11), .B(n_20));
  NAND2XL g535(.Y(n_21), .A(n_11), .B(n_8));
  OAI2BB1X1 g536(.Y(n_20), .A0N(n_7), .A1N(n_2), .B0(n_8));
  AOI21X1 g537(.Y(n_19), .A0(n_1), .A1(n_3), .B0(n_13));
  AOI21X1 g538(.Y(n_18), .A0(n_5), .A1(n_4), .B0(n_12));
  OA21X1 g539(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_11));
  OAI2BB1X1 g540(.Y(n_16), .A0N(in_3[1]), .A1N(in_3[4]), .B0(n_14));
  AOI21X1 g541(.Y(n_15), .A0(in_3[6]), .A1(n_4), .B0(n_9));
  NAND2X1 g542(.Y(n_14), .A(n_7), .B(n_6));
  NOR2X1 g543(.Y(n_13), .A(n_1), .B(n_3));
  NOR2X1 g544(.Y(n_12), .A(n_5), .B(n_4));
  NAND2X1 g545(.Y(n_11), .A(in_3[0]), .B(in_3[1]));
  INVXL g546(.Y(n_10), .A(n_9));
  NOR2X1 g547(.Y(n_9), .A(in_3[6]), .B(n_4));
  NAND2X1 g548(.Y(n_8), .A(in_3[1]), .B(in_3[2]));
  INVX1 g549(.Y(n_7), .A(in_3[1]));
  INVX1 g550(.Y(n_6), .A(in_3[4]));
  INVX1 g551(.Y(n_5), .A(in_3[5]));
  INVX1 g552(.Y(n_4), .A(in_3[7]));
  INVX1 g553(.Y(n_3), .A(in_3[0]));
  INVX1 g554(.Y(n_2), .A(in_3[2]));
  INVX1 g555(.Y(n_1), .A(in_3[3]));
endmodule

module csa_tree_SUB_TC_OP_4_group_1752_2(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [12:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
    n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_35, n_33, n_31, n_29, n_27, 
    n_25, n_23, n_21, n_20, n_19, n_18, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [12:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[11] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_004_1(.CO(n_53), .S(n_46), .A(in_3[3]), .B(n_3), .CI(n_13));
  ADDFX1 cdnfadd_005_0(.CO(n_45), .S(n_44), .A(n_7), .B(in_3[5]), .CI(in_3[4]));
  ADDFX1 cdnfadd_005_1(.CO(n_54), .S(n_47), .A(in_3[2]), .B(n_14), .CI(n_44));
  ADDFX1 cdnfadd_006_0(.CO(n_43), .S(n_42), .A(n_2), .B(in_3[6]), .CI(in_3[5]));
  ADDFX1 cdnfadd_006_1(.CO(n_55), .S(n_48), .A(in_3[3]), .B(n_45), .CI(n_42));
  ADDFX1 cdnfadd_007_0(.CO(n_41), .S(n_40), .A(n_1), .B(in_3[7]), .CI(in_3[6]));
  ADDFX1 cdnfadd_007_1(.CO(n_56), .S(n_49), .A(in_3[4]), .B(n_43), .CI(n_40));
  ADDFX1 cdnfadd_008_1(.CO(n_51), .S(n_50), .A(n_6), .B(n_41), .CI(n_18));
  ADDFX1 cdnfadd_009_0(.CO(n_52), .S(n_57), .A(n_5), .B(in_3[6]), .CI(n_12));
  OAI2BB1X1 g525(.Y(out_0[13]), .A0N(in_3[7]), .A1N(n_10), .B0(n_37));
  ADDFX1 g526(.CO(n_37), .S(out_0[10]), .A(n_15), .B(n_52), .CI(n_35));
  ADDFX1 g527(.CO(n_35), .S(out_0[9]), .A(n_57), .B(n_51), .CI(n_33));
  ADDFX1 g528(.CO(n_33), .S(out_0[8]), .A(n_56), .B(n_50), .CI(n_31));
  ADDFX1 g529(.CO(n_31), .S(out_0[7]), .A(n_55), .B(n_49), .CI(n_29));
  ADDFX1 g530(.CO(n_29), .S(out_0[6]), .A(n_54), .B(n_48), .CI(n_27));
  ADDFX1 g531(.CO(n_27), .S(out_0[5]), .A(n_53), .B(n_25), .CI(n_47));
  ADDFX1 g532(.CO(n_25), .S(out_0[4]), .A(n_16), .B(n_23), .CI(n_46));
  ADDFX1 g533(.CO(n_23), .S(out_0[3]), .A(in_3[2]), .B(n_19), .CI(n_21));
  XOR2XL g534(.Y(out_0[2]), .A(n_11), .B(n_20));
  NAND2X1 g535(.Y(n_21), .A(n_11), .B(n_8));
  OAI2BB1X1 g536(.Y(n_20), .A0N(n_7), .A1N(n_2), .B0(n_8));
  AOI21X1 g537(.Y(n_19), .A0(n_1), .A1(n_3), .B0(n_13));
  AOI21X1 g538(.Y(n_18), .A0(n_5), .A1(n_4), .B0(n_12));
  OA21X1 g539(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_11));
  OAI2BB1X1 g540(.Y(n_16), .A0N(in_3[4]), .A1N(in_3[1]), .B0(n_14));
  AOI21X1 g541(.Y(n_15), .A0(in_3[6]), .A1(n_4), .B0(n_9));
  NAND2X1 g542(.Y(n_14), .A(n_6), .B(n_7));
  NOR2X1 g543(.Y(n_13), .A(n_1), .B(n_3));
  NOR2X1 g544(.Y(n_12), .A(n_5), .B(n_4));
  NAND2X1 g545(.Y(n_11), .A(in_3[0]), .B(in_3[1]));
  INVXL g546(.Y(n_10), .A(n_9));
  NOR2X1 g547(.Y(n_9), .A(in_3[6]), .B(n_4));
  NAND2X1 g548(.Y(n_8), .A(in_3[1]), .B(in_3[2]));
  INVX1 g549(.Y(n_7), .A(in_3[1]));
  INVX1 g550(.Y(n_6), .A(in_3[4]));
  INVX1 g551(.Y(n_5), .A(in_3[5]));
  INVX1 g552(.Y(n_4), .A(in_3[7]));
  INVX1 g553(.Y(n_3), .A(in_3[0]));
  INVX1 g554(.Y(n_2), .A(in_3[2]));
  INVX1 g555(.Y(n_1), .A(in_3[3]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_2(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_34, n_32, n_30, 
    n_28, n_26, n_24, n_22, n_20, n_18, n_17, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_44), .S(n_40), .A(n_7), .B(in_3[2]), .CI(n_6));
  ADDFX1 cdnfadd_006_0(.CO(n_45), .S(n_41), .A(n_5), .B(in_3[3]), .CI(n_3));
  ADDFX1 cdnfadd_007_0(.CO(n_46), .S(n_42), .A(n_2), .B(in_3[4]), .CI(n_1));
  ADDFX1 cdnfadd_008_0(.CO(n_47), .S(n_43), .A(n_0), .B(in_3[5]), .CI(n_4));
  NAND3BXL g510(.Y(out_0[13]), .AN(in_3[8]), .B(n_1), .C(n_37));
  XOR2XL g511(.Y(out_0[12]), .A(n_11), .B(n_37));
  ADDFX1 g512(.CO(n_37), .S(out_0[11]), .A(n_9), .B(n_17), .CI(n_34));
  ADDFX1 g513(.CO(n_34), .S(out_0[10]), .A(n_12), .B(n_13), .CI(n_32));
  ADDFX1 g514(.CO(n_32), .S(out_0[9]), .A(n_15), .B(n_47), .CI(n_30));
  ADDFX1 g515(.CO(n_30), .S(out_0[8]), .A(n_46), .B(n_43), .CI(n_28));
  ADDFX1 g516(.CO(n_28), .S(out_0[7]), .A(n_45), .B(n_42), .CI(n_26));
  ADDFX1 g517(.CO(n_26), .S(out_0[6]), .A(n_44), .B(n_41), .CI(n_24));
  ADDFX1 g518(.CO(n_24), .S(out_0[5]), .A(n_10), .B(n_40), .CI(n_22));
  ADDFX1 g519(.CO(n_22), .S(out_0[4]), .A(in_3[1]), .B(n_14), .CI(n_20));
  ADDFX1 g520(.CO(n_20), .S(out_0[3]), .A(n_2), .B(in_3[0]), .CI(n_18));
  AOI2BB1XL g521(.Y(out_0[2]), .A0N(n_5), .A1N(n_8), .B0(n_18));
  AND2XL g522(.Y(n_18), .A(n_5), .B(n_8));
  AOI21X1 g523(.Y(n_17), .A0(in_3[7]), .A1(in_3[8]), .B0(n_11));
  AOI21X1 g524(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_8));
  OAI2BB1X1 g525(.Y(n_15), .A0N(in_3[6]), .A1N(n_6), .B0(n_12));
  OAI21X1 g526(.Y(n_14), .A0(in_3[4]), .A1(in_3[0]), .B0(n_10));
  OAI2BB1X1 g527(.Y(n_13), .A0N(in_3[7]), .A1N(n_3), .B0(n_9));
  NAND2X1 g528(.Y(n_12), .A(in_3[5]), .B(n_3));
  NOR2X1 g529(.Y(n_11), .A(in_3[7]), .B(in_3[8]));
  NAND2X1 g530(.Y(n_10), .A(in_3[4]), .B(in_3[0]));
  NAND2X1 g531(.Y(n_9), .A(in_3[6]), .B(n_1));
  NOR2X1 g532(.Y(n_8), .A(in_3[1]), .B(in_3[0]));
  INVX1 g533(.Y(n_7), .A(in_3[1]));
  INVX1 g534(.Y(n_6), .A(in_3[5]));
  INVX1 g535(.Y(n_5), .A(in_3[2]));
  INVX1 g536(.Y(n_4), .A(in_3[8]));
  INVX1 g537(.Y(n_3), .A(in_3[6]));
  INVX1 g538(.Y(n_2), .A(in_3[3]));
  INVX1 g539(.Y(n_1), .A(in_3[7]));
  INVX1 g540(.Y(n_0), .A(in_3[4]));
endmodule

module csa_tree_SUB_TC_OP_3_group_11408_1(in_0, in_1, in_2, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
output  [13:0] out_0;
wire  n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, 
    n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_17, n_16, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_1, n_0;
wire   [13:0] out_0;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[1] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd3(.CO(n_26), .S(out_0[3]), .A(in_2[2]), .B(in_2[3]), .CI(n_11));
  ADDFX1 cdnfadd4(.CO(n_25), .S(out_0[4]), .A(in_2[4]), .B(n_14), .CI(n_26));
  ADDFX1 cdnfadd5(.CO(n_24), .S(out_0[5]), .A(n_10), .B(n_27), .CI(n_25));
  ADDFX1 cdnfadd6(.CO(n_23), .S(out_0[6]), .A(n_35), .B(n_28), .CI(n_24));
  ADDFX1 cdnfadd7(.CO(n_22), .S(out_0[7]), .A(n_36), .B(n_29), .CI(n_23));
  ADDFX1 cdnfadd8(.CO(n_21), .S(out_0[8]), .A(n_37), .B(n_30), .CI(n_22));
  ADDFX1 cdnfadd9(.CO(n_34), .S(out_0[9]), .A(n_38), .B(n_31), .CI(n_21));
  ADDFX1 cdnfadd10(.CO(n_33), .S(out_0[10]), .A(n_13), .B(n_32), .CI(n_34));
  ADDFX1 cdnfadd11(.CO(n_20), .S(out_0[11]), .A(n_6), .B(n_12), .CI(n_33));
  ADDFX1 cdnfadd_005_0(.CO(n_35), .S(n_27), .A(n_7), .B(in_2[5]), .CI(in_2[4]));
  ADDFX1 cdnfadd_006_0(.CO(n_36), .S(n_28), .A(n_8), .B(in_2[6]), .CI(in_2[5]));
  ADDFX1 cdnfadd_007_0(.CO(n_37), .S(n_29), .A(n_9), .B(in_2[7]), .CI(in_2[6]));
  ADDFX1 cdnfadd_008_0(.CO(n_38), .S(n_30), .A(n_4), .B(in_2[8]), .CI(in_2[7]));
  ADDFX1 cdnfadd_009_0(.CO(n_32), .S(n_31), .A(n_5), .B(in_2[9]), .CI(in_2[8]));
  AOI21X1 g230(.Y(out_0[12]), .A0(in_2[9]), .A1(n_16), .B0(n_17));
  INVX1 g231(.Y(out_0[13]), .A(n_17));
  NOR2X1 g232(.Y(n_17), .A(in_2[9]), .B(n_16));
  INVX1 g233(.Y(n_16), .A(n_20));
  AOI2BB1X1 g234(.Y(out_0[2]), .A0N(in_2[2]), .A1N(n_1), .B0(n_11));
  OAI21X1 g235(.Y(n_14), .A0(n_8), .A1(n_1), .B0(n_10));
  AOI21X1 g236(.Y(n_13), .A0(in_2[7]), .A1(n_3), .B0(n_12));
  NOR2X1 g237(.Y(n_12), .A(in_2[7]), .B(n_3));
  AND2XL g238(.Y(n_11), .A(in_2[2]), .B(n_1));
  NAND2X1 g239(.Y(n_10), .A(n_8), .B(n_1));
  INVX1 g240(.Y(n_9), .A(in_2[4]));
  INVX1 g241(.Y(n_8), .A(in_2[3]));
  INVX1 g242(.Y(n_7), .A(in_2[2]));
  INVX1 g243(.Y(n_6), .A(in_2[8]));
  INVX1 g244(.Y(n_5), .A(in_2[6]));
  INVX1 g245(.Y(n_4), .A(in_2[5]));
  INVX1 g246(.Y(n_3), .A(in_2[9]));
  INVX1 drc_bufs(.Y(n_1), .A(n_0));
  INVX1 drc_bufs248(.Y(n_0), .A(in_2[1]));
endmodule

module csa_tree_SUB_TC_OP_3_group_11408_2(in_0, in_1, in_2, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
output  [13:0] out_0;
wire  n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_15, n_14, n_12, n_11, n_10, 
    n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[1] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd3(.CO(n_24), .S(out_0[3]), .A(in_2[2]), .B(in_2[3]), .CI(n_9));
  ADDFX1 cdnfadd4(.CO(n_23), .S(out_0[4]), .A(in_2[4]), .B(n_12), .CI(n_24));
  ADDFX1 cdnfadd5(.CO(n_22), .S(out_0[5]), .A(n_8), .B(n_25), .CI(n_23));
  ADDFX1 cdnfadd6(.CO(n_21), .S(out_0[6]), .A(n_33), .B(n_26), .CI(n_22));
  ADDFX1 cdnfadd7(.CO(n_20), .S(out_0[7]), .A(n_34), .B(n_27), .CI(n_21));
  ADDFX1 cdnfadd8(.CO(n_19), .S(out_0[8]), .A(n_35), .B(n_28), .CI(n_20));
  ADDFX1 cdnfadd9(.CO(n_32), .S(out_0[9]), .A(n_36), .B(n_29), .CI(n_19));
  ADDFX1 cdnfadd10(.CO(n_31), .S(out_0[10]), .A(n_11), .B(n_30), .CI(n_32));
  ADDFX1 cdnfadd11(.CO(n_18), .S(out_0[11]), .A(n_4), .B(n_10), .CI(n_31));
  ADDFX1 cdnfadd_005_0(.CO(n_33), .S(n_25), .A(n_5), .B(in_2[5]), .CI(in_2[4]));
  ADDFX1 cdnfadd_006_0(.CO(n_34), .S(n_26), .A(n_6), .B(in_2[6]), .CI(in_2[5]));
  ADDFX1 cdnfadd_007_0(.CO(n_35), .S(n_27), .A(n_7), .B(in_2[7]), .CI(in_2[6]));
  ADDFX1 cdnfadd_008_0(.CO(n_36), .S(n_28), .A(n_2), .B(in_2[8]), .CI(in_2[7]));
  ADDFX1 cdnfadd_009_0(.CO(n_30), .S(n_29), .A(n_3), .B(in_2[9]), .CI(in_2[8]));
  AOI21X1 g230(.Y(out_0[12]), .A0(in_2[9]), .A1(n_14), .B0(n_15));
  INVX1 g231(.Y(out_0[13]), .A(n_15));
  NOR2X1 g232(.Y(n_15), .A(in_2[9]), .B(n_14));
  INVX1 g233(.Y(n_14), .A(n_18));
  AOI2BB1X1 g234(.Y(out_0[2]), .A0N(in_2[2]), .A1N(in_2[1]), .B0(n_9));
  OAI21X1 g235(.Y(n_12), .A0(in_2[1]), .A1(n_6), .B0(n_8));
  AOI21X1 g236(.Y(n_11), .A0(in_2[7]), .A1(n_1), .B0(n_10));
  NOR2X1 g237(.Y(n_10), .A(in_2[7]), .B(n_1));
  AND2XL g238(.Y(n_9), .A(in_2[2]), .B(in_2[1]));
  NAND2X1 g239(.Y(n_8), .A(n_6), .B(in_2[1]));
  INVX1 g240(.Y(n_7), .A(in_2[4]));
  INVX1 g241(.Y(n_6), .A(in_2[3]));
  INVX1 g242(.Y(n_5), .A(in_2[2]));
  INVX1 g243(.Y(n_4), .A(in_2[8]));
  INVX1 g244(.Y(n_3), .A(in_2[6]));
  INVX1 g245(.Y(n_2), .A(in_2[5]));
  INVX1 g246(.Y(n_1), .A(in_2[9]));
endmodule

module csa_tree_SUB_TC_OP_3_group_11408_3(in_0, in_1, in_2, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
output  [13:0] out_0;
wire  n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, 
    n_20, n_19, n_18, n_17, n_15, n_13, n_12, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[1] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd3(.CO(n_22), .S(out_0[3]), .A(in_2[2]), .B(in_2[3]), .CI(n_9));
  ADDFX1 cdnfadd4(.CO(n_21), .S(out_0[4]), .A(in_2[4]), .B(n_12), .CI(n_22));
  ADDFX1 cdnfadd5(.CO(n_20), .S(out_0[5]), .A(n_8), .B(n_23), .CI(n_21));
  ADDFX1 cdnfadd6(.CO(n_19), .S(out_0[6]), .A(n_29), .B(n_24), .CI(n_20));
  ADDFX1 cdnfadd7(.CO(n_18), .S(out_0[7]), .A(n_30), .B(n_25), .CI(n_19));
  ADDFX1 cdnfadd8(.CO(n_17), .S(out_0[8]), .A(n_31), .B(n_26), .CI(n_18));
  ADDFX1 cdnfadd9(.CO(n_28), .S(out_0[9]), .A(n_32), .B(n_10), .CI(n_17));
  ADDFX1 cdnfadd10(.CO(n_27), .S(out_0[10]), .A(n_2), .B(n_7), .CI(n_28));
  ADDFX1 cdnfadd_005_0(.CO(n_29), .S(n_23), .A(n_4), .B(in_2[5]), .CI(in_2[4]));
  ADDFX1 cdnfadd_006_0(.CO(n_30), .S(n_24), .A(n_5), .B(in_2[6]), .CI(in_2[5]));
  ADDFX1 cdnfadd_007_0(.CO(n_31), .S(n_25), .A(n_6), .B(in_2[7]), .CI(in_2[6]));
  ADDFX1 cdnfadd_008_0(.CO(n_32), .S(n_26), .A(n_1), .B(in_2[8]), .CI(in_2[7]));
  AOI21X1 g294(.Y(out_0[11]), .A0(in_2[8]), .A1(n_13), .B0(n_15));
  INVX1 g295(.Y(n_15), .A(out_0[13]));
  OR2X1 g296(.Y(out_0[13]), .A(in_2[8]), .B(n_13));
  INVX1 g297(.Y(n_13), .A(n_27));
  OAI21X1 g298(.Y(n_12), .A0(in_2[1]), .A1(n_5), .B0(n_8));
  AOI2BB1X1 g299(.Y(out_0[2]), .A0N(in_2[2]), .A1N(in_2[1]), .B0(n_9));
  AOI21X1 g300(.Y(n_10), .A0(in_2[6]), .A1(n_3), .B0(n_7));
  AND2XL g301(.Y(n_9), .A(in_2[2]), .B(in_2[1]));
  NAND2X1 g302(.Y(n_8), .A(n_5), .B(in_2[1]));
  NOR2X1 g303(.Y(n_7), .A(in_2[6]), .B(n_3));
  INVX1 g304(.Y(n_6), .A(in_2[4]));
  INVX1 g305(.Y(n_5), .A(in_2[3]));
  INVX1 g306(.Y(n_4), .A(in_2[2]));
  INVX1 g307(.Y(n_3), .A(in_2[8]));
  INVX1 g308(.Y(n_2), .A(in_2[7]));
  INVX1 g309(.Y(n_1), .A(in_2[5]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_3(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g507(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g508(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g509(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g510(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g511(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g512(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g513(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g514(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g515(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g516(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1XL g517(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g518(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g519(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g520(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g521(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g522(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g523(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g524(.Y(n_11), .A(in_3[4]), .B(in_3[0]));
  NOR2X1 g525(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g526(.Y(n_9), .A(in_3[4]), .B(n_2));
  NAND2X1 g527(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2X1 g528(.Y(n_7), .A(in_3[0]), .B(in_3[1]));
  INVX1 g529(.Y(n_6), .A(in_3[2]));
  INVX1 g530(.Y(n_5), .A(in_3[6]));
  INVX1 g531(.Y(n_4), .A(in_3[3]));
  INVX1 g532(.Y(n_3), .A(in_3[7]));
  INVX1 g533(.Y(n_2), .A(in_3[5]));
  INVX1 g534(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_4(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g507(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g508(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g509(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g510(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g511(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g512(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g513(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g514(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g515(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g516(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1XL g517(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g518(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g519(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g520(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g521(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g522(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g523(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g524(.Y(n_11), .A(in_3[4]), .B(in_3[0]));
  NOR2X1 g525(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g526(.Y(n_9), .A(in_3[4]), .B(n_2));
  NAND2X1 g527(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2X1 g528(.Y(n_7), .A(in_3[0]), .B(in_3[1]));
  INVX1 g529(.Y(n_6), .A(in_3[2]));
  INVX1 g530(.Y(n_5), .A(in_3[6]));
  INVX1 g531(.Y(n_4), .A(in_3[3]));
  INVX1 g532(.Y(n_3), .A(in_3[7]));
  INVX1 g533(.Y(n_2), .A(in_3[5]));
  INVX1 g534(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_5(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g516(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g517(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g518(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g519(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g520(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g521(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g522(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g523(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g524(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g525(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1X1 g526(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g527(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g528(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g529(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g530(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g531(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g532(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g533(.Y(n_11), .A(in_3[4]), .B(in_3[0]));
  NOR2X1 g534(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g535(.Y(n_9), .A(in_3[4]), .B(n_2));
  NAND2X1 g536(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2X1 g537(.Y(n_7), .A(in_3[1]), .B(in_3[0]));
  INVX1 g538(.Y(n_6), .A(in_3[2]));
  INVX1 g539(.Y(n_5), .A(in_3[6]));
  INVX1 g540(.Y(n_4), .A(in_3[3]));
  INVX1 g541(.Y(n_3), .A(in_3[7]));
  INVX1 g542(.Y(n_2), .A(in_3[5]));
  INVX1 g543(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_6(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_39, n_36, n_34, n_32, 
    n_30, n_28, n_26, n_24, n_22, n_20, n_19, n_17, n_16, n_15, n_14, n_13, 
    n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_46), .S(n_42), .A(n_9), .B(in_3[2]), .CI(n_8));
  ADDFX1 cdnfadd_006_0(.CO(n_47), .S(n_43), .A(n_7), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_48), .S(n_44), .A(n_4), .B(in_3[4]), .CI(n_3));
  ADDFX1 cdnfadd_008_0(.CO(n_49), .S(n_45), .A(n_2), .B(in_3[5]), .CI(n_6));
  NAND3BXL g510(.Y(out_0[13]), .AN(in_3[8]), .B(n_3), .C(n_39));
  XOR2XL g511(.Y(out_0[12]), .A(n_13), .B(n_39));
  ADDFX1 g512(.CO(n_39), .S(out_0[11]), .A(n_11), .B(n_19), .CI(n_36));
  ADDFX1 g513(.CO(n_36), .S(out_0[10]), .A(n_14), .B(n_15), .CI(n_34));
  ADDFX1 g514(.CO(n_34), .S(out_0[9]), .A(n_17), .B(n_49), .CI(n_32));
  ADDFX1 g515(.CO(n_32), .S(out_0[8]), .A(n_48), .B(n_45), .CI(n_30));
  ADDFX1 g516(.CO(n_30), .S(out_0[7]), .A(n_47), .B(n_44), .CI(n_28));
  ADDFX1 g517(.CO(n_28), .S(out_0[6]), .A(n_46), .B(n_43), .CI(n_26));
  ADDFX1 g518(.CO(n_26), .S(out_0[5]), .A(n_12), .B(n_42), .CI(n_24));
  ADDFX1 g519(.CO(n_24), .S(out_0[4]), .A(in_3[1]), .B(n_16), .CI(n_22));
  ADDFX1 g520(.CO(n_22), .S(out_0[3]), .A(n_4), .B(n_1), .CI(n_20));
  AOI2BB1X1 g521(.Y(out_0[2]), .A0N(n_7), .A1N(n_10), .B0(n_20));
  AND2XL g522(.Y(n_20), .A(n_7), .B(n_10));
  AOI21X1 g523(.Y(n_19), .A0(in_3[7]), .A1(in_3[8]), .B0(n_13));
  AOI21X1 g524(.Y(out_0[1]), .A0(in_3[1]), .A1(n_1), .B0(n_10));
  OAI2BB1X1 g525(.Y(n_17), .A0N(in_3[6]), .A1N(n_8), .B0(n_14));
  OAI21X1 g526(.Y(n_16), .A0(in_3[4]), .A1(n_1), .B0(n_12));
  OAI2BB1X1 g527(.Y(n_15), .A0N(in_3[7]), .A1N(n_5), .B0(n_11));
  NAND2X1 g528(.Y(n_14), .A(in_3[5]), .B(n_5));
  NOR2X1 g529(.Y(n_13), .A(in_3[7]), .B(in_3[8]));
  NAND2X1 g530(.Y(n_12), .A(in_3[4]), .B(n_1));
  NAND2X1 g531(.Y(n_11), .A(in_3[6]), .B(n_3));
  NOR2X1 g532(.Y(n_10), .A(in_3[1]), .B(n_1));
  INVX1 g533(.Y(n_9), .A(in_3[1]));
  INVX1 g534(.Y(n_8), .A(in_3[5]));
  INVX1 g535(.Y(n_7), .A(in_3[2]));
  INVX1 g536(.Y(n_6), .A(in_3[8]));
  INVX1 g537(.Y(n_5), .A(in_3[6]));
  INVX1 g538(.Y(n_4), .A(in_3[3]));
  INVX1 g539(.Y(n_3), .A(in_3[7]));
  INVX1 g540(.Y(n_2), .A(in_3[4]));
  INVX1 drc_bufs541(.Y(n_1), .A(n_0));
  INVX1 drc_bufs542(.Y(n_0), .A(in_3[0]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_7(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_34, n_32, n_30, 
    n_28, n_26, n_24, n_22, n_20, n_18, n_17, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_44), .S(n_40), .A(n_7), .B(in_3[2]), .CI(n_6));
  ADDFX1 cdnfadd_006_0(.CO(n_45), .S(n_41), .A(n_5), .B(in_3[3]), .CI(n_3));
  ADDFX1 cdnfadd_007_0(.CO(n_46), .S(n_42), .A(n_2), .B(in_3[4]), .CI(n_1));
  ADDFX1 cdnfadd_008_0(.CO(n_47), .S(n_43), .A(n_0), .B(in_3[5]), .CI(n_4));
  NAND3BXL g510(.Y(out_0[13]), .AN(in_3[8]), .B(n_1), .C(n_37));
  XOR2XL g511(.Y(out_0[12]), .A(n_11), .B(n_37));
  ADDFX1 g512(.CO(n_37), .S(out_0[11]), .A(n_9), .B(n_17), .CI(n_34));
  ADDFX1 g513(.CO(n_34), .S(out_0[10]), .A(n_12), .B(n_13), .CI(n_32));
  ADDFX1 g514(.CO(n_32), .S(out_0[9]), .A(n_15), .B(n_47), .CI(n_30));
  ADDFX1 g515(.CO(n_30), .S(out_0[8]), .A(n_46), .B(n_43), .CI(n_28));
  ADDFX1 g516(.CO(n_28), .S(out_0[7]), .A(n_45), .B(n_42), .CI(n_26));
  ADDFX1 g517(.CO(n_26), .S(out_0[6]), .A(n_44), .B(n_41), .CI(n_24));
  ADDFX1 g518(.CO(n_24), .S(out_0[5]), .A(n_10), .B(n_40), .CI(n_22));
  ADDFX1 g519(.CO(n_22), .S(out_0[4]), .A(in_3[1]), .B(n_14), .CI(n_20));
  ADDFX1 g520(.CO(n_20), .S(out_0[3]), .A(n_2), .B(in_3[0]), .CI(n_18));
  AOI2BB1X1 g521(.Y(out_0[2]), .A0N(n_5), .A1N(n_8), .B0(n_18));
  AND2XL g522(.Y(n_18), .A(n_5), .B(n_8));
  AOI21X1 g523(.Y(n_17), .A0(in_3[7]), .A1(in_3[8]), .B0(n_11));
  AOI21X1 g524(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_8));
  OAI2BB1X1 g525(.Y(n_15), .A0N(in_3[6]), .A1N(n_6), .B0(n_12));
  OAI21X1 g526(.Y(n_14), .A0(in_3[4]), .A1(in_3[0]), .B0(n_10));
  OAI2BB1X1 g527(.Y(n_13), .A0N(in_3[7]), .A1N(n_3), .B0(n_9));
  NAND2X1 g528(.Y(n_12), .A(in_3[5]), .B(n_3));
  NOR2XL g529(.Y(n_11), .A(in_3[8]), .B(in_3[7]));
  NAND2X1 g530(.Y(n_10), .A(in_3[4]), .B(in_3[0]));
  NAND2X1 g531(.Y(n_9), .A(in_3[6]), .B(n_1));
  NOR2XL g532(.Y(n_8), .A(in_3[1]), .B(in_3[0]));
  INVX1 g533(.Y(n_7), .A(in_3[1]));
  INVX1 g534(.Y(n_6), .A(in_3[5]));
  INVX1 g535(.Y(n_5), .A(in_3[2]));
  INVX1 g536(.Y(n_4), .A(in_3[8]));
  INVX1 g537(.Y(n_3), .A(in_3[6]));
  INVX1 g538(.Y(n_2), .A(in_3[3]));
  INVX1 g539(.Y(n_1), .A(in_3[7]));
  INVX1 g540(.Y(n_0), .A(in_3[4]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_8(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g507(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g508(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g509(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g510(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g511(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g512(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g513(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g514(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g515(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g516(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1X1 g517(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g518(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g519(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g520(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g521(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g522(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g523(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g524(.Y(n_11), .A(in_3[0]), .B(in_3[4]));
  NOR2X1 g525(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g526(.Y(n_9), .A(n_2), .B(in_3[4]));
  NAND2X1 g527(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2X1 g528(.Y(n_7), .A(in_3[0]), .B(in_3[1]));
  INVX1 g529(.Y(n_6), .A(in_3[2]));
  INVX1 g530(.Y(n_5), .A(in_3[6]));
  INVX1 g531(.Y(n_4), .A(in_3[3]));
  INVX1 g532(.Y(n_3), .A(in_3[7]));
  INVX1 g533(.Y(n_2), .A(in_3[5]));
  INVX1 g534(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_1752_3(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [12:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_37, n_35, 
    n_33, n_31, n_29, n_27, n_25, n_23, n_21, n_19, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [12:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_004_1(.CO(n_56), .S(n_48), .A(in_3[3]), .B(n_6), .CI(n_11));
  ADDFX1 cdnfadd_005_0(.CO(n_47), .S(n_46), .A(n_1), .B(in_3[5]), .CI(in_3[4]));
  ADDFX1 cdnfadd_005_1(.CO(n_57), .S(n_49), .A(in_3[2]), .B(n_7), .CI(n_46));
  ADDFX1 cdnfadd_006_0(.CO(n_45), .S(n_44), .A(n_2), .B(in_3[6]), .CI(in_3[5]));
  ADDFX1 cdnfadd_006_1(.CO(n_58), .S(n_50), .A(in_3[3]), .B(n_47), .CI(n_44));
  ADDFX1 cdnfadd_007_0(.CO(n_43), .S(n_42), .A(n_3), .B(in_3[7]), .CI(in_3[6]));
  ADDFX1 cdnfadd_007_1(.CO(n_59), .S(n_51), .A(in_3[4]), .B(n_45), .CI(n_42));
  ADDFX1 cdnfadd_008_0(.CO(n_41), .S(n_40), .A(n_4), .B(in_3[8]), .CI(in_3[7]));
  ADDFX1 cdnfadd_008_1(.CO(n_53), .S(n_52), .A(in_3[5]), .B(n_43), .CI(n_40));
  ADDFX1 cdnfadd_009_0(.CO(n_54), .S(n_60), .A(in_3[8]), .B(n_13), .CI(n_41));
  ADDFX1 cdnfadd_010_0(.CO(n_55), .S(n_61), .A(n_5), .B(in_3[7]), .CI(n_10));
  NAND2X1 g473(.Y(out_0[13]), .A(n_9), .B(n_37));
  ADDFX1 g474(.CO(n_37), .S(out_0[11]), .A(n_17), .B(n_55), .CI(n_35));
  ADDFX1 g475(.CO(n_35), .S(out_0[10]), .A(n_54), .B(n_61), .CI(n_33));
  ADDFX1 g476(.CO(n_33), .S(out_0[9]), .A(n_60), .B(n_53), .CI(n_31));
  ADDFX1 g477(.CO(n_31), .S(out_0[8]), .A(n_59), .B(n_52), .CI(n_29));
  ADDFX1 g478(.CO(n_29), .S(out_0[7]), .A(n_58), .B(n_51), .CI(n_27));
  ADDFX1 g479(.CO(n_27), .S(out_0[6]), .A(n_57), .B(n_50), .CI(n_25));
  ADDFX1 g480(.CO(n_25), .S(out_0[5]), .A(n_56), .B(n_23), .CI(n_49));
  ADDFX1 g481(.CO(n_23), .S(out_0[4]), .A(n_16), .B(n_21), .CI(n_48));
  ADDFX1 g482(.CO(n_21), .S(out_0[3]), .A(in_3[2]), .B(n_14), .CI(n_19));
  XOR2XL g483(.Y(out_0[2]), .A(n_8), .B(n_15));
  NAND2XL g484(.Y(n_19), .A(n_12), .B(n_8));
  OA21X1 g485(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_8));
  OAI21X1 g486(.Y(n_17), .A0(in_3[8]), .A1(in_3[7]), .B0(n_9));
  OAI2BB1X1 g487(.Y(n_16), .A0N(in_3[4]), .A1N(in_3[1]), .B0(n_7));
  OAI2BB1X1 g488(.Y(n_15), .A0N(n_1), .A1N(n_2), .B0(n_12));
  AOI21X1 g489(.Y(n_14), .A0(n_3), .A1(n_6), .B0(n_11));
  AOI21X1 g490(.Y(n_13), .A0(in_3[5]), .A1(n_5), .B0(n_10));
  NAND2X1 g491(.Y(n_12), .A(in_3[1]), .B(in_3[2]));
  NOR2X1 g492(.Y(n_11), .A(n_3), .B(n_6));
  NOR2X1 g493(.Y(n_10), .A(in_3[5]), .B(n_5));
  NAND2X1 g494(.Y(n_9), .A(in_3[7]), .B(in_3[8]));
  NAND2X1 g495(.Y(n_8), .A(in_3[1]), .B(in_3[0]));
  NAND2X1 g496(.Y(n_7), .A(n_4), .B(n_1));
  INVX1 g497(.Y(n_6), .A(in_3[0]));
  INVX1 g498(.Y(n_5), .A(in_3[6]));
  INVX1 g499(.Y(n_4), .A(in_3[4]));
  INVX1 g500(.Y(n_3), .A(in_3[3]));
  INVX1 g501(.Y(n_2), .A(in_3[2]));
  INVX1 g502(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_9(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g507(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g508(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g509(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g510(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g511(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g512(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g513(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g514(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g515(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g516(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1X1 g517(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g518(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g519(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g520(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g521(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g522(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g523(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g524(.Y(n_11), .A(in_3[4]), .B(in_3[0]));
  NOR2X1 g525(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g526(.Y(n_9), .A(in_3[4]), .B(n_2));
  NAND2X1 g527(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2XL g528(.Y(n_7), .A(in_3[1]), .B(in_3[0]));
  INVX1 g529(.Y(n_6), .A(in_3[2]));
  INVX1 g530(.Y(n_5), .A(in_3[6]));
  INVX1 g531(.Y(n_4), .A(in_3[3]));
  INVX1 g532(.Y(n_3), .A(in_3[7]));
  INVX1 g533(.Y(n_2), .A(in_3[5]));
  INVX1 g534(.Y(n_1), .A(in_3[1]));
endmodule

module csa_tree_SUB_TC_OP_4_group_54_10(in_0, in_1, in_2, in_3, out_0);
input   [13:0] in_0;
input   [11:0] in_1;
input   [10:0] in_2;
input   [9:0] in_3;
output  [13:0] out_0;
wire  n_42, n_41, n_40, n_39, n_38, n_37, n_34, n_31, n_29, n_27, n_25, n_23, 
    n_21, n_19, n_17, n_16, n_15, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
    n_5, n_4, n_3, n_2, n_1;
wire   [13:0] out_0;
wire   [9:0] in_3;
wire   [10:0] in_2;
wire   [11:0] in_1;
wire   [13:0] in_0;
  assign out_0[12] = 1'b0;
  assign out_0[0] = 1'b0;
  ADDFX1 cdnfadd_005_0(.CO(n_40), .S(n_37), .A(n_1), .B(in_3[2]), .CI(n_2));
  ADDFX1 cdnfadd_006_0(.CO(n_41), .S(n_38), .A(n_6), .B(in_3[3]), .CI(n_5));
  ADDFX1 cdnfadd_007_0(.CO(n_42), .S(n_39), .A(n_4), .B(in_3[4]), .CI(n_3));
  XOR2XL g528(.Y(out_0[11]), .A(n_10), .B(n_34));
  NAND2X1 g529(.Y(out_0[13]), .A(n_10), .B(n_34));
  ADDFX1 g530(.CO(n_34), .S(out_0[10]), .A(n_8), .B(n_16), .CI(n_31));
  ADDFX1 g531(.CO(n_31), .S(out_0[9]), .A(n_9), .B(n_12), .CI(n_29));
  ADDFX1 g532(.CO(n_29), .S(out_0[8]), .A(n_13), .B(n_42), .CI(n_27));
  ADDFX1 g533(.CO(n_27), .S(out_0[7]), .A(n_41), .B(n_39), .CI(n_25));
  ADDFX1 g534(.CO(n_25), .S(out_0[6]), .A(n_40), .B(n_38), .CI(n_23));
  ADDFX1 g535(.CO(n_23), .S(out_0[5]), .A(n_11), .B(n_37), .CI(n_21));
  ADDFX1 g536(.CO(n_21), .S(out_0[4]), .A(in_3[1]), .B(n_15), .CI(n_19));
  ADDFX1 g537(.CO(n_19), .S(out_0[3]), .A(n_4), .B(in_3[0]), .CI(n_17));
  AOI2BB1X1 g538(.Y(out_0[2]), .A0N(n_6), .A1N(n_7), .B0(n_17));
  AND2XL g539(.Y(n_17), .A(n_6), .B(n_7));
  AOI21X1 g540(.Y(n_16), .A0(in_3[6]), .A1(in_3[7]), .B0(n_10));
  OAI21X1 g541(.Y(n_15), .A0(in_3[4]), .A1(in_3[0]), .B0(n_11));
  AOI21X1 g542(.Y(out_0[1]), .A0(in_3[1]), .A1(in_3[0]), .B0(n_7));
  OAI21X1 g543(.Y(n_13), .A0(in_3[4]), .A1(n_2), .B0(n_9));
  OAI2BB1X1 g544(.Y(n_12), .A0N(in_3[6]), .A1N(n_2), .B0(n_8));
  NAND2X1 g545(.Y(n_11), .A(in_3[0]), .B(in_3[4]));
  NOR2X1 g546(.Y(n_10), .A(in_3[6]), .B(in_3[7]));
  NAND2X1 g547(.Y(n_9), .A(n_2), .B(in_3[4]));
  NAND2X1 g548(.Y(n_8), .A(in_3[5]), .B(n_5));
  NOR2XL g549(.Y(n_7), .A(in_3[1]), .B(in_3[0]));
  INVX1 g550(.Y(n_6), .A(in_3[2]));
  INVX1 g551(.Y(n_5), .A(in_3[6]));
  INVX1 g552(.Y(n_4), .A(in_3[3]));
  INVX1 g553(.Y(n_3), .A(in_3[7]));
  INVX1 g554(.Y(n_2), .A(in_3[5]));
  INVX1 g555(.Y(n_1), .A(in_3[1]));
endmodule

module mytop(in, clk, rst_n, updown, out_activehigh, done);
input  clk, rst_n, updown;
output done;
input   [127:0] in;
output  [0:9] out_activehigh;
wire  n_568, n_567, n_566, n_565, n_564, n_563, n_562, n_561, n_560, n_559, 
    n_558, n_557, n_556, n_555, n_554, n_553, n_552, n_551, n_550, n_549, 
    n_548, n_547, n_546, n_545, n_544, n_543, n_542, n_541, n_540, n_539, 
    n_538, n_537, n_536, n_535, n_534, n_533, n_532, n_531, n_530, n_529, 
    n_528, n_527, n_526, n_525, n_524, n_523, n_522, n_521, n_520, n_519, 
    n_518, n_517, n_516, n_515, n_514, n_513, n_512, n_511, n_510, n_509, 
    n_508, n_507, n_506, n_505, n_504, n_503, n_502, n_501, n_500, n_499, 
    n_498, n_497, n_496, n_495, n_494, n_493, n_492, n_491, n_490, n_489, 
    n_488, n_487, n_486, n_485, n_484, n_483, n_482, n_481, n_480, n_479, 
    n_478, n_477, n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, 
    n_468, n_467, n_466, n_465, n_464, n_463, n_462, n_461, n_460, n_459, 
    n_458, n_457, n_456, n_455, n_454, n_453, n_452, n_451, n_450, n_449, 
    n_448, n_447, n_446, n_445, n_444, n_443, n_442, n_441, n_440, n_439, 
    n_438, n_437, n_436, n_435, n_434, n_433, n_432, n_431, n_430, n_429, 
    n_428, n_427, n_426, n_425, n_424, n_423, n_422, n_421, n_420, n_419, 
    n_418, n_417, n_416, n_415, n_414, n_413, n_412, n_411, n_410, n_409, 
    n_408, n_407, n_406, n_405, n_404, n_403, n_402, n_401, n_400, n_399, 
    n_398, n_397, n_396, n_395, n_394, n_393, n_392, n_391, n_390, n_389, 
    n_388, n_387, n_386, n_385, n_384, n_383, n_382, n_381, n_380, n_379, 
    n_378, n_377, n_376, n_375, n_374, n_373, n_372, n_371, n_370, n_369, 
    n_368, n_367, n_366, n_365, n_364, n_363, n_362, n_361, n_360, n_359, 
    n_358, n_357, n_356, n_355, n_354, n_353, n_352, n_351, n_350, n_349, 
    n_348, n_347, n_346, n_345, n_344, n_343, n_342, n_341, n_340, n_339, 
    n_338, n_337, n_336, n_335, n_334, n_333, n_332, n_331, n_330, n_329, 
    n_328, n_327, n_326, n_325, n_324, n_323, n_322, n_321, n_320, n_319, 
    n_318, n_317, n_316, n_315, n_314, n_313, n_312, n_311, n_310, n_309, 
    n_308, n_307, n_306, n_305, n_304, n_303, n_302, n_301, n_300, n_299, 
    n_298, n_297, n_296, n_295, n_294, n_293, n_292, n_291, n_290, n_289, 
    n_288, n_287, n_286, n_285, n_284, n_283, n_282, n_281, n_280, n_279, 
    n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, 
    n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, 
    n_258, n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, n_249, 
    n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
    n_238, n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, 
    n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, 
    n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, 
    n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, 
    n_198, n_197, n_196, n_195, n_194, n_193, n_192, n_191, n_190, n_189, 
    n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, 
    n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, 
    n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, 
    n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, 
    n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, 
    n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, 
    n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
    n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
    n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, 
    n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
    n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, 
    n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
    n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, 
    \instanceL2_prod_terms[7][9][12] , \instanceL2_prod_terms[7][9][11] , 
    \instanceL2_prod_terms[7][9][10] , \instanceL2_prod_terms[7][9][9] , 
    \instanceL2_prod_terms[7][9][8] , \instanceL2_prod_terms[7][9][7] , 
    \instanceL2_prod_terms[7][9][6] , \instanceL2_prod_terms[7][9][5] , 
    \instanceL2_prod_terms[7][9][4] , \instanceL2_prod_terms[7][9][3] , 
    \instanceL2_prod_terms[2][11][11] , \instanceL2_prod_terms[2][11][10] , 
    \instanceL2_prod_terms[2][11][9] , \instanceL2_prod_terms[2][11][8] , 
    \instanceL2_prod_terms[2][11][7] , \instanceL2_prod_terms[2][11][6] , 
    \instanceL2_prod_terms[2][11][5] , \instanceL2_prod_terms[2][11][4] , 
    \instanceL2_prod_terms[2][11][2] , \instanceL2_prod_terms[2][8][11] , 
    \instanceL2_prod_terms[2][8][10] , \instanceL2_prod_terms[2][8][9] , 
    \instanceL2_prod_terms[2][8][8] , \instanceL2_prod_terms[2][8][7] , 
    \instanceL2_prod_terms[2][8][6] , \instanceL2_prod_terms[2][8][5] , 
    \instanceL2_prod_terms[2][8][4] , \instanceL2_prod_terms[2][8][3] , 
    \instanceL2_prod_terms[2][8][2] , \instanceL2_prod_terms[1][10][10] , 
    \instanceL2_prod_terms[1][10][9] , \instanceL2_prod_terms[1][10][8] , 
    \instanceL2_prod_terms[1][10][7] , \instanceL2_prod_terms[1][10][6] , 
    \instanceL2_prod_terms[1][10][5] , \instanceL2_prod_terms[1][10][4] , 
    \instanceL2_prod_terms[1][10][3] , \instanceL2_prod_terms[1][10][2] , 
    \instanceL2_prod_terms[1][8][13] , \instanceL2_prod_terms[1][8][9] , 
    \instanceL2_prod_terms[1][8][8] , \instanceL2_prod_terms[1][8][7] , 
    \instanceL2_prod_terms[1][8][6] , \instanceL2_prod_terms[1][8][5] , 
    \instanceL2_prod_terms[1][8][4] , \instanceL2_prod_terms[1][8][3] , 
    \instanceL2_prod_terms[1][8][2] , \instanceL2_prod_terms[1][2][12] , 
    \instanceL2_prod_terms[1][2][11] , \instanceL2_prod_terms[1][2][10] , 
    \instanceL2_prod_terms[1][2][9] , \instanceL2_prod_terms[1][2][8] , 
    \instanceL2_prod_terms[1][2][7] , \instanceL2_prod_terms[1][2][6] , 
    \instanceL2_prod_terms[1][2][5] , \instanceL2_prod_terms[1][2][4] , 
    \instanceL2_prod_terms[1][2][3] , \instanceL2_prod_terms[1][1][9] , 
    \instanceL2_prod_terms[1][1][8] , \instanceL2_prod_terms[1][1][7] , 
    \instanceL2_prod_terms[1][1][6] , \instanceL2_prod_terms[1][1][5] , 
    \instanceL2_prod_terms[1][1][4] , \instanceL2_prod_terms[1][1][3] , 
    \instanceL2_prod_terms[1][1][2] , \instanceL2_prod_terms[0][19][13] , 
    \instanceL2_prod_terms[0][19][10] , \instanceL2_prod_terms[0][19][9] , 
    \instanceL2_prod_terms[0][19][8] , \instanceL2_prod_terms[0][19][7] , 
    \instanceL2_prod_terms[0][19][6] , \instanceL2_prod_terms[0][19][5] , 
    \instanceL2_prod_terms[0][19][4] , \instanceL2_prod_terms[0][19][3] , 
    \instanceL2_prod_terms[0][19][2] , \instanceL2_prod_terms[0][19][1] , 
    \instanceL2_prod_terms[0][17][10] , \instanceL2_prod_terms[0][17][9] , 
    \instanceL2_prod_terms[0][17][8] , \instanceL2_prod_terms[0][17][7] , 
    \instanceL2_prod_terms[0][17][6] , \instanceL2_prod_terms[0][17][5] , 
    \instanceL2_prod_terms[0][17][4] , \instanceL2_prod_terms[0][17][3] , 
    \instanceL2_prod_terms[0][17][2] , \instanceL2_prod_terms[0][16][13] , 
    \instanceL2_prod_terms[0][16][7] , \instanceL2_prod_terms[0][16][6] , 
    \instanceL2_prod_terms[0][16][5] , \instanceL2_prod_terms[0][16][4] , 
    \instanceL2_prod_terms[0][16][3] , \instanceL2_prod_terms[0][16][2] , 
    \instanceL2_prod_terms[0][16][1] , \instanceL2_prod_terms[0][14][9] , 
    \instanceL2_prod_terms[0][14][8] , \instanceL2_prod_terms[0][14][7] , 
    \instanceL2_prod_terms[0][14][6] , \instanceL2_prod_terms[0][14][5] , 
    \instanceL2_prod_terms[0][14][4] , \instanceL2_prod_terms[0][14][3] , 
    \instanceL2_prod_terms[0][14][2] , \instanceL2_prod_terms[0][11][13] , 
    \instanceL2_prod_terms[0][11][7] , \instanceL2_prod_terms[0][11][6] , 
    \instanceL2_prod_terms[0][11][5] , \instanceL2_prod_terms[0][11][4] , 
    \instanceL2_prod_terms[0][11][3] , \instanceL2_prod_terms[0][11][2] , 
    \instanceL2_prod_terms[0][11][1] , \instanceL2_prod_terms[0][10][13] , 
    \instanceL2_prod_terms[0][10][8] , \instanceL2_prod_terms[0][10][7] , 
    \instanceL2_prod_terms[0][10][6] , \instanceL2_prod_terms[0][10][5] , 
    \instanceL2_prod_terms[0][10][4] , \instanceL2_prod_terms[0][10][3] , 
    \instanceL2_prod_terms[0][10][2] , \instanceL2_prod_terms[0][9][13] , 
    \instanceL2_prod_terms[0][9][12] , \instanceL2_prod_terms[0][9][11] , 
    \instanceL2_prod_terms[0][9][10] , \instanceL2_prod_terms[0][9][9] , 
    \instanceL2_prod_terms[0][9][8] , \instanceL2_prod_terms[0][9][7] , 
    \instanceL2_prod_terms[0][9][6] , \instanceL2_prod_terms[0][9][5] , 
    \instanceL2_prod_terms[0][9][4] , \instanceL2_prod_terms[0][9][3] , 
    \instanceL2_prod_terms[0][9][2] , \instanceL2_prod_terms[0][9][1] , 
    \instanceL2_prod_terms[0][5][9] , \instanceL2_prod_terms[0][5][8] , 
    \instanceL2_prod_terms[0][5][7] , \instanceL2_prod_terms[0][5][6] , 
    \instanceL2_prod_terms[0][5][5] , \instanceL2_prod_terms[0][5][4] , 
    \instanceL2_prod_terms[0][5][3] , \instanceL2_prod_terms[0][4][10] , 
    \instanceL2_prod_terms[0][4][9] , \instanceL2_prod_terms[0][4][8] , 
    \instanceL2_prod_terms[0][4][7] , \instanceL2_prod_terms[0][4][6] , 
    \instanceL2_prod_terms[0][4][5] , \instanceL2_prod_terms[0][4][4] , 
    \instanceL2_prod_terms[0][3][9] , \instanceL2_prod_terms[0][3][8] , 
    \instanceL2_prod_terms[0][3][7] , \instanceL2_prod_terms[0][3][6] , 
    \instanceL2_prod_terms[0][3][5] , \instanceL2_prod_terms[0][3][4] , 
    \instanceL2_prod_terms[0][3][3] , \instanceL2_prod_terms[0][3][2] , 
    \instanceL2_prod_terms[0][2][10] , \instanceL2_prod_terms[0][2][9] , 
    \instanceL2_prod_terms[0][2][8] , \instanceL2_prod_terms[0][2][7] , 
    \instanceL2_prod_terms[0][2][6] , \instanceL2_prod_terms[0][2][5] , 
    \instanceL2_prod_terms[0][2][4] , \instanceL2_prod_terms[0][2][3] , 
    \instanceL2_prod_terms[0][1][8] , \instanceL2_prod_terms[0][1][4] , 
    \instanceL2_prod_terms[0][0][13] , \instanceL2_prod_terms[0][0][8] , 
    \instanceL2_prod_terms[0][0][7] , \instanceL2_prod_terms[0][0][6] , 
    \instanceL2_prod_terms[0][0][5] , \instanceL2_prod_terms[0][0][4] , 
    \instanceL2_prod_terms[0][0][3] , \instanceL2_prod_terms[0][0][2] , 
    instanceL2_n_12646, instanceL2_n_12645, instanceL2_n_12644, 
    instanceL2_n_12643, instanceL2_n_12642, instanceL2_n_12641, 
    instanceL2_n_12640, instanceL2_n_12639, instanceL2_n_12638, 
    instanceL2_n_12637, instanceL2_n_12636, instanceL2_n_12635, 
    instanceL2_n_12634, instanceL2_n_12633, instanceL2_n_12632, 
    instanceL2_n_12631, instanceL2_n_12630, instanceL2_n_12629, 
    instanceL2_n_12628, instanceL2_n_12627, instanceL2_n_12626, 
    instanceL2_n_12625, instanceL2_n_12624, instanceL2_n_12623, 
    instanceL2_n_12622, instanceL2_n_12621, instanceL2_n_12620, 
    instanceL2_n_12619, instanceL2_n_12618, instanceL2_n_12617, 
    instanceL2_n_12616, instanceL2_n_12615, instanceL2_n_12614, 
    instanceL2_n_12613, instanceL2_n_12612, instanceL2_n_12611, 
    instanceL2_n_12610, instanceL2_n_12609, instanceL2_n_12608, 
    instanceL2_n_12607, instanceL2_n_12606, instanceL2_n_12605, 
    instanceL2_n_12604, instanceL2_n_12603, instanceL2_n_12602, 
    instanceL2_n_12601, instanceL2_n_12600, instanceL2_n_12599, 
    instanceL2_n_12598, instanceL2_n_12597, instanceL2_n_12596, 
    instanceL2_n_12595, instanceL2_n_12594, instanceL2_n_12593, 
    instanceL2_n_12592, instanceL2_n_12591, instanceL2_n_12590, 
    instanceL2_n_12589, instanceL2_n_12588, instanceL2_n_12587, 
    instanceL2_n_12586, instanceL2_n_12585, instanceL2_n_12584, 
    instanceL2_n_12583, instanceL2_n_12582, instanceL2_n_12581, 
    instanceL2_n_12580, instanceL2_n_12579, instanceL2_n_12578, 
    instanceL2_n_12577, instanceL2_n_12576, instanceL2_n_12575, 
    instanceL2_n_12574, instanceL2_n_12573, instanceL2_n_12572, 
    instanceL2_n_12571, instanceL2_n_12570, instanceL2_n_12569, 
    instanceL2_n_12568, instanceL2_n_12567, instanceL2_n_12566, 
    instanceL2_n_12565, instanceL2_n_12564, instanceL2_n_12563, 
    instanceL2_n_12562, instanceL2_n_12561, instanceL2_n_12560, 
    instanceL2_n_12559, instanceL2_n_12558, instanceL2_n_12557, 
    instanceL2_n_12556, instanceL2_n_12555, instanceL2_n_12554, 
    instanceL2_n_12553, instanceL2_n_12552, instanceL2_n_12551, 
    instanceL2_n_12550, instanceL2_n_12549, instanceL2_n_12548, 
    instanceL2_n_12547, instanceL2_n_12546, instanceL2_n_12545, 
    instanceL2_n_12544, instanceL2_n_12543, instanceL2_n_12542, 
    instanceL2_n_12541, instanceL2_n_12540, instanceL2_n_12539, 
    instanceL2_n_12538, instanceL2_n_12537, instanceL2_n_12536, 
    instanceL2_n_12535, instanceL2_n_12534, instanceL2_n_12533, 
    instanceL2_n_12532, instanceL2_n_12531, instanceL2_n_12530, 
    instanceL2_n_12529, instanceL2_n_12528, instanceL2_n_12527, 
    instanceL2_n_12526, instanceL2_n_12525, instanceL2_n_12524, 
    instanceL2_n_12523, instanceL2_n_12522, instanceL2_n_12521, 
    instanceL2_n_12520, instanceL2_n_12519, instanceL2_n_12518, 
    instanceL2_n_12517, instanceL2_n_12516, instanceL2_n_12515, 
    instanceL2_n_12514, instanceL2_n_12513, instanceL2_n_12512, 
    instanceL2_n_12511, instanceL2_n_12510, instanceL2_n_12509, 
    instanceL2_n_12508, instanceL2_n_12507, instanceL2_n_12506, 
    instanceL2_n_12505, instanceL2_n_12504, instanceL2_n_12503, 
    instanceL2_n_12502, instanceL2_n_12501, instanceL2_n_12500, 
    instanceL2_n_12499, instanceL2_n_12498, instanceL2_n_12497, 
    instanceL2_n_12496, instanceL2_n_12495, instanceL2_n_12494, 
    instanceL2_n_12493, instanceL2_n_12492, instanceL2_n_12491, 
    instanceL2_n_12490, instanceL2_n_12489, instanceL2_n_12488, 
    instanceL2_n_12487, instanceL2_n_12486, instanceL2_n_12485, 
    instanceL2_n_12484, instanceL2_n_12483, instanceL2_n_12482, 
    instanceL2_n_12481, instanceL2_n_12480, instanceL2_n_12479, 
    instanceL2_n_12478, instanceL2_n_12477, instanceL2_n_12476, 
    instanceL2_n_12475, instanceL2_n_12474, instanceL2_n_12473, 
    instanceL2_n_12472, instanceL2_n_12471, instanceL2_n_12470, 
    instanceL2_n_12469, instanceL2_n_12468, instanceL2_n_12467, 
    instanceL2_n_12466, instanceL2_n_12465, instanceL2_n_12464, 
    instanceL2_n_12463, instanceL2_n_12462, instanceL2_n_12461, 
    instanceL2_n_12460, instanceL2_n_12459, instanceL2_n_12458, 
    instanceL2_n_12457, instanceL2_n_12456, instanceL2_n_12455, 
    instanceL2_n_12454, instanceL2_n_12453, instanceL2_n_12452, 
    instanceL2_n_12451, instanceL2_n_12450, instanceL2_n_12449, 
    instanceL2_n_12448, instanceL2_n_12447, instanceL2_n_12446, 
    instanceL2_n_12445, instanceL2_n_12444, instanceL2_n_12443, 
    instanceL2_n_12442, instanceL2_n_12441, instanceL2_n_12440, 
    instanceL2_n_12439, instanceL2_n_12438, instanceL2_n_12437, 
    instanceL2_n_12436, instanceL2_n_12435, instanceL2_n_12434, 
    instanceL2_n_12433, instanceL2_n_12432, instanceL2_n_12431, 
    instanceL2_n_12430, instanceL2_n_12429, instanceL2_n_12428, 
    instanceL2_n_12427, instanceL2_n_12426, instanceL2_n_12425, 
    instanceL2_n_12424, instanceL2_n_12423, instanceL2_n_12422, 
    instanceL2_n_12421, instanceL2_n_12420, instanceL2_n_12419, 
    instanceL2_n_12418, instanceL2_n_12417, instanceL2_n_12416, 
    instanceL2_n_12415, instanceL2_n_12414, instanceL2_n_12413, 
    instanceL2_n_12412, instanceL2_n_12411, instanceL2_n_12410, 
    instanceL2_n_12409, instanceL2_n_12408, instanceL2_n_12407, 
    instanceL2_n_12406, instanceL2_n_12405, instanceL2_n_12404, 
    instanceL2_n_12403, instanceL2_n_12402, instanceL2_n_12401, 
    instanceL2_n_12400, instanceL2_n_12399, instanceL2_n_12398, 
    instanceL2_n_12397, instanceL2_n_12396, instanceL2_n_12395, 
    instanceL2_n_12394, instanceL2_n_12393, instanceL2_n_12392, 
    instanceL2_n_12391, instanceL2_n_12390, instanceL2_n_12389, 
    instanceL2_n_12388, instanceL2_n_12387, instanceL2_n_12386, 
    instanceL2_n_12385, instanceL2_n_12384, instanceL2_n_12383, 
    instanceL2_n_12382, instanceL2_n_12381, instanceL2_n_12380, 
    instanceL2_n_12379, instanceL2_n_12378, instanceL2_n_12377, 
    instanceL2_n_12376, instanceL2_n_12375, instanceL2_n_12374, 
    instanceL2_n_12373, instanceL2_n_12372, instanceL2_n_12371, 
    instanceL2_n_12370, instanceL2_n_12369, instanceL2_n_12368, 
    instanceL2_n_12367, instanceL2_n_12366, instanceL2_n_12365, 
    instanceL2_n_12364, instanceL2_n_12363, instanceL2_n_12362, 
    instanceL2_n_12361, instanceL2_n_12360, instanceL2_n_12359, 
    instanceL2_n_12358, instanceL2_n_12357, instanceL2_n_12356, 
    instanceL2_n_12355, instanceL2_n_12354, instanceL2_n_12353, 
    instanceL2_n_12352, instanceL2_n_12351, instanceL2_n_12350, 
    instanceL2_n_12349, instanceL2_n_12348, instanceL2_n_12347, 
    instanceL2_n_12346, instanceL2_n_12345, instanceL2_n_12344, 
    instanceL2_n_12343, instanceL2_n_12342, instanceL2_n_12341, 
    instanceL2_n_12340, instanceL2_n_12339, instanceL2_n_12338, 
    instanceL2_n_12337, instanceL2_n_12336, instanceL2_n_12335, 
    instanceL2_n_12334, instanceL2_n_12333, instanceL2_n_12332, 
    instanceL2_n_12331, instanceL2_n_12330, instanceL2_n_12329, 
    instanceL2_n_12328, instanceL2_n_12327, instanceL2_n_12326, 
    instanceL2_n_12325, instanceL2_n_12324, instanceL2_n_12323, 
    instanceL2_n_12322, instanceL2_n_12321, instanceL2_n_12320, 
    instanceL2_n_12319, instanceL2_n_12318, instanceL2_n_12317, 
    instanceL2_n_12316, instanceL2_n_12315, instanceL2_n_12314, 
    instanceL2_n_12313, instanceL2_n_12312, instanceL2_n_12311, 
    instanceL2_n_12310, instanceL2_n_12309, instanceL2_n_12308, 
    instanceL2_n_12307, instanceL2_n_12306, instanceL2_n_12305, 
    instanceL2_n_12304, instanceL2_n_12303, instanceL2_n_12302, 
    instanceL2_n_12301, instanceL2_n_12300, instanceL2_n_12299, 
    instanceL2_n_12298, instanceL2_n_12297, instanceL2_n_12296, 
    instanceL2_n_12295, instanceL2_n_12294, instanceL2_n_12293, 
    instanceL2_n_12292, instanceL2_n_12291, instanceL2_n_12290, 
    instanceL2_n_12289, instanceL2_n_12288, instanceL2_n_12287, 
    instanceL2_n_12286, instanceL2_n_12285, instanceL2_n_12284, 
    instanceL2_n_12283, instanceL2_n_12282, instanceL2_n_12281, 
    instanceL2_n_12280, instanceL2_n_12279, instanceL2_n_12278, 
    instanceL2_n_12277, instanceL2_n_12276, instanceL2_n_12275, 
    instanceL2_n_12274, instanceL2_n_12273, instanceL2_n_12272, 
    instanceL2_n_12271, instanceL2_n_12270, instanceL2_n_12269, 
    instanceL2_n_12268, instanceL2_n_12267, instanceL2_n_12266, 
    instanceL2_n_12265, instanceL2_n_12264, instanceL2_n_12263, 
    instanceL2_n_12262, instanceL2_n_12261, instanceL2_n_12260, 
    instanceL2_n_12259, instanceL2_n_12258, instanceL2_n_12257, 
    instanceL2_n_12256, instanceL2_n_12255, instanceL2_n_12254, 
    instanceL2_n_12253, instanceL2_n_12252, instanceL2_n_12251, 
    instanceL2_n_12250, instanceL2_n_12249, instanceL2_n_12248, 
    instanceL2_n_12247, instanceL2_n_12246, instanceL2_n_12245, 
    instanceL2_n_12244, instanceL2_n_12243, instanceL2_n_12242, 
    instanceL2_n_12241, instanceL2_n_12240, instanceL2_n_12239, 
    instanceL2_n_12238, instanceL2_n_12237, instanceL2_n_12236, 
    instanceL2_n_12235, instanceL2_n_12234, instanceL2_n_12233, 
    instanceL2_n_12232, instanceL2_n_12231, instanceL2_n_12230, 
    instanceL2_n_12229, instanceL2_n_12228, instanceL2_n_12227, 
    instanceL2_n_12226, instanceL2_n_12225, instanceL2_n_12224, 
    instanceL2_n_12223, instanceL2_n_12222, instanceL2_n_12221, 
    instanceL2_n_12220, instanceL2_n_12219, instanceL2_n_12218, 
    instanceL2_n_12217, instanceL2_n_12216, instanceL2_n_12215, 
    instanceL2_n_12214, instanceL2_n_12213, instanceL2_n_12212, 
    instanceL2_n_12211, instanceL2_n_12210, instanceL2_n_12209, 
    instanceL2_n_12208, instanceL2_n_12207, instanceL2_n_12206, 
    instanceL2_n_12205, instanceL2_n_12204, instanceL2_n_12203, 
    instanceL2_n_12202, instanceL2_n_12201, instanceL2_n_12200, 
    instanceL2_n_12199, instanceL2_n_12198, instanceL2_n_12197, 
    instanceL2_n_12196, instanceL2_n_12195, instanceL2_n_12194, 
    instanceL2_n_12193, instanceL2_n_12192, instanceL2_n_12191, 
    instanceL2_n_12190, instanceL2_n_12189, instanceL2_n_12188, 
    instanceL2_n_12187, instanceL2_n_12186, instanceL2_n_12185, 
    instanceL2_n_12184, instanceL2_n_12183, instanceL2_n_12182, 
    instanceL2_n_12181, instanceL2_n_12180, instanceL2_n_12179, 
    instanceL2_n_12178, instanceL2_n_12177, instanceL2_n_12176, 
    instanceL2_n_12175, instanceL2_n_12174, instanceL2_n_12173, 
    instanceL2_n_12172, instanceL2_n_12171, instanceL2_n_12170, 
    instanceL2_n_12169, instanceL2_n_12168, instanceL2_n_12167, 
    instanceL2_n_12166, instanceL2_n_12165, instanceL2_n_12164, 
    instanceL2_n_12163, instanceL2_n_12162, instanceL2_n_12161, 
    instanceL2_n_12160, instanceL2_n_12159, instanceL2_n_12158, 
    instanceL2_n_12157, instanceL2_n_12156, instanceL2_n_12155, 
    instanceL2_n_12154, instanceL2_n_12153, instanceL2_n_12152, 
    instanceL2_n_12151, instanceL2_n_12150, instanceL2_n_12149, 
    instanceL2_n_12148, instanceL2_n_12147, instanceL2_n_12146, 
    instanceL2_n_12145, instanceL2_n_12144, instanceL2_n_12143, 
    instanceL2_n_12142, instanceL2_n_12141, instanceL2_n_12140, 
    instanceL2_n_12139, instanceL2_n_12138, instanceL2_n_12137, 
    instanceL2_n_12136, instanceL2_n_12135, instanceL2_n_12134, 
    instanceL2_n_12133, instanceL2_n_12132, instanceL2_n_12131, 
    instanceL2_n_12130, instanceL2_n_12129, instanceL2_n_12128, 
    instanceL2_n_12127, instanceL2_n_12126, instanceL2_n_12125, 
    instanceL2_n_12124, instanceL2_n_12123, instanceL2_n_12122, 
    instanceL2_n_12121, instanceL2_n_12120, instanceL2_n_12119, 
    instanceL2_n_12118, instanceL2_n_12117, instanceL2_n_12116, 
    instanceL2_n_12115, instanceL2_n_12114, instanceL2_n_12113, 
    instanceL2_n_12112, instanceL2_n_12111, instanceL2_n_12110, 
    instanceL2_n_12109, instanceL2_n_12108, instanceL2_n_12107, 
    instanceL2_n_12106, instanceL2_n_12105, instanceL2_n_12104, 
    instanceL2_n_12103, instanceL2_n_12102, instanceL2_n_12101, 
    instanceL2_n_12100, instanceL2_n_12099, instanceL2_n_12098, 
    instanceL2_n_12097, instanceL2_n_12096, instanceL2_n_12095, 
    instanceL2_n_12094, instanceL2_n_12093, instanceL2_n_12092, 
    instanceL2_n_12091, instanceL2_n_12090, instanceL2_n_12089, 
    instanceL2_n_12088, instanceL2_n_12087, instanceL2_n_12086, 
    instanceL2_n_12085, instanceL2_n_12084, instanceL2_n_12083, 
    instanceL2_n_12082, instanceL2_n_12081, instanceL2_n_12080, 
    instanceL2_n_12079, instanceL2_n_12078, instanceL2_n_12077, 
    instanceL2_n_12076, instanceL2_n_12075, instanceL2_n_12074, 
    instanceL2_n_12073, instanceL2_n_12072, instanceL2_n_12071, 
    instanceL2_n_12070, instanceL2_n_12069, instanceL2_n_12068, 
    instanceL2_n_12067, instanceL2_n_12066, instanceL2_n_12065, 
    instanceL2_n_12064, instanceL2_n_12063, instanceL2_n_12062, 
    instanceL2_n_12061, instanceL2_n_12060, instanceL2_n_12059, 
    instanceL2_n_12058, instanceL2_n_12057, instanceL2_n_12056, 
    instanceL2_n_12055, instanceL2_n_12054, instanceL2_n_12053, 
    instanceL2_n_12052, instanceL2_n_12051, instanceL2_n_12050, 
    instanceL2_n_12049, instanceL2_n_12048, instanceL2_n_12047, 
    instanceL2_n_12046, instanceL2_n_12045, instanceL2_n_12044, 
    instanceL2_n_12043, instanceL2_n_12042, instanceL2_n_12041, 
    instanceL2_n_12040, instanceL2_n_12039, instanceL2_n_12038, 
    instanceL2_n_12037, instanceL2_n_12036, instanceL2_n_12035, 
    instanceL2_n_12034, instanceL2_n_12033, instanceL2_n_12032, 
    instanceL2_n_12031, instanceL2_n_12030, instanceL2_n_12029, 
    instanceL2_n_12028, instanceL2_n_12027, instanceL2_n_12026, 
    instanceL2_n_12025, instanceL2_n_12024, instanceL2_n_12023, 
    instanceL2_n_12022, instanceL2_n_12021, instanceL2_n_12020, 
    instanceL2_n_12019, instanceL2_n_12018, instanceL2_n_12017, 
    instanceL2_n_12016, instanceL2_n_12015, instanceL2_n_12014, 
    instanceL2_n_12013, instanceL2_n_12012, instanceL2_n_12011, 
    instanceL2_n_12010, instanceL2_n_12009, instanceL2_n_12008, 
    instanceL2_n_12007, instanceL2_n_12006, instanceL2_n_12005, 
    instanceL2_n_12004, instanceL2_n_12003, instanceL2_n_12002, 
    instanceL2_n_12001, instanceL2_n_12000, instanceL2_n_11999, 
    instanceL2_n_11998, instanceL2_n_11997, instanceL2_n_11996, 
    instanceL2_n_11995, instanceL2_n_11994, instanceL2_n_11993, 
    instanceL2_n_11992, instanceL2_n_11991, instanceL2_n_11990, 
    instanceL2_n_11989, instanceL2_n_11988, instanceL2_n_11987, 
    instanceL2_n_11986, instanceL2_n_11985, instanceL2_n_11984, 
    instanceL2_n_11983, instanceL2_n_11982, instanceL2_n_11981, 
    instanceL2_n_11980, instanceL2_n_11979, instanceL2_n_11978, 
    instanceL2_n_11977, instanceL2_n_11976, instanceL2_n_11975, 
    instanceL2_n_11974, instanceL2_n_11973, instanceL2_n_11972, 
    instanceL2_n_11971, instanceL2_n_11970, instanceL2_n_11969, 
    instanceL2_n_11968, instanceL2_n_11967, instanceL2_n_11966, 
    instanceL2_n_11965, instanceL2_n_11964, instanceL2_n_11963, 
    instanceL2_n_11962, instanceL2_n_11961, instanceL2_n_11960, 
    instanceL2_n_11959, instanceL2_n_11958, instanceL2_n_11957, 
    instanceL2_n_11956, instanceL2_n_11955, instanceL2_n_11954, 
    instanceL2_n_11953, instanceL2_n_11952, instanceL2_n_11951, 
    instanceL2_n_11950, instanceL2_n_11949, instanceL2_n_11948, 
    instanceL2_n_11947, instanceL2_n_11946, instanceL2_n_11945, 
    instanceL2_n_11944, instanceL2_n_11943, instanceL2_n_11942, 
    instanceL2_n_11941, instanceL2_n_11940, instanceL2_n_11939, 
    instanceL2_n_11938, instanceL2_n_11937, instanceL2_n_11936, 
    instanceL2_n_11935, instanceL2_n_11934, instanceL2_n_11933, 
    instanceL2_n_11932, instanceL2_n_11931, instanceL2_n_11930, 
    instanceL2_n_11929, instanceL2_n_11928, instanceL2_n_11927, 
    instanceL2_n_11926, instanceL2_n_11925, instanceL2_n_11924, 
    instanceL2_n_11923, instanceL2_n_11922, instanceL2_n_11921, 
    instanceL2_n_11920, instanceL2_n_11919, instanceL2_n_11918, 
    instanceL2_n_11917, instanceL2_n_11916, instanceL2_n_11915, 
    instanceL2_n_11914, instanceL2_n_11913, instanceL2_n_11912, 
    instanceL2_n_11911, instanceL2_n_11910, instanceL2_n_11909, 
    instanceL2_n_11908, instanceL2_n_11907, instanceL2_n_11906, 
    instanceL2_n_11905, instanceL2_n_11904, instanceL2_n_11903, 
    instanceL2_n_11902, instanceL2_n_11901, instanceL2_n_11900, 
    instanceL2_n_11899, instanceL2_n_11898, instanceL2_n_11897, 
    instanceL2_n_11896, instanceL2_n_11895, instanceL2_n_11894, 
    instanceL2_n_11893, instanceL2_n_11892, instanceL2_n_11891, 
    instanceL2_n_11890, instanceL2_n_11889, instanceL2_n_11888, 
    instanceL2_n_11887, instanceL2_n_11886, instanceL2_n_11885, 
    instanceL2_n_11884, instanceL2_n_11883, instanceL2_n_11882, 
    instanceL2_n_11881, instanceL2_n_11880, instanceL2_n_11879, 
    instanceL2_n_11878, instanceL2_n_11877, instanceL2_n_11876, 
    instanceL2_n_11875, instanceL2_n_11874, instanceL2_n_11873, 
    instanceL2_n_11872, instanceL2_n_11871, instanceL2_n_11870, 
    instanceL2_n_11869, instanceL2_n_11868, instanceL2_n_11867, 
    instanceL2_n_11866, instanceL2_n_11865, instanceL2_n_11864, 
    instanceL2_n_11863, instanceL2_n_11862, instanceL2_n_11861, 
    instanceL2_n_11860, instanceL2_n_11859, instanceL2_n_11858, 
    instanceL2_n_11857, instanceL2_n_11856, instanceL2_n_11855, 
    instanceL2_n_11854, instanceL2_n_11853, instanceL2_n_11852, 
    instanceL2_n_11851, instanceL2_n_11850, instanceL2_n_11849, 
    instanceL2_n_11848, instanceL2_n_11847, instanceL2_n_11846, 
    instanceL2_n_11845, instanceL2_n_11844, instanceL2_n_11843, 
    instanceL2_n_11842, instanceL2_n_11841, instanceL2_n_11840, 
    instanceL2_n_11839, instanceL2_n_11838, instanceL2_n_11837, 
    instanceL2_n_11836, instanceL2_n_11835, instanceL2_n_11834, 
    instanceL2_n_11833, instanceL2_n_11832, instanceL2_n_11831, 
    instanceL2_n_11830, instanceL2_n_11829, instanceL2_n_11828, 
    instanceL2_n_11827, instanceL2_n_11826, instanceL2_n_11825, 
    instanceL2_n_11824, instanceL2_n_11823, instanceL2_n_11822, 
    instanceL2_n_11821, instanceL2_n_11820, instanceL2_n_11819, 
    instanceL2_n_11818, instanceL2_n_11817, instanceL2_n_11816, 
    instanceL2_n_11815, instanceL2_n_11814, instanceL2_n_11813, 
    instanceL2_n_11812, instanceL2_n_11811, instanceL2_n_11810, 
    instanceL2_n_11809, instanceL2_n_11808, instanceL2_n_11807, 
    instanceL2_n_11806, instanceL2_n_11805, instanceL2_n_11804, 
    instanceL2_n_11803, instanceL2_n_11802, instanceL2_n_11801, 
    instanceL2_n_11800, instanceL2_n_11799, instanceL2_n_11798, 
    instanceL2_n_11797, instanceL2_n_11796, instanceL2_n_11795, 
    instanceL2_n_11794, instanceL2_n_11793, instanceL2_n_11792, 
    instanceL2_n_11791, instanceL2_n_11790, instanceL2_n_11789, 
    instanceL2_n_11788, instanceL2_n_11787, instanceL2_n_11786, 
    instanceL2_n_11785, instanceL2_n_11784, instanceL2_n_11783, 
    instanceL2_n_11782, instanceL2_n_11781, instanceL2_n_11780, 
    instanceL2_n_11779, instanceL2_n_11778, instanceL2_n_11777, 
    instanceL2_n_11776, instanceL2_n_11775, instanceL2_n_11774, 
    instanceL2_n_11773, instanceL2_n_11772, instanceL2_n_11771, 
    instanceL2_n_11770, instanceL2_n_11769, instanceL2_n_11768, 
    instanceL2_n_11767, instanceL2_n_11766, instanceL2_n_11765, 
    instanceL2_n_11764, instanceL2_n_11763, instanceL2_n_11762, 
    instanceL2_n_11761, instanceL2_n_11760, instanceL2_n_11759, 
    instanceL2_n_11758, instanceL2_n_11757, instanceL2_n_11413, 
    instanceL2_n_11411, instanceL2_n_11409, instanceL2_n_11406, 
    instanceL2_n_11404, instanceL2_n_11403, instanceL2_n_11402, 
    instanceL2_n_11400, instanceL2_n_11398, instanceL2_n_11397, 
    instanceL2_n_11396, instanceL2_n_11395, instanceL2_n_11394, 
    instanceL2_n_11393, instanceL2_n_11392, instanceL2_n_11391, 
    instanceL2_n_11390, instanceL2_n_11389, instanceL2_n_11388, 
    instanceL2_n_11387, instanceL2_n_11386, instanceL2_n_11385, 
    instanceL2_n_11384, instanceL2_n_11383, instanceL2_n_11382, 
    instanceL2_n_11381, instanceL2_n_11380, instanceL2_n_11379, 
    instanceL2_n_11378, instanceL2_n_11377, instanceL2_n_11376, 
    instanceL2_n_11375, instanceL2_n_11374, instanceL2_n_11373, 
    instanceL2_n_11372, instanceL2_n_11371, instanceL2_n_11370, 
    instanceL2_n_11369, instanceL2_n_11368, instanceL2_n_11367, 
    instanceL2_n_11366, instanceL2_n_11365, instanceL2_n_11364, 
    instanceL2_n_11363, instanceL2_n_11362, instanceL2_n_11361, 
    instanceL2_n_11360, instanceL2_n_11359, instanceL2_n_11358, 
    instanceL2_n_11357, instanceL2_n_11356, instanceL2_n_11351, 
    instanceL2_n_11349, instanceL2_n_11348, instanceL2_n_11347, 
    instanceL2_n_11346, instanceL2_n_11345, instanceL2_n_11344, 
    instanceL2_n_11343, instanceL2_n_11341, instanceL2_n_11340, 
    instanceL2_n_11339, instanceL2_n_11338, instanceL2_n_11337, 
    instanceL2_n_11336, instanceL2_n_11334, instanceL2_n_11333, 
    instanceL2_n_11332, instanceL2_n_11331, instanceL2_n_11330, 
    instanceL2_n_11329, instanceL2_n_11328, instanceL2_n_11327, 
    instanceL2_n_11326, instanceL2_n_11325, instanceL2_n_11324, 
    instanceL2_n_11323, instanceL2_n_11322, instanceL2_n_11321, 
    instanceL2_n_11320, instanceL2_n_11319, instanceL2_n_11318, 
    instanceL2_n_11317, instanceL2_n_11316, instanceL2_n_11315, 
    instanceL2_n_11314, instanceL2_n_11313, instanceL2_n_11312, 
    instanceL2_n_11311, instanceL2_n_11310, instanceL2_n_11309, 
    instanceL2_n_11308, instanceL2_n_11307, instanceL2_n_11306, 
    instanceL2_n_11305, instanceL2_n_11304, instanceL2_n_11303, 
    instanceL2_n_11302, instanceL2_n_11301, instanceL2_n_11300, 
    instanceL2_n_11299, instanceL2_n_11298, instanceL2_n_11297, 
    instanceL2_n_11296, instanceL2_n_11295, instanceL2_n_11294, 
    instanceL2_n_11293, instanceL2_n_11292, instanceL2_n_11291, 
    instanceL2_n_11290, instanceL2_n_11289, instanceL2_n_11288, 
    instanceL2_n_11287, instanceL2_n_11286, instanceL2_n_11285, 
    instanceL2_n_11284, instanceL2_n_11283, instanceL2_n_11282, 
    instanceL2_n_11281, instanceL2_n_11280, instanceL2_n_11279, 
    instanceL2_n_11278, instanceL2_n_11277, instanceL2_n_11276, 
    instanceL2_n_11275, instanceL2_n_11274, instanceL2_n_11273, 
    instanceL2_n_11272, instanceL2_n_11271, instanceL2_n_11270, 
    instanceL2_n_11269, instanceL2_n_11268, instanceL2_n_11267, 
    instanceL2_n_11266, instanceL2_n_11265, instanceL2_n_11264, 
    instanceL2_n_11263, instanceL2_n_11262, instanceL2_n_11261, 
    instanceL2_n_11260, instanceL2_n_11259, instanceL2_n_11258, 
    instanceL2_n_11257, instanceL2_n_11256, instanceL2_n_11255, 
    instanceL2_n_11254, instanceL2_n_11253, instanceL2_n_11252, 
    instanceL2_n_11251, instanceL2_n_11250, instanceL2_n_11249, 
    instanceL2_n_11248, instanceL2_n_11247, instanceL2_n_11246, 
    instanceL2_n_11245, instanceL2_n_11244, instanceL2_n_11243, 
    instanceL2_n_11242, instanceL2_n_11241, instanceL2_n_11240, 
    instanceL2_n_11239, instanceL2_n_11238, instanceL2_n_11237, 
    instanceL2_n_11236, instanceL2_n_11235, instanceL2_n_11234, 
    instanceL2_n_11233, instanceL2_n_11232, instanceL2_n_11231, 
    instanceL2_n_11230, instanceL2_n_11229, instanceL2_n_11228, 
    instanceL2_n_11227, instanceL2_n_11226, instanceL2_n_11225, 
    instanceL2_n_11224, instanceL2_n_11223, instanceL2_n_11222, 
    instanceL2_n_11221, instanceL2_n_11220, instanceL2_n_11219, 
    instanceL2_n_11218, instanceL2_n_11217, instanceL2_n_11216, 
    instanceL2_n_11215, instanceL2_n_11214, instanceL2_n_11213, 
    instanceL2_n_11212, instanceL2_n_11211, instanceL2_n_11210, 
    instanceL2_n_11209, instanceL2_n_11208, instanceL2_n_11207, 
    instanceL2_n_11206, instanceL2_n_11205, instanceL2_n_11204, 
    instanceL2_n_11203, instanceL2_n_11202, instanceL2_n_11201, 
    instanceL2_n_11200, instanceL2_n_11199, instanceL2_n_11198, 
    instanceL2_n_11197, instanceL2_n_11196, instanceL2_n_11195, 
    instanceL2_n_11194, instanceL2_n_11193, instanceL2_n_11192, 
    instanceL2_n_11191, instanceL2_n_11190, instanceL2_n_11189, 
    instanceL2_n_11188, instanceL2_n_11187, instanceL2_n_11186, 
    instanceL2_n_11185, instanceL2_n_11184, instanceL2_n_11183, 
    instanceL2_n_11182, instanceL2_n_11181, instanceL2_n_11180, 
    instanceL2_n_11179, instanceL2_n_11178, instanceL2_n_11177, 
    instanceL2_n_11176, instanceL2_n_11175, instanceL2_n_11174, 
    instanceL2_n_11173, instanceL2_n_11172, instanceL2_n_11171, 
    instanceL2_n_11170, instanceL2_n_11169, instanceL2_n_11168, 
    instanceL2_n_11167, instanceL2_n_11166, instanceL2_n_11165, 
    instanceL2_n_11164, instanceL2_n_11163, instanceL2_n_11162, 
    instanceL2_n_11161, instanceL2_n_11160, instanceL2_n_11159, 
    instanceL2_n_11158, instanceL2_n_11157, instanceL2_n_11156, 
    instanceL2_n_11155, instanceL2_n_11154, instanceL2_n_11153, 
    instanceL2_n_11152, instanceL2_n_11151, instanceL2_n_11150, 
    instanceL2_n_11149, instanceL2_n_11148, instanceL2_n_11147, 
    instanceL2_n_11146, instanceL2_n_11145, instanceL2_n_11144, 
    instanceL2_n_11143, instanceL2_n_11142, instanceL2_n_11141, 
    instanceL2_n_11140, instanceL2_n_11139, instanceL2_n_11138, 
    instanceL2_n_11137, instanceL2_n_11136, instanceL2_n_11135, 
    instanceL2_n_11134, instanceL2_n_11133, instanceL2_n_11132, 
    instanceL2_n_11131, instanceL2_n_11130, instanceL2_n_11129, 
    instanceL2_n_11128, instanceL2_n_11127, instanceL2_n_11126, 
    instanceL2_n_11125, instanceL2_n_11124, instanceL2_n_11123, 
    instanceL2_n_11121, instanceL2_n_11120, instanceL2_n_11119, 
    instanceL2_n_11118, instanceL2_n_11117, instanceL2_n_11116, 
    instanceL2_n_11115, instanceL2_n_11114, instanceL2_n_11113, 
    instanceL2_n_11112, instanceL2_n_11111, instanceL2_n_11110, 
    instanceL2_n_11109, instanceL2_n_11108, instanceL2_n_11107, 
    instanceL2_n_11106, instanceL2_n_11105, instanceL2_n_11104, 
    instanceL2_n_11103, instanceL2_n_11102, instanceL2_n_11101, 
    instanceL2_n_11100, instanceL2_n_11099, instanceL2_n_11098, 
    instanceL2_n_11097, instanceL2_n_11096, instanceL2_n_11095, 
    instanceL2_n_11094, instanceL2_n_11092, instanceL2_n_11091, 
    instanceL2_n_11090, instanceL2_n_11089, instanceL2_n_11088, 
    instanceL2_n_11086, instanceL2_n_11085, instanceL2_n_11084, 
    instanceL2_n_11083, instanceL2_n_11080, instanceL2_n_11079, 
    instanceL2_n_11078, instanceL2_n_11077, instanceL2_n_11076, 
    instanceL2_n_11075, instanceL2_n_11074, instanceL2_n_11073, 
    instanceL2_n_11072, instanceL2_n_11071, instanceL2_n_11070, 
    instanceL2_n_11069, instanceL2_n_11068, instanceL2_n_11067, 
    instanceL2_n_11066, instanceL2_n_11065, instanceL2_n_11064, 
    instanceL2_n_11063, instanceL2_n_11062, instanceL2_n_11060, 
    instanceL2_n_11059, instanceL2_n_11058, instanceL2_n_11057, 
    instanceL2_n_11056, instanceL2_n_11055, instanceL2_n_11053, 
    instanceL2_n_11052, instanceL2_n_11051, instanceL2_n_11050, 
    instanceL2_n_11049, instanceL2_n_11048, instanceL2_n_11047, 
    instanceL2_n_11046, instanceL2_n_11045, instanceL2_n_11044, 
    instanceL2_n_11042, instanceL2_n_11041, instanceL2_n_11040, 
    instanceL2_n_11039, instanceL2_n_11038, instanceL2_n_11037, 
    instanceL2_n_11036, instanceL2_n_11035, instanceL2_n_11034, 
    instanceL2_n_11033, instanceL2_n_11032, instanceL2_n_11031, 
    instanceL2_n_11030, instanceL2_n_11029, instanceL2_n_11028, 
    instanceL2_n_11027, instanceL2_n_11026, instanceL2_n_11025, 
    instanceL2_n_11024, instanceL2_n_11023, instanceL2_n_11022, 
    instanceL2_n_11021, instanceL2_n_11020, instanceL2_n_11019, 
    instanceL2_n_11018, instanceL2_n_11017, instanceL2_n_11015, 
    instanceL2_n_11013, instanceL2_n_11012, instanceL2_n_11011, 
    instanceL2_n_11009, instanceL2_n_11008, instanceL2_n_11006, 
    instanceL2_n_11005, instanceL2_n_11004, instanceL2_n_11003, 
    instanceL2_n_11002, instanceL2_n_11001, instanceL2_n_11000, 
    instanceL2_n_10999, instanceL2_n_10997, instanceL2_n_10996, 
    instanceL2_n_10995, instanceL2_n_10994, instanceL2_n_10993, 
    instanceL2_n_10992, instanceL2_n_10991, instanceL2_n_10989, 
    instanceL2_n_10988, instanceL2_n_10987, instanceL2_n_10986, 
    instanceL2_n_10985, instanceL2_n_10984, instanceL2_n_10983, 
    instanceL2_n_10982, instanceL2_n_10981, instanceL2_n_10980, 
    instanceL2_n_10979, instanceL2_n_10978, instanceL2_n_10977, 
    instanceL2_n_10976, instanceL2_n_10975, instanceL2_n_10974, 
    instanceL2_n_10973, instanceL2_n_10972, instanceL2_n_10971, 
    instanceL2_n_10970, instanceL2_n_10969, instanceL2_n_10968, 
    instanceL2_n_10967, instanceL2_n_10966, instanceL2_n_10965, 
    instanceL2_n_10964, instanceL2_n_10963, instanceL2_n_10962, 
    instanceL2_n_10961, instanceL2_n_10960, instanceL2_n_10959, 
    instanceL2_n_10958, instanceL2_n_10957, instanceL2_n_10956, 
    instanceL2_n_10955, instanceL2_n_10954, instanceL2_n_10953, 
    instanceL2_n_10952, instanceL2_n_10951, instanceL2_n_10950, 
    instanceL2_n_10949, instanceL2_n_10948, instanceL2_n_10947, 
    instanceL2_n_10946, instanceL2_n_10945, instanceL2_n_10944, 
    instanceL2_n_10943, instanceL2_n_10942, instanceL2_n_10941, 
    instanceL2_n_10940, instanceL2_n_10939, instanceL2_n_10938, 
    instanceL2_n_10937, instanceL2_n_10936, instanceL2_n_10935, 
    instanceL2_n_10934, instanceL2_n_10933, instanceL2_n_10932, 
    instanceL2_n_10931, instanceL2_n_10929, instanceL2_n_10928, 
    instanceL2_n_10927, instanceL2_n_10926, instanceL2_n_10925, 
    instanceL2_n_10924, instanceL2_n_10923, instanceL2_n_10922, 
    instanceL2_n_10921, instanceL2_n_10920, instanceL2_n_10919, 
    instanceL2_n_10918, instanceL2_n_10917, instanceL2_n_10916, 
    instanceL2_n_10915, instanceL2_n_10914, instanceL2_n_10913, 
    instanceL2_n_10912, instanceL2_n_10911, instanceL2_n_10910, 
    instanceL2_n_10909, instanceL2_n_10908, instanceL2_n_10907, 
    instanceL2_n_10906, instanceL2_n_10905, instanceL2_n_10904, 
    instanceL2_n_10903, instanceL2_n_10902, instanceL2_n_10901, 
    instanceL2_n_10900, instanceL2_n_10899, instanceL2_n_10898, 
    instanceL2_n_10897, instanceL2_n_10896, instanceL2_n_10895, 
    instanceL2_n_10894, instanceL2_n_10893, instanceL2_n_10892, 
    instanceL2_n_10891, instanceL2_n_10890, instanceL2_n_10889, 
    instanceL2_n_10888, instanceL2_n_10887, instanceL2_n_10886, 
    instanceL2_n_10885, instanceL2_n_10884, instanceL2_n_10883, 
    instanceL2_n_10882, instanceL2_n_10881, instanceL2_n_10880, 
    instanceL2_n_10879, instanceL2_n_10878, instanceL2_n_10877, 
    instanceL2_n_10876, instanceL2_n_10875, instanceL2_n_10874, 
    instanceL2_n_10873, instanceL2_n_10872, instanceL2_n_10871, 
    instanceL2_n_10870, instanceL2_n_10869, instanceL2_n_10868, 
    instanceL2_n_10867, instanceL2_n_10866, instanceL2_n_10865, 
    instanceL2_n_10864, instanceL2_n_10863, instanceL2_n_10862, 
    instanceL2_n_10861, instanceL2_n_10860, instanceL2_n_10859, 
    instanceL2_n_10858, instanceL2_n_10857, instanceL2_n_10856, 
    instanceL2_n_10855, instanceL2_n_10854, instanceL2_n_10853, 
    instanceL2_n_10852, instanceL2_n_10851, instanceL2_n_10850, 
    instanceL2_n_10849, instanceL2_n_10848, instanceL2_n_10847, 
    instanceL2_n_10846, instanceL2_n_10845, instanceL2_n_10844, 
    instanceL2_n_10843, instanceL2_n_10842, instanceL2_n_10841, 
    instanceL2_n_10840, instanceL2_n_10839, instanceL2_n_10838, 
    instanceL2_n_10836, instanceL2_n_10835, instanceL2_n_10834, 
    instanceL2_n_10833, instanceL2_n_10832, instanceL2_n_10831, 
    instanceL2_n_10830, instanceL2_n_10829, instanceL2_n_10828, 
    instanceL2_n_10827, instanceL2_n_10826, instanceL2_n_10825, 
    instanceL2_n_10824, instanceL2_n_10823, instanceL2_n_10821, 
    instanceL2_n_10820, instanceL2_n_10817, instanceL2_n_10816, 
    instanceL2_n_10815, instanceL2_n_10814, instanceL2_n_10812, 
    instanceL2_n_10811, instanceL2_n_10810, instanceL2_n_10809, 
    instanceL2_n_10808, instanceL2_n_10807, instanceL2_n_10806, 
    instanceL2_n_10805, instanceL2_n_10804, instanceL2_n_10802, 
    instanceL2_n_10801, instanceL2_n_10800, instanceL2_n_10797, 
    instanceL2_n_10795, instanceL2_n_10794, instanceL2_n_10793, 
    instanceL2_n_10791, instanceL2_n_10790, instanceL2_n_10787, 
    instanceL2_n_10786, instanceL2_n_10785, instanceL2_n_10784, 
    instanceL2_n_10783, instanceL2_n_10780, instanceL2_n_10779, 
    instanceL2_n_10775, instanceL2_n_10773, instanceL2_n_10772, 
    instanceL2_n_10771, instanceL2_n_10770, instanceL2_n_10768, 
    instanceL2_n_10766, instanceL2_n_10763, instanceL2_n_10757, 
    instanceL2_n_10755, instanceL2_n_10753, instanceL2_n_10751, 
    instanceL2_n_10750, instanceL2_n_10740, instanceL2_n_10738, 
    instanceL2_n_10734, instanceL2_n_10730, instanceL2_n_10725, 
    instanceL2_n_10723, instanceL2_n_10719, instanceL2_n_10716, 
    instanceL2_n_10711, instanceL2_n_10708, instanceL2_n_10704, 
    instanceL2_n_10701, UNCONNECTED412, UNCONNECTED411, UNCONNECTED410, 
    UNCONNECTED409, UNCONNECTED408, UNCONNECTED407, UNCONNECTED406, 
    UNCONNECTED405, UNCONNECTED404, UNCONNECTED403, UNCONNECTED402, 
    UNCONNECTED401, UNCONNECTED400, UNCONNECTED399, UNCONNECTED398, 
    UNCONNECTED397, UNCONNECTED396, UNCONNECTED395, UNCONNECTED394, 
    UNCONNECTED393, UNCONNECTED392, UNCONNECTED391, UNCONNECTED390, 
    UNCONNECTED389, UNCONNECTED388, UNCONNECTED387, UNCONNECTED386, 
    UNCONNECTED385, UNCONNECTED384, UNCONNECTED383, UNCONNECTED382, 
    UNCONNECTED381, UNCONNECTED380, UNCONNECTED379, UNCONNECTED378, 
    UNCONNECTED377, UNCONNECTED376, UNCONNECTED375, UNCONNECTED374, 
    UNCONNECTED373, UNCONNECTED372, UNCONNECTED371, UNCONNECTED370, 
    UNCONNECTED369, UNCONNECTED368, UNCONNECTED367, UNCONNECTED366, 
    UNCONNECTED365, UNCONNECTED364, UNCONNECTED363, UNCONNECTED362, 
    UNCONNECTED361, UNCONNECTED360, UNCONNECTED359, done, updown, rst_n, clk;
wire   [18:0] \instanceL2_row_sums[0] ;
wire   [18:0] \instanceL2_row_sums[1] ;
wire   [13:0] \instanceL2_prod_terms[1][3] ;
wire   [13:0] \instanceL2_prod_terms[1][4] ;
wire   [13:0] \instanceL2_prod_terms[1][5] ;
wire   [13:0] \instanceL2_prod_terms[1][6] ;
wire   [13:0] \instanceL2_prod_terms[1][11] ;
wire   [13:0] \instanceL2_prod_terms[1][13] ;
wire   [13:0] \instanceL2_prod_terms[1][14] ;
wire   [13:0] \instanceL2_prod_terms[1][16] ;
wire   [18:0] \instanceL2_row_sums[2] ;
wire   [13:0] \instanceL2_prod_terms[2][0] ;
wire   [13:0] \instanceL2_prod_terms[2][16] ;
wire   [18:0] \instanceL2_row_sums[3] ;
wire   [13:0] \instanceL2_prod_terms[3][6] ;
wire   [13:0] \instanceL2_prod_terms[3][8] ;
wire   [13:0] \instanceL2_prod_terms[3][9] ;
wire   [13:0] \instanceL2_prod_terms[3][17] ;
wire   [13:0] \instanceL2_prod_terms[3][18] ;
wire   [18:0] \instanceL2_row_sums[4] ;
wire   [13:0] \instanceL2_prod_terms[4][2] ;
wire   [13:0] \instanceL2_prod_terms[4][6] ;
wire   [13:0] \instanceL2_prod_terms[4][11] ;
wire   [18:0] \instanceL2_row_sums[5] ;
wire   [13:0] \instanceL2_prod_terms[2][3] ;
wire   [13:0] \instanceL2_prod_terms[5][12] ;
wire   [13:0] \instanceL2_prod_terms[5][17] ;
wire   [13:0] \instanceL2_prod_terms[5][19] ;
wire   [18:0] \instanceL2_row_sums[6] ;
wire   [13:0] \instanceL2_prod_terms[6][2] ;
wire   [13:0] \instanceL2_prod_terms[6][5] ;
wire   [13:0] \instanceL2_prod_terms[3][7] ;
wire   [13:0] \instanceL2_prod_terms[2][9] ;
wire   [13:0] \instanceL2_prod_terms[6][10] ;
wire   [13:0] \instanceL2_prod_terms[6][11] ;
wire   [13:0] \instanceL2_prod_terms[4][12] ;
wire   [13:0] \instanceL2_prod_terms[6][13] ;
wire   [13:0] \instanceL2_prod_terms[6][15] ;
wire   [18:0] \instanceL2_row_sums[7] ;
wire   [13:0] \instanceL2_prod_terms[6][1] ;
wire   [13:0] \instanceL2_prod_terms[7][3] ;
wire   [13:0] \instanceL2_prod_terms[7][4] ;
wire   [13:0] \instanceL2_prod_terms[5][4] ;
wire   [13:0] \instanceL2_prod_terms[7][5] ;
wire   [13:0] \instanceL2_prod_terms[2][6] ;
wire   [13:0] \instanceL2_prod_terms[3][12] ;
wire   [13:0] \instanceL2_prod_terms[7][12] ;
wire   [13:0] \instanceL2_prod_terms[7][15] ;
wire   [13:0] \instanceL2_prod_terms[7][17] ;
wire   [13:0] \instanceL2_prod_terms[7][18] ;
wire   [18:0] \instanceL2_row_sums[8] ;
wire   [13:0] \instanceL2_prod_terms[8][0] ;
wire   [13:0] \instanceL2_prod_terms[8][2] ;
wire   [13:0] \instanceL2_prod_terms[7][2] ;
wire   [13:0] \instanceL2_prod_terms[8][7] ;
wire   [13:0] \instanceL2_prod_terms[6][8] ;
wire   [13:0] \instanceL2_prod_terms[8][11] ;
wire   [13:0] \instanceL2_prod_terms[8][14] ;
wire   [13:0] \instanceL2_prod_terms[4][14] ;
wire   [13:0] \instanceL2_prod_terms[1][15] ;
wire   [13:0] \instanceL2_prod_terms[8][15] ;
wire   [13:0] \instanceL2_prod_terms[8][18] ;
wire   [13:0] \instanceL2_prod_terms[4][18] ;
wire   [13:0] \instanceL2_prod_terms[8][19] ;
wire   [13:0] \instanceL2_prod_terms[1][19] ;
wire   [18:0] \instanceL2_row_sums[9] ;
wire   [13:0] \instanceL2_prod_terms[2][1] ;
wire   [13:0] \instanceL2_prod_terms[9][1] ;
wire   [13:0] \instanceL2_prod_terms[9][2] ;
wire   [13:0] \instanceL2_prod_terms[9][3] ;
wire   [13:0] \instanceL2_prod_terms[9][4] ;
wire   [13:0] \instanceL2_prod_terms[5][5] ;
wire   [13:0] \instanceL2_prod_terms[2][5] ;
wire   [13:0] \instanceL2_prod_terms[9][5] ;
wire   [13:0] \instanceL2_prod_terms[4][7] ;
wire   [13:0] \instanceL2_prod_terms[0][7] ;
wire   [13:0] \instanceL2_prod_terms[9][8] ;
wire   [13:0] \instanceL2_prod_terms[9][12] ;
wire   [13:0] \instanceL2_prod_terms[2][13] ;
wire   [13:0] \instanceL2_prod_terms[5][13] ;
wire   [13:0] \instanceL2_prod_terms[9][13] ;
wire   [13:0] \instanceL2_prod_terms[3][14] ;
wire   [13:0] \instanceL2_prod_terms[9][15] ;
wire   [13:0] \instanceL2_prod_terms[9][16] ;
wire   [13:0] \instanceL2_prod_terms[4][17] ;
wire   [13:0] \instanceL2_prod_terms[9][17] ;
wire   [13:0] \instanceL2_prod_terms[9][18] ;
wire   [1:0] counter;
wire   [179:0] layer2_out;
wire   [3:0] out;
wire   [179:0] layer1_out;
wire   [0:9] out_activehigh;
wire   [127:0] in;
  layer1 instanceL1(.clk(clk), .rst_n(rst_n), .updown(updown), .in({ in[127:0] }), .out({
    UNCONNECTED373,  layer1_out[178:171] , UNCONNECTED372,  layer1_out[169:153] , UNCONNECTED371,  layer1_out[151:144] , UNCONNECTED370,  layer1_out[142:135] , 
    UNCONNECTED369,  layer1_out[133:126] , UNCONNECTED368,  layer1_out[124:117] , UNCONNECTED367,  layer1_out[115:108] , UNCONNECTED366,  layer1_out[106:99] , 
    UNCONNECTED365,  layer1_out[97:72] , UNCONNECTED364,  layer1_out[70:54] , UNCONNECTED363,  layer1_out[52:45] , UNCONNECTED362,  layer1_out[43:36] , 
    UNCONNECTED361,  layer1_out[34:18] , UNCONNECTED360,  layer1_out[16:9] , UNCONNECTED359,  layer1_out[7:0] }));
  csa_tree_ADD_TC_OP_19_group_17897 instanceL2_csa_tree_ADD_TC_OP_19_groupi(
    .in_0({1'b0, 1'b0, \instanceL2_prod_terms[0][19][13] , 
    \instanceL2_prod_terms[0][19][10] , \instanceL2_prod_terms[0][19][9] , 
    \instanceL2_prod_terms[0][19][8] , \instanceL2_prod_terms[0][19][7] , 
    \instanceL2_prod_terms[0][19][6] , \instanceL2_prod_terms[0][19][5] , 
    \instanceL2_prod_terms[0][19][4] , \instanceL2_prod_terms[0][19][3] , 
    \instanceL2_prod_terms[0][19][2] , \instanceL2_prod_terms[0][19][1] , 
    layer1_out[171]}), .in_1({1'b0, \instanceL2_prod_terms[9][18] [13],  \instanceL2_prod_terms[9][18] [11:1] , 
    layer1_out[162]}), .in_2({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[9][17] [10:2] , 
    \instanceL2_prod_terms[4][17] [1], layer1_out[153]}), .in_3({1'b0, 1'b0,  \instanceL2_prod_terms[9][16] [11:3] ,  layer1_out[145:144] , 
    1'b0}), .in_4({1'b0, 1'b0,  \instanceL2_prod_terms[9][15] [11:3] ,  layer1_out[137:135] }), .in_5({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[3][14] [10:2] ,  layer1_out[127:126] }), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, \instanceL2_prod_terms[9][13] [13], 
    \instanceL2_prod_terms[9][13] [8],  \instanceL2_prod_terms[5][13] [8:5] ,  \instanceL2_prod_terms[2][13] [2:1] , layer1_out[117], 1'b0}), .in_7({1'b0, 
    \instanceL2_prod_terms[9][12] [13],  \instanceL2_prod_terms[9][12] [11:1] , layer1_out[108]}), .in_8({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[97:90] , 1'b0}), .in_10({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0,  layer1_out[89:81] }), .in_11({1'b0, \instanceL2_prod_terms[9][8] [13],  \instanceL2_prod_terms[9][8] [11:1] , 
    layer1_out[72]}), .in_12({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , 
    layer1_out[63], 1'b0, 1'b0}), .in_13({1'b0, 1'b0, 1'b0,  layer1_out[62:54] , 1'b0, 1'b0}),
     .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[9][5] [13],  \instanceL2_prod_terms[2][5] [8:6] , 
    \instanceL2_prod_terms[5][5] [6],  \instanceL2_prod_terms[2][5] [4:2] , layer1_out[45]}), .in_15({1'b0, 
    \instanceL2_prod_terms[9][4] [13],  \instanceL2_prod_terms[9][4] [11:1] , layer1_out[36]}), .in_16({1'b0, 1'b0,  \instanceL2_prod_terms[9][3] [11:3] ,  layer1_out[29:27] }),
     .in_17({ \instanceL2_prod_terms[9][2] [13:1] , layer1_out[18]}), .in_18({1'b0, 1'b0, 
    \instanceL2_prod_terms[0][0][13] , \instanceL2_prod_terms[0][0][8] , 
    \instanceL2_prod_terms[0][0][7] , \instanceL2_prod_terms[0][0][6] , 
    \instanceL2_prod_terms[0][0][5] , \instanceL2_prod_terms[0][0][4] , 
    \instanceL2_prod_terms[0][0][3] , \instanceL2_prod_terms[0][0][2] , 
    layer1_out[0], 1'b0, 1'b0, 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[9][1] [10], \instanceL2_prod_terms[0][1][8] ,  \instanceL2_prod_terms[9][1] [8:6] , 
    \instanceL2_prod_terms[0][1][4] ,  \instanceL2_prod_terms[9][1] [4:3] , \instanceL2_prod_terms[2][1] [1], 
    layer1_out[9], 1'b0}), .out_0({ \instanceL2_row_sums[9] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_8228_1 instanceL2_csa_tree_ADD_TC_OP_19_groupi823(
    .in_0({1'b0, \instanceL2_prod_terms[1][19] [13],  \instanceL2_prod_terms[8][19] [11:2] , 
    \instanceL2_prod_terms[1][19] [3], layer1_out[171]}), .in_1({1'b0, 1'b0, 
    \instanceL2_prod_terms[4][18] [13],  \instanceL2_prod_terms[8][18] [10:3] ,  layer1_out[163:162] , 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[4][17] [13],  \instanceL2_prod_terms[4][17] [8:1] , layer1_out[153]}), .in_3({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][16][13] , 
    \instanceL2_prod_terms[0][16][7] , \instanceL2_prod_terms[0][16][6] , 
    \instanceL2_prod_terms[0][16][5] , \instanceL2_prod_terms[0][16][4] , 
    \instanceL2_prod_terms[0][16][3] , \instanceL2_prod_terms[0][16][2] , 
    \instanceL2_prod_terms[0][16][1] , layer1_out[144]}), .in_4({1'b0, 1'b0, 
    1'b0,  \instanceL2_prod_terms[8][15] [10:3] , \instanceL2_prod_terms[1][15] [1], layer1_out[135], 1'b0}), .in_5({
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[4][14] [13],  \instanceL2_prod_terms[8][14] [9:3] , 
    \instanceL2_prod_terms[3][14] [2],  layer1_out[127:126] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[124:117] , 
    1'b0}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_8({1'b0, \instanceL2_prod_terms[0][11][13] ,  \instanceL2_prod_terms[8][11] [11:5] , 
    \instanceL2_prod_terms[2][11][2] ,  layer1_out[100:99] , 1'b0, 1'b0}), .in_9({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_10({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[89:81] }), .in_11({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[6][8] [10:2] , 
    \instanceL2_prod_terms[1][8][2] , layer1_out[72]}), .in_12({1'b0, 1'b0,  \instanceL2_prod_terms[8][7] [11:3] ,  layer1_out[64:63] , 
    1'b0}), .in_13({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[62:54] , 1'b0}), .in_14({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0,  layer1_out[52:45] }), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[34:27] , 
    1'b0}), .in_17({1'b0, 1'b0, \instanceL2_prod_terms[7][2] [13],  \instanceL2_prod_terms[7][2] [8:7] ,  \instanceL2_prod_terms[8][2] [8:4] , 
    \instanceL2_prod_terms[7][2] [1], layer1_out[18], 1'b0, 1'b0}), .in_18({
    1'b0, 1'b0, \instanceL2_prod_terms[0][0][13] ,  \instanceL2_prod_terms[8][0] [10:3] ,  layer1_out[2:0] }), .in_19({1'b0, 1'b0, 1'b0, 
    1'b0,  layer1_out[16:9] , 1'b0, 1'b0}), .out_0({ \instanceL2_row_sums[8] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_14031 instanceL2_csa_tree_ADD_TC_OP_19_groupi824(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[7][18] [9:2] , 
    \instanceL2_prod_terms[4][18] [3], layer1_out[162]}), .in_2({ \instanceL2_prod_terms[7][17] [13:1] , 
    layer1_out[153]}), .in_3({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[151:144] , 1'b0, 1'b0}), .in_4({
    1'b0, \instanceL2_prod_terms[7][15] [13],  \instanceL2_prod_terms[7][15] [11:1] , layer1_out[135]}), .in_5({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[133:126] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_7({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[7][12] [10:3] , 
    \instanceL2_prod_terms[3][12] [3], layer1_out[108], 1'b0}), .in_8({1'b0, 
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][11][13] , 
    \instanceL2_prod_terms[0][11][7] , \instanceL2_prod_terms[0][11][6] , 
    \instanceL2_prod_terms[0][11][5] , \instanceL2_prod_terms[0][11][4] , 
    \instanceL2_prod_terms[0][11][3] , \instanceL2_prod_terms[0][11][2] , 
    \instanceL2_prod_terms[0][11][1] , layer1_out[99], 1'b0}), .in_9({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0}), .in_10({1'b0, \instanceL2_prod_terms[7][9][12] , 
    \instanceL2_prod_terms[7][9][11] , \instanceL2_prod_terms[7][9][10] , 
    \instanceL2_prod_terms[7][9][9] , \instanceL2_prod_terms[7][9][8] , 
    \instanceL2_prod_terms[7][9][7] , \instanceL2_prod_terms[7][9][6] , 
    \instanceL2_prod_terms[7][9][5] , \instanceL2_prod_terms[7][9][4] , 
    \instanceL2_prod_terms[7][9][3] ,  layer1_out[83:81] }), .in_11({1'b0, 1'b0, 
    \instanceL2_prod_terms[2][8][11] , \instanceL2_prod_terms[2][8][10] , 
    \instanceL2_prod_terms[2][8][9] , \instanceL2_prod_terms[2][8][8] , 
    \instanceL2_prod_terms[2][8][7] , \instanceL2_prod_terms[2][8][6] , 
    \instanceL2_prod_terms[2][8][5] , \instanceL2_prod_terms[2][8][4] , 
    \instanceL2_prod_terms[2][8][3] , \instanceL2_prod_terms[2][8][2] ,  layer1_out[73:72] }),
     .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , 
    \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , layer1_out[63]}), .in_13({1'b0, 
    \instanceL2_prod_terms[2][6] [13],  \instanceL2_prod_terms[2][6] [11:3] ,  layer1_out[55:54] , 1'b0}), .in_14({1'b0, 1'b0, 
    \instanceL2_prod_terms[9][5] [13],  \instanceL2_prod_terms[7][5] [10:3] ,  layer1_out[47:45] }), .in_15({1'b0, 1'b0, 
    \instanceL2_prod_terms[5][4] [13],  \instanceL2_prod_terms[7][4] [10:3] ,  layer1_out[38:36] }), .in_16({1'b0, 
    \instanceL2_prod_terms[7][3] [13],  \instanceL2_prod_terms[7][3] [11:1] , layer1_out[27]}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, \instanceL2_prod_terms[7][2] [13],  \instanceL2_prod_terms[7][2] [8:7] ,  \instanceL2_prod_terms[8][2] [8:4] , 
    \instanceL2_prod_terms[7][2] [1], layer1_out[18]}), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .in_19({1'b0, 1'b0,  \instanceL2_prod_terms[6][1] [11:3] ,  layer1_out[11:9] }), .out_0({ \instanceL2_row_sums[7] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_12094 instanceL2_csa_tree_ADD_TC_OP_19_groupi825(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[178:171] }), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0,  layer1_out[169:162] }), .in_2({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[4][17] [13],  \instanceL2_prod_terms[4][17] [8:1] , 
    layer1_out[153], 1'b0}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][16][13] , \instanceL2_prod_terms[0][16][7] , 
    \instanceL2_prod_terms[0][16][6] , \instanceL2_prod_terms[0][16][5] , 
    \instanceL2_prod_terms[0][16][4] , \instanceL2_prod_terms[0][16][3] , 
    \instanceL2_prod_terms[0][16][2] , \instanceL2_prod_terms[0][16][1] , 
    layer1_out[144]}), .in_4({1'b0, \instanceL2_prod_terms[6][15] [13],  \instanceL2_prod_terms[6][15] [11:4] ,  \instanceL2_prod_terms[8][15] [4:3] , 
    \instanceL2_prod_terms[1][15] [1], layer1_out[135]}), .in_5({1'b0, 1'b0, 
    1'b0, \instanceL2_prod_terms[4][14] [13],  \instanceL2_prod_terms[4][14] [7:1] , layer1_out[126], 1'b0, 1'b0}),
     .in_6({1'b0, 1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[6][13] [9:2] , \instanceL2_prod_terms[2][13] [1], 
    layer1_out[117]}), .in_7({1'b0, 1'b0, \instanceL2_prod_terms[3][12] [13],  \instanceL2_prod_terms[4][12] [10:3] ,  layer1_out[110:108] }),
     .in_8({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[6][11] [10:3] , \instanceL2_prod_terms[0][11][1] , layer1_out[99], 
    1'b0}), .in_9({1'b0, \instanceL2_prod_terms[6][10] [13],  \instanceL2_prod_terms[6][10] [11:1] , layer1_out[90]}),
     .in_10({1'b0, 1'b0, \instanceL2_prod_terms[2][9] [13],  \instanceL2_prod_terms[2][9] [10:3] , layer1_out[81], 
    1'b0, 1'b0}), .in_11({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[6][8] [10:2] , \instanceL2_prod_terms[1][8][2] , 
    layer1_out[72]}), .in_12({1'b0, 1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[3][7] [9:2] , 
    \instanceL2_prod_terms[0][7] [2], layer1_out[63]}), .in_13({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .in_14({1'b0, \instanceL2_prod_terms[6][5] [13],  \instanceL2_prod_terms[6][5] [11:2] , layer1_out[45], 1'b0}),
     .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[43:36] }), .in_16({1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0,  layer1_out[34:27] }), .in_17({ \instanceL2_prod_terms[6][2] [13:2] , layer1_out[18], 1'b0}), .in_18({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0,  layer1_out[7:0] , 1'b0}), .in_19({1'b0, 1'b0,  \instanceL2_prod_terms[6][1] [11:3] ,  layer1_out[11:9] }), .out_0({ \instanceL2_row_sums[6] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_10152 instanceL2_csa_tree_ADD_TC_OP_19_groupi826(
    .in_0({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[5][19] [10:3] ,  \instanceL2_prod_terms[1][19] [4:3] , layer1_out[171]}), .in_1({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[4][18] [13],  \instanceL2_prod_terms[4][18] [9:3] , layer1_out[162], 1'b0, 1'b0}), .in_2({ \instanceL2_prod_terms[5][17] [13:2] , 
    layer1_out[153], 1'b0}), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][16][13] , \instanceL2_prod_terms[0][16][7] , 
    \instanceL2_prod_terms[0][16][6] , \instanceL2_prod_terms[0][16][5] , 
    \instanceL2_prod_terms[0][16][4] , \instanceL2_prod_terms[0][16][3] , 
    \instanceL2_prod_terms[0][16][2] , \instanceL2_prod_terms[0][16][1] , 
    layer1_out[144], 1'b0}), .in_4({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[1][15] [10:1] , layer1_out[135]}), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][14][9] , 
    \instanceL2_prod_terms[0][14][8] , \instanceL2_prod_terms[0][14][7] , 
    \instanceL2_prod_terms[0][14][6] , \instanceL2_prod_terms[0][14][5] , 
    \instanceL2_prod_terms[0][14][4] , \instanceL2_prod_terms[0][14][3] , 
    \instanceL2_prod_terms[0][14][2] , \instanceL2_prod_terms[4][14] [1], 
    layer1_out[126]}), .in_6({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[9][13] [13], \instanceL2_prod_terms[9][13] [8],  \instanceL2_prod_terms[5][13] [8:5] ,  \instanceL2_prod_terms[2][13] [2:1] , 
    layer1_out[117], 1'b0, 1'b0}), .in_7({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[3][12] [13],  \instanceL2_prod_terms[5][12] [9:2] ,  layer1_out[109:108] }), .in_8({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][11][13] , \instanceL2_prod_terms[0][11][7] , 
    \instanceL2_prod_terms[0][11][6] , \instanceL2_prod_terms[0][11][5] , 
    \instanceL2_prod_terms[0][11][4] , \instanceL2_prod_terms[0][11][3] , 
    \instanceL2_prod_terms[0][11][2] , \instanceL2_prod_terms[0][11][1] , 
    layer1_out[99], 1'b0, 1'b0}), .in_9({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[97:90] , 1'b0, 1'b0}),
     .in_10({1'b0, 1'b0, \instanceL2_prod_terms[2][9] [13],  \instanceL2_prod_terms[2][9] [10:3] , layer1_out[81], 
    1'b0, 1'b0}), .in_11({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[1][8][13] , 
    \instanceL2_prod_terms[1][8][9] , \instanceL2_prod_terms[1][8][8] , 
    \instanceL2_prod_terms[1][8][7] , \instanceL2_prod_terms[1][8][6] , 
    \instanceL2_prod_terms[1][8][5] , \instanceL2_prod_terms[1][8][4] , 
    \instanceL2_prod_terms[1][8][3] , \instanceL2_prod_terms[1][8][2] , 
    layer1_out[72], 1'b0}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_13({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[62:54] , 
    1'b0}), .in_14({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[9][5] [13],  \instanceL2_prod_terms[2][5] [8:6] , 
    \instanceL2_prod_terms[5][5] [6],  \instanceL2_prod_terms[2][5] [4:2] , layer1_out[45], 1'b0, 1'b0}), .in_15({
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[5][4] [13],  \instanceL2_prod_terms[5][4] [9:3] , layer1_out[36], 1'b0, 
    1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[2][3] [13],  \instanceL2_prod_terms[2][3] [7:1] , layer1_out[27]}), .in_17({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0,  layer1_out[26:18] }), .in_18({1'b0, 1'b0, 1'b0,  layer1_out[7:0] , 1'b0, 1'b0, 1'b0}), .in_19({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[16:9] , 1'b0}), .out_0({ \instanceL2_row_sums[5] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_8228 instanceL2_csa_tree_ADD_TC_OP_19_groupi827(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[178:171] , 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[4][18] [13],  \instanceL2_prod_terms[4][18] [9:3] , layer1_out[162], 1'b0, 1'b0}), .in_2({
    1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[4][17] [13],  \instanceL2_prod_terms[4][17] [8:1] , layer1_out[153]}),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][16][13] , 
    \instanceL2_prod_terms[0][16][7] , \instanceL2_prod_terms[0][16][6] , 
    \instanceL2_prod_terms[0][16][5] , \instanceL2_prod_terms[0][16][4] , 
    \instanceL2_prod_terms[0][16][3] , \instanceL2_prod_terms[0][16][2] , 
    \instanceL2_prod_terms[0][16][1] , layer1_out[144], 1'b0}), .in_4({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[142:135] , 1'b0}), .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[4][14] [13],  \instanceL2_prod_terms[4][14] [7:1] , layer1_out[126]}), .in_6({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[124:117] }), .in_7({1'b0, 1'b0, 
    \instanceL2_prod_terms[3][12] [13],  \instanceL2_prod_terms[4][12] [10:3] ,  layer1_out[110:108] }), .in_8({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[4][11] [10:3] , 
    \instanceL2_prod_terms[2][11][2] ,  layer1_out[100:99] }), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_10({1'b0, 1'b0, 
    1'b0, \instanceL2_prod_terms[2][9] [13],  \instanceL2_prod_terms[2][9] [10:3] , layer1_out[81], 1'b0}), .in_11({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[80:72] }), .in_12({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , 
    layer1_out[63], 1'b0, 1'b0}), .in_13({1'b0, 1'b0,  \instanceL2_prod_terms[4][6] [11:3] , 
    \instanceL2_prod_terms[2][6] [3],  layer1_out[55:54] }), .in_14({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[52:45] , 
    1'b0}), .in_15({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[43:36] , 1'b0, 1'b0}), .in_16({1'b0, 1'b0, 
    1'b0, \instanceL2_prod_terms[2][3] [13], \instanceL2_prod_terms[0][3][9] , 
    \instanceL2_prod_terms[0][3][8] , \instanceL2_prod_terms[0][3][7] , 
    \instanceL2_prod_terms[0][3][6] , \instanceL2_prod_terms[0][3][5] , 
    \instanceL2_prod_terms[0][3][4] , \instanceL2_prod_terms[0][3][3] , 
    \instanceL2_prod_terms[0][3][2] ,  layer1_out[28:27] }), .in_17({1'b0,  \instanceL2_prod_terms[4][2] [12:3] ,  layer1_out[19:18] , 1'b0}), .in_18({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[16:9] , 1'b0}), .out_0({ \instanceL2_row_sums[4] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_6301 instanceL2_csa_tree_ADD_TC_OP_19_groupi828(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[178:171] , 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[3][18] [10:3] ,  \instanceL2_prod_terms[4][18] [4:3] , 
    layer1_out[162]}), .in_2({1'b0, 1'b0,  \instanceL2_prod_terms[3][17] [11:3] , \instanceL2_prod_terms[0][17][2] ,  layer1_out[154:153] }),
     .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[151:144] }), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_5({1'b0, 
    1'b0, 1'b0,  \instanceL2_prod_terms[3][14] [10:2] ,  layer1_out[127:126] }), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_7({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[3][12] [13],  \instanceL2_prod_terms[3][12] [9:3] , layer1_out[108], 1'b0, 1'b0}), .in_8({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[106:99] , 1'b0}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_10({1'b0, 1'b0, 
    1'b0,  \instanceL2_prod_terms[3][9] [10:2] , \instanceL2_prod_terms[2][9] [3], layer1_out[81]}), .in_11({ \instanceL2_prod_terms[3][8] [13:1] , 
    layer1_out[72]}), .in_12({1'b0, 1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[3][7] [9:2] , 
    \instanceL2_prod_terms[0][7] [2], layer1_out[63]}), .in_13({1'b0, 1'b0, 
    \instanceL2_prod_terms[2][6] [13],  \instanceL2_prod_terms[3][6] [10:3] , layer1_out[54], 1'b0, 1'b0}), .in_14({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[52:45] , 1'b0}), .in_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[43:36] , 
    1'b0}), .in_16({1'b0, 1'b0, \instanceL2_prod_terms[2][3] [13],  \instanceL2_prod_terms[2][3] [7:1] , 
    layer1_out[27], 1'b0, 1'b0, 1'b0}), .in_17({1'b0, 
    \instanceL2_prod_terms[7][2] [13],  \instanceL2_prod_terms[7][2] [8:7] ,  \instanceL2_prod_terms[8][2] [8:4] , \instanceL2_prod_terms[7][2] [1], 
    layer1_out[18], 1'b0, 1'b0, 1'b0}), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0,  layer1_out[7:0] }), .in_19({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[2][1] [13],  \instanceL2_prod_terms[2][1] [7:1] , 
    layer1_out[9], 1'b0, 1'b0}), .out_0({ \instanceL2_row_sums[3] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_4361 instanceL2_csa_tree_ADD_TC_OP_19_groupi829(
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[178:171] }), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 
    1'b0, 1'b0,  layer1_out[161:153] , 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  \instanceL2_prod_terms[2][16] [11:2] , 
    \instanceL2_prod_terms[0][16][1] , layer1_out[144]}), .in_4({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .in_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[133:126] }), .in_6({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[2][13] [10:1] , 
    layer1_out[117]}), .in_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_8({1'b0, 
    \instanceL2_prod_terms[0][11][13] , \instanceL2_prod_terms[2][11][11] , 
    \instanceL2_prod_terms[2][11][10] , \instanceL2_prod_terms[2][11][9] , 
    \instanceL2_prod_terms[2][11][8] , \instanceL2_prod_terms[2][11][7] , 
    \instanceL2_prod_terms[2][11][6] , \instanceL2_prod_terms[2][11][5] , 
    \instanceL2_prod_terms[2][11][4] , \instanceL2_prod_terms[4][11] [3], 
    \instanceL2_prod_terms[2][11][2] ,  layer1_out[100:99] }), .in_9({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[1][10][10] , \instanceL2_prod_terms[1][10][9] , 
    \instanceL2_prod_terms[1][10][8] , \instanceL2_prod_terms[1][10][7] , 
    \instanceL2_prod_terms[1][10][6] , \instanceL2_prod_terms[1][10][5] , 
    \instanceL2_prod_terms[1][10][4] , \instanceL2_prod_terms[1][10][3] , 
    \instanceL2_prod_terms[1][10][2] ,  layer1_out[91:90] }), .in_10({1'b0, 1'b0, 
    \instanceL2_prod_terms[2][9] [13],  \instanceL2_prod_terms[2][9] [10:3] , layer1_out[81], 1'b0, 1'b0}), .in_11({
    1'b0, 1'b0, \instanceL2_prod_terms[2][8][11] , 
    \instanceL2_prod_terms[2][8][10] , \instanceL2_prod_terms[2][8][9] , 
    \instanceL2_prod_terms[2][8][8] , \instanceL2_prod_terms[2][8][7] , 
    \instanceL2_prod_terms[2][8][6] , \instanceL2_prod_terms[2][8][5] , 
    \instanceL2_prod_terms[2][8][4] , \instanceL2_prod_terms[2][8][3] , 
    \instanceL2_prod_terms[2][8][2] ,  layer1_out[73:72] }), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , 
    layer1_out[63], 1'b0}), .in_13({1'b0, \instanceL2_prod_terms[2][6] [13],  \instanceL2_prod_terms[2][6] [11:3] ,  layer1_out[55:54] , 
    1'b0}), .in_14({1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[9][5] [13],  \instanceL2_prod_terms[2][5] [8:6] , 
    \instanceL2_prod_terms[5][5] [6],  \instanceL2_prod_terms[2][5] [4:2] , layer1_out[45], 1'b0}), .in_15({1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[43:36] , 1'b0}), .in_16({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[2][3] [13],  \instanceL2_prod_terms[2][3] [7:1] , layer1_out[27]}), .in_17({1'b0, 
    \instanceL2_prod_terms[7][2] [13],  \instanceL2_prod_terms[7][2] [8:7] ,  \instanceL2_prod_terms[8][2] [8:4] , \instanceL2_prod_terms[7][2] [1], 
    layer1_out[18], 1'b0, 1'b0, 1'b0}), .in_18({1'b0, 1'b0, 
    \instanceL2_prod_terms[2][0] [13],  \instanceL2_prod_terms[2][0] [10:1] , layer1_out[0]}), .in_19({1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[2][1] [13],  \instanceL2_prod_terms[2][1] [7:1] , layer1_out[9]}),
     .out_0({ \instanceL2_row_sums[2] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_2425 instanceL2_csa_tree_ADD_TC_OP_19_groupi830(
    .in_0({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[1][19] [13],  \instanceL2_prod_terms[1][19] [9:3] , 
    layer1_out[171], 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[169:162] , 1'b0}),
     .in_2({1'b0, 1'b0, \instanceL2_prod_terms[4][17] [13], 
    \instanceL2_prod_terms[0][17][10] , \instanceL2_prod_terms[0][17][9] , 
    \instanceL2_prod_terms[0][17][8] , \instanceL2_prod_terms[0][17][7] , 
    \instanceL2_prod_terms[0][17][6] , \instanceL2_prod_terms[0][17][5] , 
    \instanceL2_prod_terms[0][17][4] , \instanceL2_prod_terms[0][17][3] , 
    \instanceL2_prod_terms[0][17][2] ,  layer1_out[154:153] }), .in_3({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[1][16] [10:3] , 
    \instanceL2_prod_terms[0][16][2] , \instanceL2_prod_terms[0][16][1] , 
    layer1_out[144]}), .in_4({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[1][15] [10:1] , layer1_out[135]}), .in_5({1'b0, 
    \instanceL2_prod_terms[4][14] [13],  \instanceL2_prod_terms[1][14] [11:4] , \instanceL2_prod_terms[0][14][3] , 
    \instanceL2_prod_terms[0][14][2] , \instanceL2_prod_terms[4][14] [1], 
    layer1_out[126]}), .in_6({1'b0, 1'b0, \instanceL2_prod_terms[1][13] [13],  \instanceL2_prod_terms[1][13] [10:1] , 
    layer1_out[117]}), .in_7({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[115:108] , 1'b0, 1'b0}), .in_8({
    1'b0, \instanceL2_prod_terms[1][11] [13],  \instanceL2_prod_terms[1][11] [11:2] , layer1_out[99], 1'b0}), .in_9({
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[1][10][10] , 
    \instanceL2_prod_terms[1][10][9] , \instanceL2_prod_terms[1][10][8] , 
    \instanceL2_prod_terms[1][10][7] , \instanceL2_prod_terms[1][10][6] , 
    \instanceL2_prod_terms[1][10][5] , \instanceL2_prod_terms[1][10][4] , 
    \instanceL2_prod_terms[1][10][3] , \instanceL2_prod_terms[1][10][2] ,  layer1_out[91:90] }),
     .in_10({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[2][9] [13],  \instanceL2_prod_terms[2][9] [10:3] , 
    layer1_out[81], 1'b0}), .in_11({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[1][8][13] , \instanceL2_prod_terms[1][8][9] , 
    \instanceL2_prod_terms[1][8][8] , \instanceL2_prod_terms[1][8][7] , 
    \instanceL2_prod_terms[1][8][6] , \instanceL2_prod_terms[1][8][5] , 
    \instanceL2_prod_terms[1][8][4] , \instanceL2_prod_terms[1][8][3] , 
    \instanceL2_prod_terms[1][8][2] , layer1_out[72], 1'b0}), .in_12({1'b0, 
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , 
    \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , layer1_out[63], 1'b0}), .in_13({ \instanceL2_prod_terms[1][6] [13:1] , 
    layer1_out[54]}), .in_14({1'b0, 1'b0,  \instanceL2_prod_terms[1][5] [11:3] ,  layer1_out[46:45] , 1'b0}), .in_15({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[1][4] [10:2] ,  layer1_out[37:36] }),
     .in_16({1'b0, 1'b0, 1'b0,  \instanceL2_prod_terms[1][3] [10:3] , \instanceL2_prod_terms[0][3][2] ,  layer1_out[28:27] }), .in_17({1'b0, 
    \instanceL2_prod_terms[1][2][12] , \instanceL2_prod_terms[1][2][11] , 
    \instanceL2_prod_terms[1][2][10] , \instanceL2_prod_terms[1][2][9] , 
    \instanceL2_prod_terms[1][2][8] , \instanceL2_prod_terms[1][2][7] , 
    \instanceL2_prod_terms[1][2][6] , \instanceL2_prod_terms[1][2][5] , 
    \instanceL2_prod_terms[1][2][4] , \instanceL2_prod_terms[1][2][3] ,  layer1_out[20:18] }),
     .in_18({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[7:0] , 1'b0, 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[2][1] [13], \instanceL2_prod_terms[1][1][9] , 
    \instanceL2_prod_terms[1][1][8] , \instanceL2_prod_terms[1][1][7] , 
    \instanceL2_prod_terms[1][1][6] , \instanceL2_prod_terms[1][1][5] , 
    \instanceL2_prod_terms[1][1][4] , \instanceL2_prod_terms[1][1][3] , 
    \instanceL2_prod_terms[1][1][2] ,  layer1_out[10:9] }), .out_0({ \instanceL2_row_sums[1] [18:0] }));
  csa_tree_ADD_TC_OP_19_group_2 instanceL2_csa_tree_ADD_TC_OP_19_groupi831(.in_0({
    1'b0, 1'b0, \instanceL2_prod_terms[0][19][13] , 
    \instanceL2_prod_terms[0][19][10] , \instanceL2_prod_terms[0][19][9] , 
    \instanceL2_prod_terms[0][19][8] , \instanceL2_prod_terms[0][19][7] , 
    \instanceL2_prod_terms[0][19][6] , \instanceL2_prod_terms[0][19][5] , 
    \instanceL2_prod_terms[0][19][4] , \instanceL2_prod_terms[0][19][3] , 
    \instanceL2_prod_terms[0][19][2] , \instanceL2_prod_terms[0][19][1] , 
    layer1_out[171]}), .in_1({1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[169:162] , 1'b0, 1'b0}), .in_2({
    1'b0, 1'b0, \instanceL2_prod_terms[4][17] [13], 
    \instanceL2_prod_terms[0][17][10] , \instanceL2_prod_terms[0][17][9] , 
    \instanceL2_prod_terms[0][17][8] , \instanceL2_prod_terms[0][17][7] , 
    \instanceL2_prod_terms[0][17][6] , \instanceL2_prod_terms[0][17][5] , 
    \instanceL2_prod_terms[0][17][4] , \instanceL2_prod_terms[0][17][3] , 
    \instanceL2_prod_terms[0][17][2] ,  layer1_out[154:153] }), .in_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][16][13] , \instanceL2_prod_terms[0][16][7] , 
    \instanceL2_prod_terms[0][16][6] , \instanceL2_prod_terms[0][16][5] , 
    \instanceL2_prod_terms[0][16][4] , \instanceL2_prod_terms[0][16][3] , 
    \instanceL2_prod_terms[0][16][2] , \instanceL2_prod_terms[0][16][1] , 
    layer1_out[144]}), .in_4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[142:135] , 1'b0}), .in_5({
    1'b0, 1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[0][14][9] , 
    \instanceL2_prod_terms[0][14][8] , \instanceL2_prod_terms[0][14][7] , 
    \instanceL2_prod_terms[0][14][6] , \instanceL2_prod_terms[0][14][5] , 
    \instanceL2_prod_terms[0][14][4] , \instanceL2_prod_terms[0][14][3] , 
    \instanceL2_prod_terms[0][14][2] , \instanceL2_prod_terms[4][14] [1], 
    layer1_out[126]}), .in_6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[124:117] }), .in_7({
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[115:108] }), .in_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][11][13] , \instanceL2_prod_terms[0][11][7] , 
    \instanceL2_prod_terms[0][11][6] , \instanceL2_prod_terms[0][11][5] , 
    \instanceL2_prod_terms[0][11][4] , \instanceL2_prod_terms[0][11][3] , 
    \instanceL2_prod_terms[0][11][2] , \instanceL2_prod_terms[0][11][1] , 
    layer1_out[99]}), .in_9({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][10][13] , \instanceL2_prod_terms[0][10][8] , 
    \instanceL2_prod_terms[0][10][7] , \instanceL2_prod_terms[0][10][6] , 
    \instanceL2_prod_terms[0][10][5] , \instanceL2_prod_terms[0][10][4] , 
    \instanceL2_prod_terms[0][10][3] , \instanceL2_prod_terms[0][10][2] , 
    layer1_out[90], 1'b0}), .in_10({\instanceL2_prod_terms[0][9][13] , 
    \instanceL2_prod_terms[0][9][12] , \instanceL2_prod_terms[0][9][11] , 
    \instanceL2_prod_terms[0][9][10] , \instanceL2_prod_terms[0][9][9] , 
    \instanceL2_prod_terms[0][9][8] , \instanceL2_prod_terms[0][9][7] , 
    \instanceL2_prod_terms[0][9][6] , \instanceL2_prod_terms[0][9][5] , 
    \instanceL2_prod_terms[0][9][4] , \instanceL2_prod_terms[0][9][3] , 
    \instanceL2_prod_terms[0][9][2] , \instanceL2_prod_terms[0][9][1] , 
    layer1_out[81]}), .in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_12({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][7] [13],  \instanceL2_prod_terms[0][7] [8:6] , \instanceL2_prod_terms[4][7] [6],  \instanceL2_prod_terms[0][7] [4:2] , 
    layer1_out[63], 1'b0}), .in_13({1'b0, 1'b0, 1'b0, 1'b0, 1'b0,  layer1_out[62:54] }), .in_14({
    1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[9][5] [13], 
    \instanceL2_prod_terms[0][5][9] , \instanceL2_prod_terms[0][5][8] , 
    \instanceL2_prod_terms[0][5][7] , \instanceL2_prod_terms[0][5][6] , 
    \instanceL2_prod_terms[0][5][5] , \instanceL2_prod_terms[0][5][4] , 
    \instanceL2_prod_terms[0][5][3] , \instanceL2_prod_terms[1][5] [3],  layer1_out[46:45] }),
     .in_15({1'b0, 1'b0, \instanceL2_prod_terms[5][4] [13], 
    \instanceL2_prod_terms[0][4][10] , \instanceL2_prod_terms[0][4][9] , 
    \instanceL2_prod_terms[0][4][8] , \instanceL2_prod_terms[0][4][7] , 
    \instanceL2_prod_terms[0][4][6] , \instanceL2_prod_terms[0][4][5] , 
    \instanceL2_prod_terms[0][4][4] , \instanceL2_prod_terms[1][4] [2],  layer1_out[37:36] , 1'b0}),
     .in_16({1'b0, 1'b0, 1'b0, \instanceL2_prod_terms[2][3] [13], 
    \instanceL2_prod_terms[0][3][9] , \instanceL2_prod_terms[0][3][8] , 
    \instanceL2_prod_terms[0][3][7] , \instanceL2_prod_terms[0][3][6] , 
    \instanceL2_prod_terms[0][3][5] , \instanceL2_prod_terms[0][3][4] , 
    \instanceL2_prod_terms[0][3][3] , \instanceL2_prod_terms[0][3][2] ,  layer1_out[28:27] }),
     .in_17({1'b0, 1'b0, \instanceL2_prod_terms[7][2] [13], 
    \instanceL2_prod_terms[0][2][10] , \instanceL2_prod_terms[0][2][9] , 
    \instanceL2_prod_terms[0][2][8] , \instanceL2_prod_terms[0][2][7] , 
    \instanceL2_prod_terms[0][2][6] , \instanceL2_prod_terms[0][2][5] , 
    \instanceL2_prod_terms[0][2][4] , \instanceL2_prod_terms[0][2][3] , 
    \instanceL2_prod_terms[4][2] [3],  layer1_out[19:18] }), .in_18({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[0][0][13] , \instanceL2_prod_terms[0][0][8] , 
    \instanceL2_prod_terms[0][0][7] , \instanceL2_prod_terms[0][0][6] , 
    \instanceL2_prod_terms[0][0][5] , \instanceL2_prod_terms[0][0][4] , 
    \instanceL2_prod_terms[0][0][3] , \instanceL2_prod_terms[0][0][2] , 
    layer1_out[0], 1'b0}), .in_19({1'b0, 1'b0, 1'b0, 1'b0, 
    \instanceL2_prod_terms[9][1] [10], \instanceL2_prod_terms[0][1][8] ,  \instanceL2_prod_terms[9][1] [8:6] , 
    \instanceL2_prod_terms[0][1][4] ,  \instanceL2_prod_terms[9][1] [4:3] , \instanceL2_prod_terms[2][1] [1], 
    layer1_out[9]}), .out_0({ \instanceL2_row_sums[0] [18:0] }));
  csa_tree_SUB_TC_OP_4_group_54 
    \instanceL2_row_iteration[0].prod_calc[9].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[89:81] }), .out_0({
    \instanceL2_prod_terms[0][9][13] , \instanceL2_prod_terms[0][9][12] , 
    \instanceL2_prod_terms[0][9][11] , \instanceL2_prod_terms[0][9][10] , 
    \instanceL2_prod_terms[0][9][9] , \instanceL2_prod_terms[0][9][8] , 
    \instanceL2_prod_terms[0][9][7] , \instanceL2_prod_terms[0][9][6] , 
    \instanceL2_prod_terms[0][9][5] , \instanceL2_prod_terms[0][9][4] , 
    \instanceL2_prod_terms[0][9][3] , \instanceL2_prod_terms[0][9][2] , 
    \instanceL2_prod_terms[0][9][1] , UNCONNECTED375}));
  csa_tree_SUB_TC_OP_4_group_1752 
    \instanceL2_row_iteration[0].prod_calc[19].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[178:171] }), .out_0({
    \instanceL2_prod_terms[0][19][13] , UNCONNECTED378, UNCONNECTED377, 
    \instanceL2_prod_terms[0][19][10] , \instanceL2_prod_terms[0][19][9] , 
    \instanceL2_prod_terms[0][19][8] , \instanceL2_prod_terms[0][19][7] , 
    \instanceL2_prod_terms[0][19][6] , \instanceL2_prod_terms[0][19][5] , 
    \instanceL2_prod_terms[0][19][4] , \instanceL2_prod_terms[0][19][3] , 
    \instanceL2_prod_terms[0][19][2] , \instanceL2_prod_terms[0][19][1] , 
    UNCONNECTED376}));
  csa_tree_SUB_TC_OP_4_group_54_1 
    \instanceL2_row_iteration[1].prod_calc[6].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[62:54] }), .out_0({ \instanceL2_prod_terms[1][6] [13:1] , UNCONNECTED379}));
  csa_tree_SUB_TC_OP_3_group_11408 
    \instanceL2_row_iteration[1].prod_calc[11].mult_inst_csa_tree_SUB_TC_OP_3_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0,  layer1_out[106:99] , 1'b0}), .out_0({
    \instanceL2_prod_terms[1][11] [13], UNCONNECTED382,  \instanceL2_prod_terms[1][11] [11:2] , UNCONNECTED381, 
    UNCONNECTED380}));
  csa_tree_SUB_TC_OP_4_group_1752_1 
    \instanceL2_row_iteration[1].prod_calc[13].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[124:117] }), .out_0({
    \instanceL2_prod_terms[1][13] [13], UNCONNECTED385, UNCONNECTED384,  \instanceL2_prod_terms[1][13] [10:1] , 
    UNCONNECTED383}));
  csa_tree_SUB_TC_OP_4_group_1752_2 
    \instanceL2_row_iteration[2].prod_calc[0].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[7:0] }), .out_0({
    \instanceL2_prod_terms[2][0] [13], UNCONNECTED388, UNCONNECTED387,  \instanceL2_prod_terms[2][0] [10:1] , 
    UNCONNECTED386}));
  csa_tree_SUB_TC_OP_4_group_54_2 
    \instanceL2_row_iteration[3].prod_calc[8].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[80:72] }), .out_0({ \instanceL2_prod_terms[3][8] [13:1] , UNCONNECTED389}));
  csa_tree_SUB_TC_OP_3_group_11408_1 
    \instanceL2_row_iteration[5].prod_calc[17].mult_inst_csa_tree_SUB_TC_OP_3_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0,  layer1_out[161:153] , 1'b0}), .out_0({ \instanceL2_prod_terms[5][17] [13:2] , UNCONNECTED391, 
    UNCONNECTED390}));
  csa_tree_SUB_TC_OP_3_group_11408_2 
    \instanceL2_row_iteration[6].prod_calc[2].mult_inst_csa_tree_SUB_TC_OP_3_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0,  layer1_out[26:18] , 1'b0}), .out_0({ \instanceL2_prod_terms[6][2] [13:2] , UNCONNECTED393, 
    UNCONNECTED392}));
  csa_tree_SUB_TC_OP_3_group_11408_3 
    \instanceL2_row_iteration[6].prod_calc[5].mult_inst_csa_tree_SUB_TC_OP_3_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0,  layer1_out[52:45] , 1'b0}), .out_0({
    \instanceL2_prod_terms[6][5] [13], UNCONNECTED396,  \instanceL2_prod_terms[6][5] [11:2] , UNCONNECTED395, 
    UNCONNECTED394}));
  csa_tree_SUB_TC_OP_4_group_54_3 
    \instanceL2_row_iteration[6].prod_calc[10].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[97:90] }), .out_0({
    \instanceL2_prod_terms[6][10] [13], UNCONNECTED398,  \instanceL2_prod_terms[6][10] [11:1] , UNCONNECTED397}));
  csa_tree_SUB_TC_OP_4_group_54_4 
    \instanceL2_row_iteration[7].prod_calc[3].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[34:27] }), .out_0({
    \instanceL2_prod_terms[7][3] [13], UNCONNECTED400,  \instanceL2_prod_terms[7][3] [11:1] , UNCONNECTED399}));
  csa_tree_SUB_TC_OP_4_group_54_5 
    \instanceL2_row_iteration[7].prod_calc[15].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[142:135] }), .out_0({
    \instanceL2_prod_terms[7][15] [13], UNCONNECTED402,  \instanceL2_prod_terms[7][15] [11:1] , UNCONNECTED401}));
  csa_tree_SUB_TC_OP_4_group_54_6 
    \instanceL2_row_iteration[7].prod_calc[17].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[161:153] }), .out_0({ \instanceL2_prod_terms[7][17] [13:1] , UNCONNECTED403}));
  csa_tree_SUB_TC_OP_4_group_54_7 
    \instanceL2_row_iteration[9].prod_calc[2].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[26:18] }), .out_0({ \instanceL2_prod_terms[9][2] [13:1] , UNCONNECTED404}));
  csa_tree_SUB_TC_OP_4_group_54_8 
    \instanceL2_row_iteration[9].prod_calc[4].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[43:36] }), .out_0({
    \instanceL2_prod_terms[9][4] [13], UNCONNECTED406,  \instanceL2_prod_terms[9][4] [11:1] , UNCONNECTED405}));
  csa_tree_SUB_TC_OP_4_group_1752_3 
    \instanceL2_row_iteration[9].prod_calc[8].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0,  layer1_out[80:72] }), .out_0({
    \instanceL2_prod_terms[9][8] [13], UNCONNECTED408,  \instanceL2_prod_terms[9][8] [11:1] , UNCONNECTED407}));
  csa_tree_SUB_TC_OP_4_group_54_9 
    \instanceL2_row_iteration[9].prod_calc[12].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[115:108] }), .out_0({
    \instanceL2_prod_terms[9][12] [13], UNCONNECTED410,  \instanceL2_prod_terms[9][12] [11:1] , UNCONNECTED409}));
  csa_tree_SUB_TC_OP_4_group_54_10 
    \instanceL2_row_iteration[9].prod_calc[18].mult_inst_csa_tree_SUB_TC_OP_4_groupi (
    .in_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0}), .in_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0}), .in_3({1'b0, 1'b0,  layer1_out[169:162] }), .out_0({
    \instanceL2_prod_terms[9][18] [13], UNCONNECTED412,  \instanceL2_prod_terms[9][18] [11:1] , UNCONNECTED411}));
  SDFFRHQX1 \uut_max_index_reg[0] (.Q(out[0]), .D(n_406), .SE(n_558), .SI(n_510),
     .RN(rst_n), .CK(clk));
  DFFRHQX1 \uut_max_index_reg[1] (.Q(out[1]), .D(n_560), .RN(rst_n), .CK(clk));
  DFFRHQX1 \uut_max_index_reg[2] (.Q(out[2]), .D(n_561), .RN(rst_n), .CK(clk));
  DFFRHQX1 \uut_max_index_reg[3] (.Q(out[3]), .D(n_559), .RN(rst_n), .CK(clk));
  AND2X6 g7059(.Y(out_activehigh[7]), .A(n_565), .B(n_562));
  AND2X6 g7060(.Y(out_activehigh[1]), .A(n_567), .B(n_563));
  AND2X6 g7061(.Y(out_activehigh[0]), .A(n_568), .B(n_563));
  AND2X6 g7062(.Y(out_activehigh[8]), .A(n_564), .B(n_568));
  AND2X6 g7063(.Y(out_activehigh[2]), .A(n_566), .B(n_563));
  AND2X6 g7064(.Y(out_activehigh[6]), .A(n_566), .B(n_562));
  AND2X6 g7065(.Y(out_activehigh[4]), .A(n_562), .B(n_568));
  AND2X6 g7066(.Y(out_activehigh[3]), .A(n_565), .B(n_563));
  AND2X6 g7067(.Y(out_activehigh[5]), .A(n_567), .B(n_562));
  AND2X6 g7068(.Y(out_activehigh[9]), .A(n_564), .B(n_567));
  NOR2X1 g7069(.Y(n_568), .A(out[0]), .B(out[1]));
  NOR2BX1 g7070(.Y(n_567), .AN(out[0]), .B(out[1]));
  NOR2BX1 g7071(.Y(n_566), .AN(out[1]), .B(out[0]));
  AND2X1 g7072(.Y(n_565), .A(out[0]), .B(out[1]));
  NOR2BX1 g7073(.Y(n_564), .AN(out[3]), .B(out[2]));
  NOR2X1 g7075(.Y(n_563), .A(out[2]), .B(out[3]));
  NOR2BX1 g7076(.Y(n_562), .AN(out[2]), .B(out[3]));
  NOR2X1 g7080(.Y(n_561), .A(n_508), .B(n_559));
  NOR2X1 g7081(.Y(n_560), .A(n_509), .B(n_559));
  INVX1 g7082(.Y(n_559), .A(n_558));
  AOI221X1 g7083(.Y(n_558), .A0(n_548), .A1(n_553), .B0(n_555), .B1(n_557), .C0(
    n_556));
  OAI221X1 g7084(.Y(n_557), .A0(n_546), .A1(n_554), .B0(n_543), .B1(n_534), .C0(
    n_552));
  OAI221X1 g7085(.Y(n_556), .A0(n_541), .A1(n_539), .B0(n_536), .B1(n_545), .C0(
    n_84));
  NOR2BX1 g7086(.Y(n_555), .AN(n_548), .B(n_549));
  AOI21X1 g7087(.Y(n_554), .A0(n_412), .A1(n_513), .B0(n_551));
  OAI222X1 g7088(.Y(n_553), .A0(n_411), .A1(n_521), .B0(n_542), .B1(n_538), .C0(
    n_527), .C1(n_528));
  AOI22X1 g7089(.Y(n_552), .A0(n_420), .A1(n_532), .B0(n_524), .B1(n_540));
  INVX1 g7090(.Y(n_551), .A(n_550));
  OAI221X1 g7091(.Y(n_550), .A0(n_413), .A1(n_515), .B0(n_412), .B1(n_513), .C0(
    n_547));
  OAI211X1 g7092(.Y(n_549), .A0(n_425), .A1(n_523), .B0(n_531), .C0(n_537));
  OAI211X1 g7093(.Y(n_547), .A0(n_415), .A1(n_512), .B0(n_526), .C0(n_533));
  OAI211X1 g7094(.Y(n_546), .A0(n_416), .A1(n_516), .B0(n_529), .C0(n_535));
  AOI211XL g7095(.Y(n_548), .A0(n_421), .A1(n_520), .B0(n_530), .C0(n_536));
  INVX1 g7096(.Y(n_545), .A(n_544));
  OAI32X1 g7097(.Y(n_544), .A0(n_421), .A1(n_520), .A2(n_530), .B0(n_423), .B1(
    n_519));
  AOI32X1 g7098(.Y(n_543), .A0(n_416), .A1(n_516), .A2(n_529), .B0(n_417), .B1(
    n_511));
  AOI32X1 g7099(.Y(n_542), .A0(n_425), .A1(n_523), .A2(n_531), .B0(n_422), .B1(
    n_522));
  AOI21X1 g7100(.Y(n_541), .A0(layer2_out[176]), .A1(n_517), .B0(layer2_out[177]));
  OR2XL g7101(.Y(n_540), .A(n_420), .B(n_532));
  AOI31X1 g7102(.Y(n_539), .A0(layer2_out[176]), .A1(layer2_out[177]), .A2(n_517),
     .B0(n_166));
  INVX1 g7103(.Y(n_538), .A(n_537));
  INVX1 g7104(.Y(n_535), .A(n_534));
  OAI2BB1X1 g7105(.Y(n_533), .A0N(n_415), .A1N(n_512), .B0(n_525));
  AOI21X1 g7106(.Y(n_537), .A0(n_424), .A1(n_518), .B0(n_528));
  OAI22X1 g7107(.Y(n_536), .A0(layer2_out[176]), .A1(n_517), .B0(layer2_out[177]),
     .B1(n_166));
  OAI22X1 g7108(.Y(n_534), .A0(n_414), .A1(n_514), .B0(n_420), .B1(n_524));
  AND2X1 g7109(.Y(n_532), .A(n_514), .B(n_414));
  OR2X1 g7110(.Y(n_531), .A(n_422), .B(n_522));
  AND2XL g7111(.Y(n_530), .A(n_423), .B(n_519));
  OR2X1 g7112(.Y(n_529), .A(n_417), .B(n_511));
  OR2XL g7113(.Y(n_527), .A(n_424), .B(n_518));
  NAND2X1 g7114(.Y(n_526), .A(n_413), .B(n_515));
  OAI221X1 g7115(.Y(n_525), .A0(n_435), .A1(n_507), .B0(n_458), .B1(n_508), .C0(
    n_410));
  AND2XL g7116(.Y(n_528), .A(n_411), .B(n_521));
  AOI22X1 g7117(.Y(n_524), .A0(n_461), .A1(n_507), .B0(n_437), .B1(n_508));
  AOI22X1 g7118(.Y(n_523), .A0(n_466), .A1(n_507), .B0(n_447), .B1(n_508));
  AOI22X1 g7119(.Y(n_522), .A0(n_467), .A1(n_507), .B0(n_440), .B1(n_508));
  MX2XL g7120(.Y(n_521), .A(n_439), .B(n_465), .S0(n_507));
  MX2XL g7121(.Y(n_520), .A(n_430), .B(n_453), .S0(n_507));
  MX2XL g7122(.Y(n_519), .A(n_432), .B(n_454), .S0(n_507));
  MX2XL g7123(.Y(n_518), .A(n_444), .B(n_464), .S0(n_507));
  AOI22X1 g7124(.Y(n_517), .A0(n_427), .A1(n_508), .B0(n_459), .B1(n_507));
  AOI22X1 g7125(.Y(n_510), .A0(n_448), .A1(n_507), .B0(n_426), .B1(n_508));
  AOI22X1 g7126(.Y(n_509), .A0(n_418), .A1(n_507), .B0(n_409), .B1(n_508));
  AOI22X1 g7127(.Y(n_516), .A0(n_462), .A1(n_507), .B0(n_446), .B1(n_508));
  AOI22X1 g7128(.Y(n_515), .A0(n_452), .A1(n_507), .B0(n_429), .B1(n_508));
  AOI22X1 g7129(.Y(n_514), .A0(n_463), .A1(n_507), .B0(n_442), .B1(n_508));
  AOI22X1 g7130(.Y(n_513), .A0(n_449), .A1(n_507), .B0(n_431), .B1(n_508));
  MX2XL g7131(.Y(n_512), .A(n_433), .B(n_457), .S0(n_507));
  AOI22X1 g7132(.Y(n_511), .A0(n_455), .A1(n_507), .B0(n_441), .B1(n_508));
  INVX1 g7133(.Y(n_507), .A(n_508));
  OR2X1 g7134(.Y(n_508), .A(n_500), .B(n_506));
  NOR4X1 g7135(.Y(n_506), .A(n_469), .B(n_472), .C(n_488), .D(n_505));
  AOI21X1 g7136(.Y(n_505), .A0(n_499), .A1(n_504), .B0(n_503));
  OAI211X1 g7137(.Y(n_504), .A0(n_462), .A1(n_494), .B0(n_501), .C0(n_502));
  OAI211X1 g7138(.Y(n_503), .A0(n_466), .A1(n_495), .B0(n_491), .C0(n_497));
  OAI211X1 g7139(.Y(n_502), .A0(n_450), .A1(n_431), .B0(n_496), .C0(n_498));
  AOI32X1 g7140(.Y(n_501), .A0(n_456), .A1(n_441), .A2(n_481), .B0(n_485), .B1(
    n_490));
  OAI22X1 g7141(.Y(n_500), .A0(n_488), .A1(n_489), .B0(n_487), .B1(n_486));
  OAI31X1 g7142(.Y(n_499), .A0(n_466), .A1(n_476), .A2(n_483), .B0(n_495));
  OAI31X1 g7143(.Y(n_498), .A0(n_462), .A1(n_474), .A2(n_480), .B0(n_494));
  OAI21X1 g7144(.Y(n_497), .A0(n_439), .A1(n_475), .B0(n_493));
  NAND2X1 g7145(.Y(n_496), .A(n_479), .B(n_492));
  OAI2BB1X1 g7146(.Y(n_493), .A0N(n_439), .A1N(n_475), .B0(n_465));
  NAND3BXL g7147(.Y(n_495), .AN(n_476), .B(n_447), .C(n_482));
  NAND3BXL g7148(.Y(n_494), .AN(n_474), .B(n_446), .C(n_481));
  NAND2X1 g7149(.Y(n_492), .A(n_477), .B(n_478));
  NAND3BXL g7150(.Y(n_491), .AN(n_467), .B(n_440), .C(n_482));
  OAI2BB1X1 g7151(.Y(n_490), .A0N(n_437), .A1N(n_471), .B0(n_461));
  NOR2X1 g7152(.Y(n_489), .A(n_468), .B(n_484));
  NOR2X1 g7153(.Y(n_487), .A(layer2_out[33]), .B(n_473));
  AOI31X1 g7154(.Y(n_486), .A0(layer2_out[33]), .A1(n_460), .A2(n_427), .B0(n_95));
  OR2XL g7155(.Y(n_485), .A(n_437), .B(n_471));
  NOR3BX1 g7156(.Y(n_484), .AN(n_430), .B(n_453), .C(n_472));
  OAI22X1 g7157(.Y(n_488), .A0(n_460), .A1(n_427), .B0(layer2_out[33]), .B1(n_95));
  INVX1 g7158(.Y(n_483), .A(n_482));
  INVX1 g7159(.Y(n_480), .A(n_481));
  AOI22X1 g7160(.Y(n_479), .A0(n_451), .A1(n_429), .B0(n_450), .B1(n_431));
  NAND3BXL g7161(.Y(n_478), .AN(n_435), .B(n_458), .C(n_470));
  AOI22X1 g7162(.Y(n_477), .A0(n_434), .A1(n_457), .B0(n_428), .B1(n_452));
  AOI22X1 g7163(.Y(n_482), .A0(n_445), .A1(n_464), .B0(n_438), .B1(n_465));
  AOI22X1 g7164(.Y(n_481), .A0(n_443), .A1(n_463), .B0(n_436), .B1(n_461));
  AND2XL g7165(.Y(n_473), .A(n_460), .B(n_427));
  NOR2BX1 g7166(.Y(n_476), .AN(n_467), .B(n_440));
  NOR2X1 g7167(.Y(n_475), .A(n_445), .B(n_464));
  NOR2X1 g7168(.Y(n_474), .A(n_456), .B(n_441));
  OR2XL g7169(.Y(n_470), .A(n_434), .B(n_457));
  NOR2BX1 g7170(.Y(n_469), .AN(n_453), .B(n_430));
  NOR2BX1 g7171(.Y(n_468), .AN(n_432), .B(n_454));
  NOR2BX1 g7172(.Y(n_472), .AN(n_454), .B(n_432));
  NOR2X1 g7173(.Y(n_471), .A(n_443), .B(n_463));
  INVX1 g7174(.Y(n_460), .A(n_459));
  OAI22X1 g7175(.Y(n_467), .A0(n_339), .A1(n_419), .B0(n_302), .B1(n_418));
  OAI22X1 g7176(.Y(n_466), .A0(n_333), .A1(n_419), .B0(n_309), .B1(n_418));
  OAI22X1 g7177(.Y(n_465), .A0(n_354), .A1(n_419), .B0(n_287), .B1(n_418));
  OAI22X1 g7178(.Y(n_464), .A0(n_353), .A1(n_419), .B0(n_297), .B1(n_418));
  OAI22X1 g7179(.Y(n_463), .A0(n_342), .A1(n_419), .B0(n_293), .B1(n_418));
  OAI22X1 g7180(.Y(n_462), .A0(n_341), .A1(n_419), .B0(n_290), .B1(n_418));
  OAI22X1 g7181(.Y(n_461), .A0(n_332), .A1(n_419), .B0(n_304), .B1(n_418));
  OAI21X1 g7182(.Y(n_459), .A0(n_124), .A1(n_418), .B0(n_350));
  INVX1 g7183(.Y(n_456), .A(n_455));
  INVX1 g7184(.Y(n_451), .A(n_452));
  INVX1 g7185(.Y(n_450), .A(n_449));
  OAI22X1 g7186(.Y(n_448), .A0(n_307), .A1(n_419), .B0(n_242), .B1(n_418));
  OAI22X1 g7187(.Y(n_458), .A0(n_343), .A1(n_419), .B0(n_313), .B1(n_418));
  OAI22X1 g7188(.Y(n_457), .A0(n_336), .A1(n_419), .B0(n_299), .B1(n_418));
  OAI22X1 g7189(.Y(n_455), .A0(n_340), .A1(n_419), .B0(n_289), .B1(n_418));
  OAI22X1 g7190(.Y(n_454), .A0(n_351), .A1(n_419), .B0(n_295), .B1(n_418));
  OAI22X1 g7191(.Y(n_453), .A0(n_352), .A1(n_419), .B0(n_300), .B1(n_418));
  OAI22X1 g7192(.Y(n_452), .A0(n_338), .A1(n_419), .B0(n_312), .B1(n_418));
  OAI22X1 g7193(.Y(n_449), .A0(n_334), .A1(n_419), .B0(n_291), .B1(n_418));
  INVX1 g7194(.Y(n_445), .A(n_444));
  INVX1 g7195(.Y(n_443), .A(n_442));
  INVX1 g7196(.Y(n_438), .A(n_439));
  INVX1 g7197(.Y(n_436), .A(n_437));
  OAI22X1 g7198(.Y(n_447), .A0(n_283), .A1(n_409), .B0(n_252), .B1(n_408));
  OAI22X1 g7199(.Y(n_446), .A0(n_284), .A1(n_409), .B0(n_248), .B1(n_408));
  OAI22X1 g7200(.Y(n_444), .A0(n_271), .A1(n_409), .B0(n_249), .B1(n_408));
  OAI22X1 g7201(.Y(n_442), .A0(n_273), .A1(n_409), .B0(n_256), .B1(n_408));
  OAI22X1 g7202(.Y(n_441), .A0(n_254), .A1(n_409), .B0(n_247), .B1(n_408));
  OAI22X1 g7203(.Y(n_440), .A0(n_275), .A1(n_409), .B0(n_251), .B1(n_408));
  OAI22X1 g7204(.Y(n_439), .A0(n_272), .A1(n_409), .B0(n_245), .B1(n_408));
  OAI22X1 g7205(.Y(n_437), .A0(n_262), .A1(n_409), .B0(n_246), .B1(n_408));
  INVX1 g7206(.Y(n_434), .A(n_433));
  INVX1 g7207(.Y(n_428), .A(n_429));
  OAI22X1 g7208(.Y(n_426), .A0(n_237), .A1(n_409), .B0(n_239), .B1(n_408));
  OAI22X1 g7209(.Y(n_435), .A0(n_285), .A1(n_409), .B0(n_264), .B1(n_408));
  OAI22X1 g7210(.Y(n_433), .A0(n_276), .A1(n_409), .B0(n_258), .B1(n_408));
  OAI22X1 g7211(.Y(n_432), .A0(n_278), .A1(n_409), .B0(n_253), .B1(n_408));
  OAI22X1 g7212(.Y(n_431), .A0(n_267), .A1(n_409), .B0(n_255), .B1(n_408));
  OAI22X1 g7213(.Y(n_430), .A0(n_269), .A1(n_409), .B0(n_259), .B1(n_408));
  OAI22X1 g7214(.Y(n_429), .A0(n_282), .A1(n_409), .B0(n_260), .B1(n_408));
  OAI22X1 g7215(.Y(n_427), .A0(n_280), .A1(1'b0), .B0(n_96), .B1(n_408));
  INVX1 g7216(.Y(n_418), .A(n_419));
  MX2X1 g7217(.Y(n_425), .A(layer2_out[152]), .B(layer2_out[170]), .S0(n_406));
  AOI22X1 g7218(.Y(n_424), .A0(layer2_out[154]), .A1(n_405), .B0(layer2_out[172]),
     .B1(n_406));
  AOI21X1 g7219(.Y(n_423), .A0(layer2_out[157]), .A1(n_405), .B0(layer2_out[175]));
  MX2XL g7220(.Y(n_422), .A(layer2_out[153]), .B(layer2_out[171]), .S0(n_406));
  AOI22X1 g7221(.Y(n_421), .A0(layer2_out[156]), .A1(n_405), .B0(layer2_out[174]),
     .B1(n_406));
  MX2X1 g7222(.Y(n_420), .A(layer2_out[151]), .B(layer2_out[169]), .S0(n_406));
  OR2X1 g7223(.Y(n_419), .A(n_407), .B(n_403));
  AOI22X1 g7224(.Y(n_410), .A0(layer2_out[144]), .A1(n_405), .B0(layer2_out[162]),
     .B1(n_406));
  MX2XL g7225(.Y(n_417), .A(layer2_out[149]), .B(layer2_out[167]), .S0(n_406));
  MX2X1 g7226(.Y(n_416), .A(layer2_out[148]), .B(layer2_out[166]), .S0(n_406));
  AOI22X1 g7227(.Y(n_415), .A0(layer2_out[145]), .A1(n_405), .B0(layer2_out[163]),
     .B1(n_406));
  MX2XL g7228(.Y(n_414), .A(layer2_out[150]), .B(layer2_out[168]), .S0(n_406));
  MX2X1 g7229(.Y(n_413), .A(layer2_out[164]), .B(layer2_out[146]), .S0(n_405));
  MX2X1 g7230(.Y(n_412), .A(layer2_out[147]), .B(layer2_out[165]), .S0(n_406));
  AOI22X1 g7231(.Y(n_411), .A0(layer2_out[155]), .A1(n_405), .B0(layer2_out[173]),
     .B1(n_406));
  INVX1 g7232(.Y(n_408), .A(n_409));
  OA21X1 g7233(.Y(n_409), .A0(n_349), .A1(n_400), .B0(n_378));
  NOR4X1 g7234(.Y(n_407), .A(n_380), .B(n_379), .C(n_390), .D(n_404));
  INVX1 g7235(.Y(n_405), .A(n_406));
  NAND2X2 g7236(.Y(n_406), .A(n_84), .B(n_401));
  AOI31X1 g7237(.Y(n_404), .A0(n_385), .A1(n_388), .A2(n_395), .B0(n_402));
  OAI221X1 g7238(.Y(n_403), .A0(n_390), .A1(n_398), .B0(n_384), .B1(n_389), .C0(
    n_361));
  NAND2X1 g7239(.Y(n_402), .A(n_387), .B(n_399));
  OAI222X1 g7240(.Y(n_401), .A0(n_181), .A1(n_224), .B0(n_181), .B1(n_392), .C0(
    n_109), .C1(n_199));
  AOI221X1 g7241(.Y(n_400), .A0(n_252), .A1(n_357), .B0(n_365), .B1(n_396), .C0(
    n_381));
  OAI211X1 g7242(.Y(n_399), .A0(n_340), .A1(n_382), .B0(n_383), .C0(n_385));
  INVX1 g7243(.Y(n_398), .A(n_397));
  OAI221X1 g7244(.Y(n_397), .A0(n_379), .A1(n_386), .B0(n_287), .B1(n_371), .C0(
    n_393));
  NAND4XL g7245(.Y(n_396), .A(n_330), .B(n_346), .C(n_362), .D(n_391));
  NAND2X1 g7246(.Y(n_395), .A(n_375), .B(n_394));
  NAND2X1 g7247(.Y(n_394), .A(n_374), .B(n_373));
  OAI2BB1X1 g7248(.Y(n_393), .A0N(n_287), .A1N(n_371), .B0(n_354));
  NAND2X1 g7249(.Y(n_392), .A(n_100), .B(n_377));
  OAI211X1 g7250(.Y(n_391), .A0(n_255), .A1(n_268), .B0(n_360), .C0(n_364));
  AOI32X1 g7251(.Y(n_389), .A0(n_301), .A1(n_352), .A2(n_368), .B0(n_296), .B1(
    n_351));
  NOR2X1 g7252(.Y(n_388), .A(n_358), .B(n_376));
  AOI32X1 g7253(.Y(n_387), .A0(n_294), .A1(n_342), .A2(n_369), .B0(n_305), .B1(
    n_332));
  AOI32X1 g7254(.Y(n_386), .A0(n_310), .A1(n_333), .A2(n_370), .B0(n_303), .B1(
    n_339));
  NAND3BXL g7255(.Y(n_390), .AN(n_384), .B(n_367), .C(n_368));
  NAND2X1 g7256(.Y(n_383), .A(n_289), .B(n_372));
  NOR2X1 g7257(.Y(n_382), .A(n_289), .B(n_372));
  OAI211X1 g7258(.Y(n_381), .A0(n_272), .A1(n_327), .B0(n_326), .C0(n_347));
  OAI21X1 g7259(.Y(n_380), .A0(n_310), .A1(n_333), .B0(n_370));
  OA21X1 g7260(.Y(n_385), .A0(n_294), .A1(n_342), .B0(n_369));
  NAND2X1 g7261(.Y(n_384), .A(n_95), .B(n_366));
  AOI221X1 g7262(.Y(n_378), .A0(n_96), .A1(n_279), .B0(n_315), .B1(n_344), .C0(
    layer2_out[33]));
  AOI221X1 g7263(.Y(n_377), .A0(n_204), .A1(n_321), .B0(layer2_out[170]), .B1(
    n_42), .C0(n_151));
  OAI22X1 g7264(.Y(n_376), .A0(n_292), .A1(n_334), .B0(n_288), .B1(n_340));
  AOI22X1 g7265(.Y(n_375), .A0(n_311), .A1(n_338), .B0(n_292), .B1(n_334));
  AOI22X1 g7266(.Y(n_374), .A0(n_299), .A1(n_335), .B0(n_312), .B1(n_337));
  NAND3BXL g7267(.Y(n_373), .AN(n_343), .B(n_313), .C(n_363));
  OAI22X1 g7268(.Y(n_379), .A0(n_298), .A1(n_353), .B0(n_286), .B1(n_354));
  OR2XL g7269(.Y(n_367), .A(n_301), .B(n_352));
  NAND2BX1 g7270(.Y(n_366), .AN(n_350), .B(n_124));
  NAND2BX1 g7271(.Y(n_372), .AN(n_290), .B(n_341));
  NAND2X1 g7272(.Y(n_371), .A(n_298), .B(n_353));
  OR2XL g7273(.Y(n_370), .A(n_303), .B(n_339));
  OR2XL g7274(.Y(n_369), .A(n_305), .B(n_332));
  OR2XL g7275(.Y(n_368), .A(n_296), .B(n_351));
  INVX1 g7276(.Y(n_365), .A(n_359));
  OAI21X1 g7277(.Y(n_364), .A0(n_325), .A1(n_329), .B0(n_356));
  NAND2BXL g7278(.Y(n_363), .AN(n_299), .B(n_336));
  NAND2XL g7279(.Y(n_362), .A(n_248), .B(n_355));
  NAND3BXL g7280(.Y(n_361), .AN(n_124), .B(n_95), .C(n_350));
  NAND2X1 g7281(.Y(n_360), .A(n_323), .B(n_348));
  AOI31X1 g7282(.Y(n_359), .A0(n_252), .A1(n_316), .A2(n_324), .B0(n_357));
  NOR2BX1 g7283(.Y(n_358), .AN(n_290), .B(n_341));
  INVX1 g7284(.Y(n_357), .A(n_345));
  INVX1 g7285(.Y(n_356), .A(n_355));
  OAI211X1 g7286(.Y(n_349), .A0(n_259), .A1(n_270), .B0(n_315), .C0(n_317));
  NAND2X1 g7287(.Y(n_348), .A(n_322), .B(n_320));
  NAND3BXL g7288(.Y(n_347), .AN(n_275), .B(n_251), .C(n_324));
  NAND3BXL g7289(.Y(n_346), .AN(n_254), .B(n_247), .C(n_328));
  NAND3BXL g7290(.Y(n_345), .AN(n_283), .B(n_316), .C(n_324));
  NOR3X1 g7291(.Y(n_355), .A(n_284), .B(n_319), .C(n_329));
  AOI22X1 g7292(.Y(n_354), .A0(layer2_out[137]), .A1(n_307), .B0(layer2_out[119]),
     .B1(n_308));
  AOI22X1 g7293(.Y(n_353), .A0(layer2_out[136]), .A1(n_307), .B0(layer2_out[118]),
     .B1(n_308));
  AOI22X1 g7294(.Y(n_352), .A0(layer2_out[138]), .A1(n_307), .B0(layer2_out[120]),
     .B1(n_308));
  AOI22X1 g7295(.Y(n_351), .A0(layer2_out[139]), .A1(n_307), .B0(layer2_out[121]),
     .B1(n_308));
  AOI22X1 g7296(.Y(n_350), .A0(layer2_out[140]), .A1(n_307), .B0(layer2_out[122]),
     .B1(n_308));
  INVX1 g7297(.Y(n_344), .A(n_331));
  INVX1 g7298(.Y(n_337), .A(n_338));
  INVX1 g7299(.Y(n_335), .A(n_336));
  AOI32X1 g7300(.Y(n_331), .A0(n_259), .A1(n_270), .A2(n_317), .B0(n_253), .B1(
    n_277));
  AOI32X1 g7301(.Y(n_330), .A0(n_256), .A1(n_274), .A2(n_314), .B0(n_246), .B1(
    n_263));
  AOI22X1 g7302(.Y(n_343), .A0(layer2_out[126]), .A1(n_307), .B0(layer2_out[108]),
     .B1(n_308));
  AOI22X1 g7303(.Y(n_342), .A0(layer2_out[132]), .A1(n_307), .B0(layer2_out[114]),
     .B1(n_308));
  AOI22X1 g7304(.Y(n_341), .A0(layer2_out[130]), .A1(n_307), .B0(layer2_out[112]),
     .B1(n_308));
  AOI22X1 g7305(.Y(n_340), .A0(layer2_out[131]), .A1(n_307), .B0(layer2_out[113]),
     .B1(n_308));
  AOI22X1 g7306(.Y(n_339), .A0(layer2_out[135]), .A1(n_307), .B0(layer2_out[117]),
     .B1(n_308));
  AOI22X1 g7307(.Y(n_338), .A0(layer2_out[128]), .A1(n_307), .B0(layer2_out[110]),
     .B1(n_308));
  AOI22X1 g7308(.Y(n_336), .A0(layer2_out[127]), .A1(n_307), .B0(layer2_out[109]),
     .B1(n_308));
  AOI22X1 g7309(.Y(n_334), .A0(layer2_out[129]), .A1(n_307), .B0(layer2_out[111]),
     .B1(n_308));
  AOI22X1 g7310(.Y(n_333), .A0(layer2_out[134]), .A1(n_307), .B0(layer2_out[116]),
     .B1(n_308));
  AOI22X1 g7311(.Y(n_332), .A0(layer2_out[133]), .A1(n_307), .B0(layer2_out[115]),
     .B1(n_308));
  INVXL g7312(.Y(n_328), .A(n_329));
  NOR2X1 g7313(.Y(n_327), .A(n_245), .B(n_318));
  NAND2X1 g7314(.Y(n_326), .A(n_245), .B(n_318));
  NAND2BXL g7315(.Y(n_325), .AN(n_319), .B(n_248));
  OAI21X1 g7316(.Y(n_329), .A0(n_256), .A1(n_274), .B0(n_314));
  AOI22XL g7317(.Y(n_323), .A0(n_260), .A1(n_281), .B0(n_255), .B1(n_268));
  AOI22X1 g7318(.Y(n_322), .A0(n_276), .A1(n_257), .B0(n_282), .B1(n_261));
  OAI221X1 g7319(.Y(n_321), .A0(layer2_out[151]), .A1(n_11), .B0(layer2_out[150]),
     .B1(n_9), .C0(n_266));
  NAND3BXL g7320(.Y(n_320), .AN(n_264), .B(n_285), .C(n_306));
  AOI22X1 g7321(.Y(n_324), .A0(n_271), .A1(n_250), .B0(n_272), .B1(n_244));
  INVX1 g7322(.Y(n_311), .A(n_312));
  INVX1 g7323(.Y(n_310), .A(n_309));
  INVX1 g7324(.Y(n_307), .A(n_308));
  NAND2BXL g7325(.Y(n_306), .AN(n_276), .B(n_258));
  NOR2BX1 g7326(.Y(n_319), .AN(n_254), .B(n_247));
  NOR2X1 g7327(.Y(n_318), .A(n_271), .B(n_250));
  NAND2BX1 g7328(.Y(n_317), .AN(n_253), .B(n_278));
  NAND2BX1 g7329(.Y(n_316), .AN(n_251), .B(n_275));
  NAND2BX1 g7330(.Y(n_315), .AN(n_96), .B(n_280));
  OR2X1 g7331(.Y(n_314), .A(n_246), .B(n_263));
  AOI22X1 g7332(.Y(n_313), .A0(layer2_out[90]), .A1(n_242), .B0(layer2_out[72]),
     .B1(n_241));
  AOI22X1 g7333(.Y(n_312), .A0(layer2_out[92]), .A1(n_242), .B0(layer2_out[74]),
     .B1(n_241));
  AOI22X1 g7334(.Y(n_309), .A0(layer2_out[98]), .A1(n_242), .B0(layer2_out[80]),
     .B1(n_241));
  OR2X1 g7335(.Y(n_308), .A(n_218), .B(n_265));
  INVX1 g7336(.Y(n_305), .A(n_304));
  INVX1 g7337(.Y(n_303), .A(n_302));
  INVX1 g7338(.Y(n_301), .A(n_300));
  INVX1 g7339(.Y(n_298), .A(n_297));
  INVX1 g7340(.Y(n_296), .A(n_295));
  INVX1 g7341(.Y(n_294), .A(n_293));
  INVX1 g7342(.Y(n_292), .A(n_291));
  INVX1 g7343(.Y(n_288), .A(n_289));
  INVX1 g7344(.Y(n_286), .A(n_287));
  AOI22X1 g7345(.Y(n_304), .A0(layer2_out[97]), .A1(n_242), .B0(layer2_out[79]),
     .B1(n_241));
  AOI22X1 g7346(.Y(n_302), .A0(layer2_out[99]), .A1(n_242), .B0(layer2_out[81]),
     .B1(n_241));
  AOI22X1 g7347(.Y(n_300), .A0(layer2_out[102]), .A1(n_242), .B0(layer2_out[84]),
     .B1(n_241));
  AOI22X1 g7348(.Y(n_299), .A0(layer2_out[91]), .A1(n_242), .B0(layer2_out[73]),
     .B1(n_241));
  AOI22X1 g7349(.Y(n_297), .A0(layer2_out[100]), .A1(n_242), .B0(layer2_out[82]),
     .B1(n_241));
  AOI22X1 g7350(.Y(n_295), .A0(layer2_out[103]), .A1(n_242), .B0(layer2_out[85]),
     .B1(n_241));
  AOI22X1 g7351(.Y(n_293), .A0(layer2_out[96]), .A1(n_242), .B0(layer2_out[78]),
     .B1(n_241));
  AOI22X1 g7352(.Y(n_291), .A0(layer2_out[93]), .A1(n_242), .B0(layer2_out[75]),
     .B1(n_241));
  AOI22X1 g7353(.Y(n_290), .A0(layer2_out[94]), .A1(n_242), .B0(layer2_out[76]),
     .B1(n_241));
  AOI22X1 g7354(.Y(n_289), .A0(layer2_out[95]), .A1(n_242), .B0(layer2_out[77]),
     .B1(n_241));
  AOI22X1 g7355(.Y(n_287), .A0(layer2_out[101]), .A1(n_242), .B0(layer2_out[83]),
     .B1(n_241));
  INVX1 g7356(.Y(n_281), .A(n_282));
  INVX1 g7357(.Y(n_279), .A(n_280));
  INVX1 g7358(.Y(n_277), .A(n_278));
  INVX1 g7359(.Y(n_274), .A(n_273));
  INVX1 g7360(.Y(n_270), .A(n_269));
  INVX1 g7361(.Y(n_268), .A(n_267));
  OAI21X1 g7362(.Y(n_266), .A0(layer2_out[167]), .A1(n_232), .B0(n_243));
  NOR4X1 g7363(.Y(n_265), .A(n_119), .B(n_135), .C(n_152), .D(n_240));
  AOI22X1 g7364(.Y(n_285), .A0(layer2_out[18]), .A1(n_237), .B0(layer2_out[0]),
     .B1(n_236));
  AOI22X1 g7365(.Y(n_284), .A0(layer2_out[22]), .A1(n_237), .B0(layer2_out[4]),
     .B1(n_236));
  AOI22X1 g7366(.Y(n_283), .A0(layer2_out[26]), .A1(n_237), .B0(layer2_out[8]),
     .B1(n_236));
  AOI22X1 g7367(.Y(n_282), .A0(layer2_out[20]), .A1(n_237), .B0(layer2_out[2]),
     .B1(n_236));
  AOI21X1 g7368(.Y(n_280), .A0(layer2_out[14]), .A1(n_236), .B0(layer2_out[32]));
  AOI22X1 g7369(.Y(n_278), .A0(layer2_out[31]), .A1(n_237), .B0(layer2_out[13]),
     .B1(n_236));
  AOI22X1 g7370(.Y(n_276), .A0(layer2_out[19]), .A1(n_237), .B0(layer2_out[1]),
     .B1(n_236));
  AOI22X1 g7371(.Y(n_275), .A0(layer2_out[27]), .A1(n_237), .B0(layer2_out[9]),
     .B1(n_236));
  AOI22X1 g7372(.Y(n_273), .A0(layer2_out[24]), .A1(n_237), .B0(layer2_out[6]),
     .B1(n_236));
  AOI22X1 g7373(.Y(n_272), .A0(layer2_out[29]), .A1(n_237), .B0(layer2_out[11]),
     .B1(n_236));
  AOI22X1 g7374(.Y(n_271), .A0(layer2_out[28]), .A1(n_237), .B0(layer2_out[10]),
     .B1(n_236));
  AOI22X1 g7375(.Y(n_269), .A0(layer2_out[30]), .A1(n_237), .B0(layer2_out[12]),
     .B1(n_236));
  AOI22X1 g7376(.Y(n_267), .A0(layer2_out[21]), .A1(n_237), .B0(layer2_out[3]),
     .B1(n_236));
  INVX1 g7377(.Y(n_263), .A(n_262));
  INVX1 g7378(.Y(n_261), .A(n_260));
  INVX1 g7379(.Y(n_257), .A(n_258));
  INVX1 g7380(.Y(n_250), .A(n_249));
  INVX1 g7381(.Y(n_244), .A(n_245));
  AOI22X1 g7382(.Y(n_264), .A0(layer2_out[54]), .A1(n_239), .B0(layer2_out[36]),
     .B1(n_238));
  AOI22X1 g7383(.Y(n_262), .A0(layer2_out[25]), .A1(n_237), .B0(layer2_out[7]),
     .B1(n_236));
  AOI22X1 g7384(.Y(n_260), .A0(layer2_out[56]), .A1(n_239), .B0(layer2_out[38]),
     .B1(n_238));
  AOI22X1 g7385(.Y(n_259), .A0(layer2_out[66]), .A1(n_239), .B0(layer2_out[48]),
     .B1(n_238));
  AOI22X1 g7386(.Y(n_258), .A0(layer2_out[55]), .A1(n_239), .B0(layer2_out[37]),
     .B1(n_238));
  AOI22X1 g7387(.Y(n_256), .A0(layer2_out[60]), .A1(n_239), .B0(layer2_out[42]),
     .B1(n_238));
  AOI22X1 g7388(.Y(n_255), .A0(layer2_out[57]), .A1(n_239), .B0(layer2_out[39]),
     .B1(n_238));
  AOI22X1 g7389(.Y(n_254), .A0(layer2_out[23]), .A1(n_237), .B0(layer2_out[5]),
     .B1(n_236));
  AOI22X1 g7390(.Y(n_253), .A0(layer2_out[67]), .A1(n_239), .B0(layer2_out[49]),
     .B1(n_238));
  AOI22X1 g7391(.Y(n_252), .A0(layer2_out[62]), .A1(n_239), .B0(layer2_out[44]),
     .B1(n_238));
  AOI22X1 g7392(.Y(n_251), .A0(layer2_out[63]), .A1(n_239), .B0(layer2_out[45]),
     .B1(n_238));
  AOI22X1 g7393(.Y(n_249), .A0(layer2_out[64]), .A1(n_239), .B0(layer2_out[46]),
     .B1(n_238));
  AOI22X1 g7394(.Y(n_248), .A0(layer2_out[58]), .A1(n_239), .B0(layer2_out[40]),
     .B1(n_238));
  AOI22X1 g7395(.Y(n_247), .A0(layer2_out[59]), .A1(n_239), .B0(layer2_out[41]),
     .B1(n_238));
  AOI22X1 g7396(.Y(n_246), .A0(layer2_out[61]), .A1(n_239), .B0(layer2_out[43]),
     .B1(n_238));
  AOI22X1 g7397(.Y(n_245), .A0(layer2_out[65]), .A1(n_239), .B0(layer2_out[47]),
     .B1(n_238));
  OAI2BB1X1 g7398(.Y(n_243), .A0N(layer2_out[167]), .A1N(n_232), .B0(
    layer2_out[149]));
  INVX1 g7399(.Y(n_241), .A(n_242));
  AOI21X1 g7400(.Y(n_240), .A0(n_211), .A1(n_233), .B0(n_222));
  AND2X1 g7401(.Y(n_242), .A(n_4), .B(n_235));
  INVX1 g7402(.Y(n_238), .A(n_239));
  INVX1 g7403(.Y(n_236), .A(n_237));
  AOI21X2 g7404(.Y(n_239), .A0(n_213), .A1(n_223), .B0(n_230));
  AND4X1 g7405(.Y(n_237), .A(n_143), .B(n_206), .C(n_227), .D(n_231));
  AOI222X1 g7407(.Y(n_235), .A0(n_134), .A1(n_191), .B0(layer2_out[86]), .B1(
    n_51), .C0(n_179), .C1(n_228));
  OAI211X1 g7408(.Y(n_234), .A0(layer2_out[94]), .A1(n_195), .B0(n_214), .C0(
    n_229));
  OAI211X1 g7409(.Y(n_233), .A0(layer2_out[130]), .A1(n_194), .B0(n_221), .C0(
    n_226));
  NAND2X1 g7410(.Y(n_231), .A(n_209), .B(n_225));
  OAI222X1 g7411(.Y(n_230), .A0(n_131), .A1(n_177), .B0(n_178), .B1(n_216), .C0(
    layer2_out[68]), .C1(n_35));
  AOI32X1 g7412(.Y(n_232), .A0(n_116), .A1(n_88), .A2(n_220), .B0(
    layer2_out[148]), .B1(n_30));
  OAI211X1 g7413(.Y(n_229), .A0(layer2_out[75]), .A1(n_16), .B0(n_203), .C0(
    n_212));
  OAI222X1 g7414(.Y(n_228), .A0(n_156), .A1(n_186), .B0(layer2_out[98]), .B1(
    n_192), .C0(n_114), .C1(n_149));
  NAND2BX1 g7415(.Y(n_227), .AN(n_180), .B(n_215));
  OAI211X1 g7416(.Y(n_226), .A0(layer2_out[111]), .A1(n_59), .B0(n_201), .C0(
    n_210));
  OAI211X1 g7417(.Y(n_225), .A0(n_164), .A1(n_172), .B0(n_173), .C0(n_219));
  OA22X1 g7418(.Y(n_224), .A0(n_151), .A1(n_198), .B0(n_158), .B1(n_188));
  NAND4XL g7419(.Y(n_223), .A(n_93), .B(n_142), .C(n_197), .D(n_217));
  OAI222X1 g7420(.Y(n_222), .A0(n_159), .A1(n_190), .B0(layer2_out[134]), .B1(
    n_193), .C0(n_115), .C1(n_145));
  AOI31X1 g7421(.Y(n_221), .A0(layer2_out[113]), .A1(n_61), .A2(n_147), .B0(
    n_205));
  OAI221X1 g7422(.Y(n_220), .A0(layer2_out[164]), .A1(n_27), .B0(layer2_out[165]),
     .B1(n_56), .C0(n_196));
  NAND3BXL g7423(.Y(n_219), .AN(n_164), .B(n_169), .C(n_200));
  OAI222X1 g7424(.Y(n_218), .A0(n_121), .A1(n_132), .B0(n_152), .B1(n_176), .C0(
    layer2_out[141]), .C1(n_25));
  NAND3BXL g7425(.Y(n_217), .AN(n_168), .B(n_163), .C(n_202));
  AOI21X1 g7426(.Y(n_216), .A0(n_150), .A1(n_175), .B0(n_207));
  OAI222X1 g7427(.Y(n_215), .A0(n_118), .A1(n_127), .B0(n_153), .B1(n_171), .C0(
    layer2_out[29]), .C1(n_31));
  AOI31X1 g7428(.Y(n_214), .A0(layer2_out[77]), .A1(n_55), .A2(n_162), .B0(n_170));
  NOR2X1 g7429(.Y(n_213), .A(n_167), .B(n_178));
  OAI31X1 g7430(.Y(n_212), .A0(layer2_out[94]), .A1(n_129), .A2(n_161), .B0(
    n_195));
  OAI31X1 g7431(.Y(n_211), .A0(layer2_out[134]), .A1(n_128), .A2(n_145), .B0(
    n_193));
  OAI31X1 g7432(.Y(n_210), .A0(layer2_out[130]), .A1(n_102), .A2(n_146), .B0(
    n_194));
  NOR4X1 g7433(.Y(n_209), .A(n_92), .B(n_97), .C(n_153), .D(n_180));
  OAI31X1 g7434(.Y(n_208), .A0(layer2_out[98]), .A1(n_112), .A2(n_149), .B0(
    n_192));
  AOI21XL g7435(.Y(n_207), .A0(layer2_out[65]), .A1(n_120), .B0(n_187));
  NAND2X1 g7436(.Y(n_206), .A(n_165), .B(n_174));
  AOI21XL g7437(.Y(n_205), .A0(layer2_out[133]), .A1(n_117), .B0(n_189));
  OAI22X1 g7438(.Y(n_204), .A0(layer2_out[151]), .A1(n_160), .B0(n_11), .B1(n_94));
  OAI221X1 g7439(.Y(n_203), .A0(layer2_out[92]), .A1(n_21), .B0(layer2_out[93]),
     .B1(n_62), .C0(n_182));
  OAI221X1 g7440(.Y(n_202), .A0(layer2_out[56]), .A1(n_50), .B0(layer2_out[57]),
     .B1(n_67), .C0(n_183));
  OAI221X1 g7441(.Y(n_201), .A0(layer2_out[128]), .A1(n_72), .B0(layer2_out[129]),
     .B1(n_52), .C0(n_184));
  OAI221X1 g7442(.Y(n_200), .A0(layer2_out[20]), .A1(n_19), .B0(layer2_out[21]),
     .B1(n_23), .C0(n_185));
  AOI32X1 g7443(.Y(n_199), .A0(layer2_out[156]), .A1(n_79), .A2(n_107), .B0(
    layer2_out[157]), .B1(n_73));
  AOI32X1 g7444(.Y(n_198), .A0(layer2_out[152]), .A1(n_64), .A2(n_100), .B0(
    layer2_out[153]), .B1(n_33));
  OAI211X1 g7445(.Y(n_197), .A0(layer2_out[41]), .A1(n_155), .B0(n_163), .C0(
    n_154));
  OAI222X1 g7446(.Y(n_196), .A0(layer2_out[145]), .A1(n_70), .B0(layer2_out[144]),
     .B1(n_157), .C0(layer2_out[146]), .C1(n_58));
  OAI32X1 g7447(.Y(n_191), .A0(layer2_out[102]), .A1(n_54), .A2(n_137), .B0(
    layer2_out[103]), .B1(n_74));
  AOI21X1 g7448(.Y(n_190), .A0(layer2_out[118]), .A1(n_89), .B0(layer2_out[119]));
  AOI21XL g7449(.Y(n_189), .A0(layer2_out[114]), .A1(n_113), .B0(layer2_out[115]));
  AOI21XL g7450(.Y(n_188), .A0(layer2_out[154]), .A1(n_123), .B0(layer2_out[155]));
  AOI21XL g7451(.Y(n_187), .A0(layer2_out[46]), .A1(n_90), .B0(layer2_out[47]));
  AOI21X1 g7452(.Y(n_186), .A0(layer2_out[82]), .A1(n_86), .B0(layer2_out[83]));
  OAI221X1 g7453(.Y(n_185), .A0(layer2_out[1]), .A1(n_60), .B0(layer2_out[2]),
     .B1(n_15), .C0(n_141));
  OAI221X1 g7454(.Y(n_184), .A0(layer2_out[109]), .A1(n_75), .B0(layer2_out[110]),
     .B1(n_57), .C0(n_138));
  OAI221X1 g7455(.Y(n_183), .A0(layer2_out[37]), .A1(n_68), .B0(layer2_out[38]),
     .B1(n_22), .C0(n_139));
  OAI221X1 g7456(.Y(n_182), .A0(layer2_out[73]), .A1(n_77), .B0(layer2_out[74]),
     .B1(n_69), .C0(n_140));
  NAND3BXL g7457(.Y(n_195), .AN(n_129), .B(layer2_out[76]), .C(n_162));
  NAND3BXL g7458(.Y(n_194), .AN(n_102), .B(layer2_out[112]), .C(n_147));
  NAND3BXL g7459(.Y(n_193), .AN(n_128), .B(layer2_out[116]), .C(n_144));
  NAND3BXL g7460(.Y(n_192), .AN(n_112), .B(layer2_out[80]), .C(n_148));
  AOI32X1 g7462(.Y(n_177), .A0(layer2_out[48]), .A1(n_71), .A2(n_99), .B0(
    layer2_out[49]), .B1(n_37));
  AOI32X1 g7463(.Y(n_176), .A0(layer2_out[120]), .A1(n_44), .A2(n_136), .B0(
    layer2_out[121]), .B1(n_14));
  OAI32X1 g7464(.Y(n_175), .A0(layer2_out[62]), .A1(n_65), .A2(n_104), .B0(
    layer2_out[63]), .B1(n_28));
  OAI32X1 g7465(.Y(n_174), .A0(layer2_out[30]), .A1(n_66), .A2(n_111), .B0(
    layer2_out[31]), .B1(n_39));
  AOI32X1 g7466(.Y(n_173), .A0(layer2_out[6]), .A1(n_81), .A2(n_101), .B0(
    layer2_out[7]), .B1(n_18));
  AOI32X1 g7467(.Y(n_172), .A0(layer2_out[4]), .A1(n_47), .A2(n_106), .B0(
    layer2_out[5]), .B1(n_38));
  AOI32X1 g7468(.Y(n_171), .A0(layer2_out[8]), .A1(n_80), .A2(n_98), .B0(
    layer2_out[9]), .B1(n_17));
  OAI32X1 g7469(.Y(n_170), .A0(layer2_out[96]), .A1(n_53), .A2(n_126), .B0(
    layer2_out[97]), .B1(n_49));
  AOI221X1 g7470(.Y(n_169), .A0(layer2_out[21]), .A1(n_23), .B0(layer2_out[22]),
     .B1(n_26), .C0(n_105));
  OAI222X1 g7471(.Y(n_168), .A0(layer2_out[39]), .A1(n_41), .B0(layer2_out[41]),
     .B1(n_10), .C0(layer2_out[40]), .C1(n_13));
  OAI211X1 g7472(.Y(n_167), .A0(layer2_out[44]), .A1(n_29), .B0(n_103), .C0(
    n_150));
  OAI211X1 g7473(.Y(n_181), .A0(layer2_out[156]), .A1(n_79), .B0(n_108), .C0(
    n_107));
  OAI211X1 g7474(.Y(n_180), .A0(layer2_out[12]), .A1(n_43), .B0(n_110), .C0(
    n_165));
  AOI211XL g7475(.Y(n_179), .A0(layer2_out[102]), .A1(n_54), .B0(n_137), .C0(
    n_133));
  OAI211X1 g7476(.Y(n_178), .A0(layer2_out[48]), .A1(n_71), .B0(n_130), .C0(n_99));
  INVX1 g7477(.Y(n_161), .A(n_162));
  NOR3BX1 g7478(.Y(n_160), .AN(layer2_out[150]), .B(layer2_out[168]), .C(
    layer2_out[169]));
  OA21X1 g7479(.Y(n_159), .A0(layer2_out[136]), .A1(n_6), .B0(layer2_out[137]));
  OA21X1 g7480(.Y(n_158), .A0(layer2_out[172]), .A1(n_12), .B0(layer2_out[173]));
  OAI2BB1X1 g7481(.Y(n_157), .A0N(layer2_out[145]), .A1N(n_70), .B0(
    layer2_out[162]));
  OA21X1 g7482(.Y(n_156), .A0(layer2_out[100]), .A1(n_46), .B0(layer2_out[101]));
  NOR3BX1 g7483(.Y(n_155), .AN(layer2_out[40]), .B(layer2_out[59]), .C(
    layer2_out[58]));
  OAI2BB1X1 g7484(.Y(n_154), .A0N(layer2_out[40]), .A1N(n_13), .B0(
    layer2_out[59]));
  NOR2BX1 g7485(.Y(n_166), .AN(n_95), .B(layer2_out[33]));
  AOI21X1 g7486(.Y(n_165), .A0(layer2_out[32]), .A1(n_20), .B0(layer2_out[33]));
  OAI21X1 g7487(.Y(n_164), .A0(layer2_out[6]), .A1(n_81), .B0(n_101));
  AOI21X1 g7488(.Y(n_163), .A0(layer2_out[60]), .A1(n_78), .B0(n_125));
  AOI21X1 g7489(.Y(n_162), .A0(layer2_out[96]), .A1(n_53), .B0(n_126));
  INVX1 g7490(.Y(n_149), .A(n_148));
  INVX1 g7491(.Y(n_146), .A(n_147));
  INVX1 g7492(.Y(n_145), .A(n_144));
  NAND3BXL g7493(.Y(n_143), .AN(layer2_out[32]), .B(layer2_out[14]), .C(n_5));
  OR3XL g7494(.Y(n_142), .A(layer2_out[60]), .B(n_78), .C(n_125));
  OAI211X1 g7495(.Y(n_141), .A0(layer2_out[19]), .A1(n_24), .B0(layer2_out[18]),
     .C0(n_85));
  OAI211X1 g7496(.Y(n_140), .A0(layer2_out[91]), .A1(n_48), .B0(layer2_out[90]),
     .C0(n_82));
  OAI211X1 g7497(.Y(n_139), .A0(layer2_out[55]), .A1(n_63), .B0(layer2_out[54]),
     .C0(n_45));
  OAI211X1 g7498(.Y(n_138), .A0(layer2_out[127]), .A1(n_40), .B0(layer2_out[126]),
     .C0(n_83));
  NAND2BX1 g7499(.Y(n_153), .AN(n_127), .B(n_87));
  NAND2BX1 g7500(.Y(n_152), .AN(n_132), .B(n_122));
  OAI2BB1X1 g7501(.Y(n_151), .A0N(layer2_out[172]), .A1N(n_12), .B0(n_91));
  AOI22X1 g7502(.Y(n_150), .A0(layer2_out[64]), .A1(n_8), .B0(layer2_out[65]),
     .B1(n_76));
  AOI22X1 g7503(.Y(n_148), .A0(layer2_out[100]), .A1(n_46), .B0(layer2_out[101]),
     .B1(n_34));
  AOI22X1 g7504(.Y(n_147), .A0(layer2_out[132]), .A1(n_7), .B0(layer2_out[133]),
     .B1(n_36));
  AOI22X1 g7505(.Y(n_144), .A0(layer2_out[136]), .A1(n_6), .B0(layer2_out[137]),
     .B1(n_32));
  INVX1 g7506(.Y(n_136), .A(n_135));
  INVX1 g7507(.Y(n_134), .A(n_133));
  INVX1 g7508(.Y(n_131), .A(n_130));
  NOR2XL g7509(.Y(n_123), .A(layer2_out[173]), .B(layer2_out[172]));
  NAND2BX1 g7510(.Y(n_122), .AN(layer2_out[122]), .B(layer2_out[140]));
  NAND2BXL g7511(.Y(n_121), .AN(layer2_out[140]), .B(layer2_out[122]));
  NAND2BXL g7512(.Y(n_120), .AN(layer2_out[64]), .B(layer2_out[46]));
  NOR2X1 g7513(.Y(n_119), .A(layer2_out[120]), .B(n_44));
  NAND2BXL g7514(.Y(n_118), .AN(layer2_out[28]), .B(layer2_out[10]));
  NAND2BXL g7515(.Y(n_117), .AN(layer2_out[132]), .B(layer2_out[114]));
  NAND2XL g7516(.Y(n_116), .A(layer2_out[165]), .B(n_56));
  NAND2BXL g7517(.Y(n_115), .AN(layer2_out[135]), .B(layer2_out[117]));
  NAND2BXL g7518(.Y(n_114), .AN(layer2_out[99]), .B(layer2_out[81]));
  NOR2XL g7519(.Y(n_113), .A(layer2_out[133]), .B(layer2_out[132]));
  NOR2BX1 g7520(.Y(n_137), .AN(layer2_out[103]), .B(layer2_out[85]));
  NOR2X1 g7521(.Y(n_135), .A(layer2_out[121]), .B(n_14));
  NOR2X1 g7522(.Y(n_133), .A(layer2_out[86]), .B(n_51));
  NOR2BX1 g7523(.Y(n_132), .AN(layer2_out[141]), .B(layer2_out[123]));
  NAND2X1 g7524(.Y(n_130), .A(layer2_out[68]), .B(n_35));
  NOR2X1 g7525(.Y(n_129), .A(layer2_out[77]), .B(n_55));
  NOR2BX1 g7526(.Y(n_128), .AN(layer2_out[135]), .B(layer2_out[117]));
  NOR2BX1 g7527(.Y(n_127), .AN(layer2_out[29]), .B(layer2_out[11]));
  AND2X1 g7528(.Y(n_126), .A(n_49), .B(layer2_out[97]));
  NOR2BX1 g7529(.Y(n_125), .AN(layer2_out[61]), .B(layer2_out[43]));
  NOR2X1 g7530(.Y(n_124), .A(layer2_out[86]), .B(layer2_out[104]));
  INVX1 g7531(.Y(n_111), .A(n_110));
  INVX1 g7532(.Y(n_109), .A(n_108));
  INVX1 g7533(.Y(n_106), .A(n_105));
  INVX1 g7534(.Y(n_104), .A(n_103));
  INVX1 g7535(.Y(n_98), .A(n_97));
  NOR2BX1 g7536(.Y(n_94), .AN(layer2_out[150]), .B(layer2_out[168]));
  NAND2BXL g7537(.Y(n_93), .AN(layer2_out[61]), .B(layer2_out[43]));
  NOR2X1 g7538(.Y(n_92), .A(layer2_out[8]), .B(n_80));
  NAND2BX1 g7539(.Y(n_91), .AN(layer2_out[155]), .B(layer2_out[173]));
  NOR2XL g7540(.Y(n_90), .A(layer2_out[65]), .B(layer2_out[64]));
  NOR2X1 g7541(.Y(n_89), .A(layer2_out[136]), .B(layer2_out[137]));
  NAND2BXL g7542(.Y(n_88), .AN(layer2_out[148]), .B(layer2_out[166]));
  NAND2BX1 g7543(.Y(n_87), .AN(layer2_out[10]), .B(layer2_out[28]));
  NOR2X1 g7544(.Y(n_86), .A(layer2_out[100]), .B(layer2_out[101]));
  NOR2BX1 g7545(.Y(n_112), .AN(layer2_out[99]), .B(layer2_out[81]));
  NAND2X1 g7546(.Y(n_110), .A(layer2_out[31]), .B(n_39));
  NOR2X1 g7547(.Y(n_108), .A(layer2_out[176]), .B(layer2_out[177]));
  OR2X1 g7548(.Y(n_107), .A(layer2_out[157]), .B(n_73));
  NOR2X1 g7549(.Y(n_105), .A(layer2_out[5]), .B(n_38));
  NAND2X1 g7550(.Y(n_103), .A(layer2_out[63]), .B(n_28));
  NOR2X1 g7551(.Y(n_102), .A(layer2_out[113]), .B(n_61));
  OR2X1 g7552(.Y(n_101), .A(layer2_out[7]), .B(n_18));
  OR2X1 g7553(.Y(n_100), .A(layer2_out[153]), .B(n_33));
  OR2XL g7554(.Y(n_99), .A(layer2_out[49]), .B(n_37));
  NOR2X1 g7555(.Y(n_97), .A(layer2_out[9]), .B(n_17));
  NOR2X1 g7556(.Y(n_96), .A(layer2_out[50]), .B(layer2_out[68]));
  NOR2X1 g7557(.Y(n_95), .A(layer2_out[123]), .B(layer2_out[141]));
  INVX1 g7558(.Y(n_85), .A(layer2_out[0]));
  INVX1 g7559(.Y(n_84), .A(layer2_out[178]));
  INVX1 g7560(.Y(n_83), .A(layer2_out[108]));
  INVX1 g7561(.Y(n_82), .A(layer2_out[72]));
  INVX1 g7562(.Y(n_81), .A(layer2_out[24]));
  INVX1 g7563(.Y(n_80), .A(layer2_out[26]));
  INVX1 g7564(.Y(n_79), .A(layer2_out[174]));
  INVX1 g7565(.Y(n_78), .A(layer2_out[42]));
  INVX1 g7566(.Y(n_77), .A(layer2_out[91]));
  INVX1 g7567(.Y(n_76), .A(layer2_out[47]));
  INVX1 g7568(.Y(n_75), .A(layer2_out[127]));
  INVX1 g7569(.Y(n_74), .A(layer2_out[85]));
  INVX1 g7570(.Y(n_73), .A(layer2_out[175]));
  INVX1 g7571(.Y(n_72), .A(layer2_out[110]));
  INVX1 g7572(.Y(n_71), .A(layer2_out[66]));
  INVX1 g7573(.Y(n_70), .A(layer2_out[163]));
  INVX1 g7574(.Y(n_69), .A(layer2_out[92]));
  INVX1 g7575(.Y(n_68), .A(layer2_out[55]));
  INVX1 g7576(.Y(n_67), .A(layer2_out[39]));
  INVX1 g7577(.Y(n_66), .A(layer2_out[12]));
  INVX1 g7578(.Y(n_65), .A(layer2_out[44]));
  INVX1 g7579(.Y(n_64), .A(layer2_out[170]));
  INVX1 g7580(.Y(n_63), .A(layer2_out[37]));
  INVX1 g7581(.Y(n_62), .A(layer2_out[75]));
  INVX1 g7582(.Y(n_61), .A(layer2_out[131]));
  INVX1 g7583(.Y(n_60), .A(layer2_out[19]));
  INVX1 g7584(.Y(n_59), .A(layer2_out[129]));
  INVX1 g7585(.Y(n_58), .A(layer2_out[164]));
  INVX1 g7586(.Y(n_57), .A(layer2_out[128]));
  INVX1 g7587(.Y(n_56), .A(layer2_out[147]));
  INVX1 g7588(.Y(n_55), .A(layer2_out[95]));
  INVX1 g7589(.Y(n_54), .A(layer2_out[84]));
  INVX1 g7590(.Y(n_53), .A(layer2_out[78]));
  INVX1 g7591(.Y(n_52), .A(layer2_out[111]));
  INVX1 g7592(.Y(n_51), .A(layer2_out[104]));
  INVX1 g7593(.Y(n_50), .A(layer2_out[38]));
  INVX1 g7594(.Y(n_49), .A(layer2_out[79]));
  INVX1 g7595(.Y(n_48), .A(layer2_out[73]));
  INVX1 g7596(.Y(n_47), .A(layer2_out[22]));
  INVX1 g7597(.Y(n_46), .A(layer2_out[82]));
  INVX1 g7598(.Y(n_45), .A(layer2_out[36]));
  INVX1 g7599(.Y(n_44), .A(layer2_out[138]));
  INVX1 g7600(.Y(n_43), .A(layer2_out[30]));
  INVX1 g7601(.Y(n_42), .A(layer2_out[152]));
  INVX1 g7602(.Y(n_41), .A(layer2_out[57]));
  INVX1 g7603(.Y(n_40), .A(layer2_out[109]));
  INVX1 g7604(.Y(n_39), .A(layer2_out[13]));
  INVX1 g7605(.Y(n_38), .A(layer2_out[23]));
  INVX1 g7606(.Y(n_37), .A(layer2_out[67]));
  INVX1 g7607(.Y(n_36), .A(layer2_out[115]));
  INVX1 g7608(.Y(n_35), .A(layer2_out[50]));
  INVX1 g7609(.Y(n_34), .A(layer2_out[83]));
  INVX1 g7610(.Y(n_33), .A(layer2_out[171]));
  INVX1 g7611(.Y(n_32), .A(layer2_out[119]));
  INVX1 g7612(.Y(n_31), .A(layer2_out[11]));
  INVX1 g7613(.Y(n_30), .A(layer2_out[166]));
  INVX1 g7614(.Y(n_29), .A(layer2_out[62]));
  INVX1 g7615(.Y(n_28), .A(layer2_out[45]));
  INVX1 g7616(.Y(n_27), .A(layer2_out[146]));
  INVX1 g7617(.Y(n_26), .A(layer2_out[4]));
  INVX1 g7618(.Y(n_25), .A(layer2_out[123]));
  INVX1 g7619(.Y(n_24), .A(layer2_out[1]));
  INVX1 g7620(.Y(n_23), .A(layer2_out[3]));
  INVX1 g7621(.Y(n_22), .A(layer2_out[56]));
  INVX1 g7622(.Y(n_21), .A(layer2_out[74]));
  INVX1 g7623(.Y(n_20), .A(layer2_out[14]));
  INVX1 g7624(.Y(n_19), .A(layer2_out[2]));
  INVX1 g7625(.Y(n_18), .A(layer2_out[25]));
  INVX1 g7626(.Y(n_17), .A(layer2_out[27]));
  INVX1 g7627(.Y(n_16), .A(layer2_out[93]));
  INVX1 g7628(.Y(n_15), .A(layer2_out[20]));
  INVX1 g7629(.Y(n_14), .A(layer2_out[139]));
  INVX1 g7630(.Y(n_13), .A(layer2_out[58]));
  INVX1 g7631(.Y(n_12), .A(layer2_out[154]));
  INVX1 g7632(.Y(n_11), .A(layer2_out[169]));
  INVX1 g7633(.Y(n_10), .A(layer2_out[59]));
  INVX1 g7634(.Y(n_9), .A(layer2_out[168]));
  INVX1 g7635(.Y(n_8), .A(layer2_out[46]));
  INVX1 g7636(.Y(n_7), .A(layer2_out[114]));
  INVX1 g7637(.Y(n_6), .A(layer2_out[118]));
  INVXL g7638(.Y(n_5), .A(layer2_out[33]));
  NAND3X1 g2(.Y(n_4), .A(n_179), .B(n_208), .C(n_234));
  SDFFRHQX1 \counter_reg[0] (.Q(counter[0]), .D(counter[0]), .SE(n_2), .SI(n_0),
     .RN(updown), .CK(clk));
  DFFRX2 done_reg(.Q(done), .QN(UNCONNECTED374), .D(n_3), .RN(updown), .CK(clk));
  DFFRHQX1 \counter_reg[1] (.Q(counter[1]), .D(n_1), .RN(updown), .CK(clk));
  NAND2BXL g22(.Y(n_3), .AN(done), .B(n_2));
  NAND2X1 g23(.Y(n_2), .A(counter[1]), .B(counter[0]));
  NAND2BX1 g24(.Y(n_1), .AN(counter[1]), .B(n_0));
  INVX1 g25(.Y(n_0), .A(counter[0]));
  DFFRHQX1 \instanceL2_out_reg_reg[0][0] (.Q(layer2_out[0]), .D(
    instanceL2_n_10857), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][1] (.Q(layer2_out[1]), .D(
    instanceL2_n_10859), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][2] (.Q(layer2_out[2]), .D(
    instanceL2_n_10860), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][3] (.Q(layer2_out[3]), .D(
    instanceL2_n_10861), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][4] (.Q(layer2_out[4]), .D(
    instanceL2_n_10862), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][5] (.Q(layer2_out[5]), .D(
    instanceL2_n_10968), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][6] (.Q(layer2_out[6]), .D(
    instanceL2_n_10864), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][7] (.Q(layer2_out[7]), .D(
    instanceL2_n_10865), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][8] (.Q(layer2_out[8]), .D(
    instanceL2_n_10866), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][9] (.Q(layer2_out[9]), .D(
    instanceL2_n_10908), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][10] (.Q(layer2_out[10]), .D(
    instanceL2_n_10868), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][11] (.Q(layer2_out[11]), .D(
    instanceL2_n_10884), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][12] (.Q(layer2_out[12]), .D(
    instanceL2_n_10869), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][13] (.Q(layer2_out[13]), .D(
    instanceL2_n_10854), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[0][14] (.Q(layer2_out[14]), .D(
    instanceL2_n_10871), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][0] (.Q(layer2_out[18]), .D(
    instanceL2_n_10872), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][1] (.Q(layer2_out[19]), .D(
    instanceL2_n_10873), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][2] (.Q(layer2_out[20]), .D(
    instanceL2_n_10982), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][3] (.Q(layer2_out[21]), .D(
    instanceL2_n_10876), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][4] (.Q(layer2_out[22]), .D(
    instanceL2_n_10984), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][5] (.Q(layer2_out[23]), .D(
    instanceL2_n_10877), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][6] (.Q(layer2_out[24]), .D(
    instanceL2_n_10969), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][7] (.Q(layer2_out[25]), .D(
    instanceL2_n_10878), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][8] (.Q(layer2_out[26]), .D(
    instanceL2_n_10879), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][9] (.Q(layer2_out[27]), .D(
    instanceL2_n_10880), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][10] (.Q(layer2_out[28]), .D(
    instanceL2_n_10976), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][11] (.Q(layer2_out[29]), .D(
    instanceL2_n_10881), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][12] (.Q(layer2_out[30]), .D(
    instanceL2_n_10882), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][13] (.Q(layer2_out[31]), .D(
    instanceL2_n_10883), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][14] (.Q(layer2_out[32]), .D(
    instanceL2_n_10953), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[1][15] (.Q(layer2_out[33]), .D(
    instanceL2_n_10886), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][0] (.Q(layer2_out[36]), .D(
    instanceL2_n_10887), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][1] (.Q(layer2_out[37]), .D(
    instanceL2_n_10889), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][2] (.Q(layer2_out[38]), .D(
    instanceL2_n_10961), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][3] (.Q(layer2_out[39]), .D(
    instanceL2_n_10891), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][4] (.Q(layer2_out[40]), .D(
    instanceL2_n_10958), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][5] (.Q(layer2_out[41]), .D(
    instanceL2_n_10892), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][6] (.Q(layer2_out[42]), .D(
    instanceL2_n_10912), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][7] (.Q(layer2_out[43]), .D(
    instanceL2_n_10895), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][8] (.Q(layer2_out[44]), .D(
    instanceL2_n_10947), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][9] (.Q(layer2_out[45]), .D(
    instanceL2_n_10896), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][10] (.Q(layer2_out[46]), .D(
    instanceL2_n_10934), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][11] (.Q(layer2_out[47]), .D(
    instanceL2_n_10897), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][12] (.Q(layer2_out[48]), .D(
    instanceL2_n_10898), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][13] (.Q(layer2_out[49]), .D(
    instanceL2_n_10899), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[2][14] (.Q(layer2_out[50]), .D(
    instanceL2_n_10885), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][0] (.Q(layer2_out[54]), .D(
    instanceL2_n_10901), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][1] (.Q(layer2_out[55]), .D(
    instanceL2_n_10906), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][2] (.Q(layer2_out[56]), .D(
    instanceL2_n_10902), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][3] (.Q(layer2_out[57]), .D(
    instanceL2_n_10900), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][4] (.Q(layer2_out[58]), .D(
    instanceL2_n_10904), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][5] (.Q(layer2_out[59]), .D(
    instanceL2_n_10893), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][6] (.Q(layer2_out[60]), .D(
    instanceL2_n_10905), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][7] (.Q(layer2_out[61]), .D(
    instanceL2_n_10855), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][8] (.Q(layer2_out[62]), .D(
    instanceL2_n_10907), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][9] (.Q(layer2_out[63]), .D(
    instanceL2_n_10823), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][10] (.Q(layer2_out[64]), .D(
    instanceL2_n_10986), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][11] (.Q(layer2_out[65]), .D(
    instanceL2_n_10870), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][12] (.Q(layer2_out[66]), .D(
    instanceL2_n_10910), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][13] (.Q(layer2_out[67]), .D(
    instanceL2_n_10863), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[3][14] (.Q(layer2_out[68]), .D(
    instanceL2_n_10911), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][0] (.Q(layer2_out[72]), .D(
    instanceL2_n_10843), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][1] (.Q(layer2_out[73]), .D(
    instanceL2_n_10913), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][2] (.Q(layer2_out[74]), .D(
    instanceL2_n_10914), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][3] (.Q(layer2_out[75]), .D(
    instanceL2_n_10915), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][4] (.Q(layer2_out[76]), .D(
    instanceL2_n_10851), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][5] (.Q(layer2_out[77]), .D(
    instanceL2_n_10916), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][6] (.Q(layer2_out[78]), .D(
    instanceL2_n_10917), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][7] (.Q(layer2_out[79]), .D(
    instanceL2_n_10918), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][8] (.Q(layer2_out[80]), .D(
    instanceL2_n_10844), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][9] (.Q(layer2_out[81]), .D(
    instanceL2_n_10921), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][10] (.Q(layer2_out[82]), .D(
    instanceL2_n_10922), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][11] (.Q(layer2_out[83]), .D(
    instanceL2_n_10926), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][12] (.Q(layer2_out[84]), .D(
    instanceL2_n_10850), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][13] (.Q(layer2_out[85]), .D(
    instanceL2_n_10931), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[4][14] (.Q(layer2_out[86]), .D(
    instanceL2_n_10849), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][0] (.Q(layer2_out[90]), .D(
    instanceL2_n_10933), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][1] (.Q(layer2_out[91]), .D(
    instanceL2_n_10847), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][2] (.Q(layer2_out[92]), .D(
    instanceL2_n_10935), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][3] (.Q(layer2_out[93]), .D(
    instanceL2_n_10848), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][4] (.Q(layer2_out[94]), .D(
    instanceL2_n_10938), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][5] (.Q(layer2_out[95]), .D(
    instanceL2_n_10836), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][6] (.Q(layer2_out[96]), .D(
    instanceL2_n_10941), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][7] (.Q(layer2_out[97]), .D(
    instanceL2_n_10841), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][8] (.Q(layer2_out[98]), .D(
    instanceL2_n_10946), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][9] (.Q(layer2_out[99]), .D(
    instanceL2_n_10842), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][10] (.Q(layer2_out[100]), .D(
    instanceL2_n_10948), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][11] (.Q(layer2_out[101]), .D(
    instanceL2_n_10949), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][12] (.Q(layer2_out[102]), .D(
    instanceL2_n_10950), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][13] (.Q(layer2_out[103]), .D(
    instanceL2_n_10824), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[5][14] (.Q(layer2_out[104]), .D(
    instanceL2_n_10951), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][0] (.Q(layer2_out[108]), .D(
    instanceL2_n_10975), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][1] (.Q(layer2_out[109]), .D(
    instanceL2_n_10952), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][2] (.Q(layer2_out[110]), .D(
    instanceL2_n_10985), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][3] (.Q(layer2_out[111]), .D(
    instanceL2_n_10954), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][4] (.Q(layer2_out[112]), .D(
    instanceL2_n_10955), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][5] (.Q(layer2_out[113]), .D(
    instanceL2_n_10956), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][6] (.Q(layer2_out[114]), .D(
    instanceL2_n_10909), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][7] (.Q(layer2_out[115]), .D(
    instanceL2_n_10945), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][8] (.Q(layer2_out[116]), .D(
    instanceL2_n_10983), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][9] (.Q(layer2_out[117]), .D(
    instanceL2_n_10944), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][10] (.Q(layer2_out[118]), .D(
    instanceL2_n_10979), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][11] (.Q(layer2_out[119]), .D(
    instanceL2_n_10943), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][12] (.Q(layer2_out[120]), .D(
    instanceL2_n_10929), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][13] (.Q(layer2_out[121]), .D(
    instanceL2_n_10942), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][14] (.Q(layer2_out[122]), .D(
    instanceL2_n_10964), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[6][15] (.Q(layer2_out[123]), .D(
    instanceL2_n_10960), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][0] (.Q(layer2_out[126]), .D(
    instanceL2_n_10957), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][1] (.Q(layer2_out[127]), .D(
    instanceL2_n_10940), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][2] (.Q(layer2_out[128]), .D(
    instanceL2_n_10939), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][3] (.Q(layer2_out[129]), .D(
    instanceL2_n_10962), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][4] (.Q(layer2_out[130]), .D(
    instanceL2_n_10867), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][5] (.Q(layer2_out[131]), .D(
    instanceL2_n_10963), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][6] (.Q(layer2_out[132]), .D(
    instanceL2_n_10903), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][7] (.Q(layer2_out[133]), .D(
    instanceL2_n_10937), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][8] (.Q(layer2_out[134]), .D(
    instanceL2_n_10890), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][9] (.Q(layer2_out[135]), .D(
    instanceL2_n_10936), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][10] (.Q(layer2_out[136]), .D(
    instanceL2_n_10875), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][11] (.Q(layer2_out[137]), .D(
    instanceL2_n_10965), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][12] (.Q(layer2_out[138]), .D(
    instanceL2_n_10834), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][13] (.Q(layer2_out[139]), .D(
    instanceL2_n_10966), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][14] (.Q(layer2_out[140]), .D(
    instanceL2_n_10852), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[7][15] (.Q(layer2_out[141]), .D(
    instanceL2_n_10967), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][0] (.Q(layer2_out[144]), .D(
    instanceL2_n_10846), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][1] (.Q(layer2_out[145]), .D(
    instanceL2_n_10932), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][2] (.Q(layer2_out[146]), .D(
    instanceL2_n_10839), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][3] (.Q(layer2_out[147]), .D(
    instanceL2_n_10970), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][4] (.Q(layer2_out[148]), .D(
    instanceL2_n_10838), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][5] (.Q(layer2_out[149]), .D(
    instanceL2_n_10971), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][6] (.Q(layer2_out[150]), .D(
    instanceL2_n_10840), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][7] (.Q(layer2_out[151]), .D(
    instanceL2_n_10928), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][8] (.Q(layer2_out[152]), .D(
    instanceL2_n_10829), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][9] (.Q(layer2_out[153]), .D(
    instanceL2_n_10927), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][10] (.Q(layer2_out[154]), .D(
    instanceL2_n_10835), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][11] (.Q(layer2_out[155]), .D(
    instanceL2_n_10974), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][12] (.Q(layer2_out[156]), .D(
    instanceL2_n_10832), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[8][13] (.Q(layer2_out[157]), .D(
    instanceL2_n_10925), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][0] (.Q(layer2_out[162]), .D(
    instanceL2_n_10825), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][1] (.Q(layer2_out[163]), .D(
    instanceL2_n_10924), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][2] (.Q(layer2_out[164]), .D(
    instanceL2_n_10972), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][3] (.Q(layer2_out[165]), .D(
    instanceL2_n_10923), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][4] (.Q(layer2_out[166]), .D(
    instanceL2_n_10973), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][5] (.Q(layer2_out[167]), .D(
    instanceL2_n_10977), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][6] (.Q(layer2_out[168]), .D(
    instanceL2_n_10959), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][7] (.Q(layer2_out[169]), .D(
    instanceL2_n_10978), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][8] (.Q(layer2_out[170]), .D(
    instanceL2_n_10830), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][9] (.Q(layer2_out[171]), .D(
    instanceL2_n_10920), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][10] (.Q(layer2_out[172]), .D(
    instanceL2_n_10894), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][11] (.Q(layer2_out[173]), .D(
    instanceL2_n_10919), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][12] (.Q(layer2_out[174]), .D(
    instanceL2_n_10831), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][13] (.Q(layer2_out[175]), .D(
    instanceL2_n_10980), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][14] (.Q(layer2_out[176]), .D(
    instanceL2_n_10826), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][15] (.Q(layer2_out[177]), .D(
    instanceL2_n_10981), .RN(rst_n), .CK(clk));
  DFFRHQX1 \instanceL2_out_reg_reg[9][16] (.Q(layer2_out[178]), .D(
    instanceL2_n_10828), .RN(rst_n), .CK(clk));
  NOR2BX1 instanceL2_g10110(.Y(instanceL2_n_10823), .AN(
    \instanceL2_row_sums[3] [9]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10111(.Y(instanceL2_n_10824), .AN(
    \instanceL2_row_sums[5] [13]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10112(.Y(instanceL2_n_10825), .AN(
    \instanceL2_row_sums[9] [0]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10113(.Y(instanceL2_n_10826), .AN(
    \instanceL2_row_sums[9] [14]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10114(.Y(instanceL2_n_10828), .AN(
    \instanceL2_row_sums[9] [16]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10115(.Y(instanceL2_n_10829), .AN(
    \instanceL2_row_sums[8] [8]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10116(.Y(instanceL2_n_10830), .AN(
    \instanceL2_row_sums[9] [8]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10117(.Y(instanceL2_n_10831), .AN(
    \instanceL2_row_sums[9] [12]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10118(.Y(instanceL2_n_10832), .AN(
    \instanceL2_row_sums[8] [12]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10119(.Y(instanceL2_n_10834), .AN(
    \instanceL2_row_sums[7] [12]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10120(.Y(instanceL2_n_10835), .AN(
    \instanceL2_row_sums[8] [10]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10121(.Y(instanceL2_n_10836), .AN(
    \instanceL2_row_sums[5] [5]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10122(.Y(instanceL2_n_10838), .AN(
    \instanceL2_row_sums[8] [4]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10123(.Y(instanceL2_n_10839), .AN(
    \instanceL2_row_sums[8] [2]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10124(.Y(instanceL2_n_10840), .AN(
    \instanceL2_row_sums[8] [6]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10125(.Y(instanceL2_n_10841), .AN(
    \instanceL2_row_sums[5] [7]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10126(.Y(instanceL2_n_10842), .AN(
    \instanceL2_row_sums[5] [9]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10127(.Y(instanceL2_n_10843), .AN(
    \instanceL2_row_sums[4] [0]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10128(.Y(instanceL2_n_10844), .AN(
    \instanceL2_row_sums[4] [8]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10129(.Y(instanceL2_n_10846), .AN(
    \instanceL2_row_sums[8] [0]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10130(.Y(instanceL2_n_10847), .AN(
    \instanceL2_row_sums[5] [1]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10131(.Y(instanceL2_n_10848), .AN(
    \instanceL2_row_sums[5] [3]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10132(.Y(instanceL2_n_10849), .AN(
    \instanceL2_row_sums[4] [14]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10133(.Y(instanceL2_n_10850), .AN(
    \instanceL2_row_sums[4] [12]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10134(.Y(instanceL2_n_10851), .AN(
    \instanceL2_row_sums[4] [4]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10135(.Y(instanceL2_n_10852), .AN(
    \instanceL2_row_sums[7] [14]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10136(.Y(instanceL2_n_10854), .AN(
    \instanceL2_row_sums[0] [13]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10137(.Y(instanceL2_n_10855), .AN(
    \instanceL2_row_sums[3] [7]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10138(.Y(instanceL2_n_10857), .AN(
    \instanceL2_row_sums[0] [0]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10139(.Y(instanceL2_n_10859), .AN(
    \instanceL2_row_sums[0] [1]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10140(.Y(instanceL2_n_10860), .AN(
    \instanceL2_row_sums[0] [2]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10141(.Y(instanceL2_n_10861), .AN(
    \instanceL2_row_sums[0] [3]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10142(.Y(instanceL2_n_10862), .AN(
    \instanceL2_row_sums[0] [4]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10143(.Y(instanceL2_n_10863), .AN(
    \instanceL2_row_sums[3] [13]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10144(.Y(instanceL2_n_10864), .AN(
    \instanceL2_row_sums[0] [6]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10145(.Y(instanceL2_n_10865), .AN(
    \instanceL2_row_sums[0] [7]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10146(.Y(instanceL2_n_10866), .AN(
    \instanceL2_row_sums[0] [8]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10147(.Y(instanceL2_n_10867), .AN(
    \instanceL2_row_sums[7] [4]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10148(.Y(instanceL2_n_10868), .AN(
    \instanceL2_row_sums[0] [10]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10149(.Y(instanceL2_n_10869), .AN(
    \instanceL2_row_sums[0] [12]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10150(.Y(instanceL2_n_10870), .AN(
    \instanceL2_row_sums[3] [11]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10151(.Y(instanceL2_n_10871), .AN(
    \instanceL2_row_sums[0] [14]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10152(.Y(instanceL2_n_10872), .AN(
    \instanceL2_row_sums[1] [0]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10153(.Y(instanceL2_n_10873), .AN(
    \instanceL2_row_sums[1] [1]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10154(.Y(instanceL2_n_10875), .AN(
    \instanceL2_row_sums[7] [10]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10155(.Y(instanceL2_n_10876), .AN(
    \instanceL2_row_sums[1] [3]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10156(.Y(instanceL2_n_10877), .AN(
    \instanceL2_row_sums[1] [5]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10157(.Y(instanceL2_n_10878), .AN(
    \instanceL2_row_sums[1] [7]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10158(.Y(instanceL2_n_10879), .AN(
    \instanceL2_row_sums[1] [8]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10159(.Y(instanceL2_n_10880), .AN(
    \instanceL2_row_sums[1] [9]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10160(.Y(instanceL2_n_10881), .AN(
    \instanceL2_row_sums[1] [11]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10161(.Y(instanceL2_n_10882), .AN(
    \instanceL2_row_sums[1] [12]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10162(.Y(instanceL2_n_10883), .AN(
    \instanceL2_row_sums[1] [13]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10163(.Y(instanceL2_n_10884), .AN(
    \instanceL2_row_sums[0] [11]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10164(.Y(instanceL2_n_10885), .AN(
    \instanceL2_row_sums[2] [14]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10165(.Y(instanceL2_n_10886), .AN(
    \instanceL2_row_sums[1] [15]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10166(.Y(instanceL2_n_10887), .AN(
    \instanceL2_row_sums[2] [0]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10167(.Y(instanceL2_n_10889), .AN(
    \instanceL2_row_sums[2] [1]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10168(.Y(instanceL2_n_10890), .AN(
    \instanceL2_row_sums[7] [8]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10169(.Y(instanceL2_n_10891), .AN(
    \instanceL2_row_sums[2] [3]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10170(.Y(instanceL2_n_10892), .AN(
    \instanceL2_row_sums[2] [5]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10171(.Y(instanceL2_n_10893), .AN(
    \instanceL2_row_sums[3] [5]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10172(.Y(instanceL2_n_10894), .AN(
    \instanceL2_row_sums[9] [10]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10173(.Y(instanceL2_n_10895), .AN(
    \instanceL2_row_sums[2] [7]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10174(.Y(instanceL2_n_10896), .AN(
    \instanceL2_row_sums[2] [9]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10175(.Y(instanceL2_n_10897), .AN(
    \instanceL2_row_sums[2] [11]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10176(.Y(instanceL2_n_10898), .AN(
    \instanceL2_row_sums[2] [12]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10177(.Y(instanceL2_n_10899), .AN(
    \instanceL2_row_sums[2] [13]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10178(.Y(instanceL2_n_10900), .AN(
    \instanceL2_row_sums[3] [3]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10179(.Y(instanceL2_n_10901), .AN(
    \instanceL2_row_sums[3] [0]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10180(.Y(instanceL2_n_10902), .AN(
    \instanceL2_row_sums[3] [2]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10181(.Y(instanceL2_n_10903), .AN(
    \instanceL2_row_sums[7] [6]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10182(.Y(instanceL2_n_10904), .AN(
    \instanceL2_row_sums[3] [4]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10183(.Y(instanceL2_n_10905), .AN(
    \instanceL2_row_sums[3] [6]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10184(.Y(instanceL2_n_10906), .AN(
    \instanceL2_row_sums[3] [1]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10185(.Y(instanceL2_n_10907), .AN(
    \instanceL2_row_sums[3] [8]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10186(.Y(instanceL2_n_10908), .AN(
    \instanceL2_row_sums[0] [9]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10187(.Y(instanceL2_n_10909), .AN(
    \instanceL2_row_sums[6] [6]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10188(.Y(instanceL2_n_10910), .AN(
    \instanceL2_row_sums[3] [12]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10189(.Y(instanceL2_n_10911), .AN(
    \instanceL2_row_sums[3] [14]), .B(\instanceL2_row_sums[3] [18]));
  NOR2BX1 instanceL2_g10190(.Y(instanceL2_n_10912), .AN(
    \instanceL2_row_sums[2] [6]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10191(.Y(instanceL2_n_10913), .AN(
    \instanceL2_row_sums[4] [1]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10192(.Y(instanceL2_n_10914), .AN(
    \instanceL2_row_sums[4] [2]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10193(.Y(instanceL2_n_10915), .AN(
    \instanceL2_row_sums[4] [3]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10194(.Y(instanceL2_n_10916), .AN(
    \instanceL2_row_sums[4] [5]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10195(.Y(instanceL2_n_10917), .AN(
    \instanceL2_row_sums[4] [6]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10196(.Y(instanceL2_n_10918), .AN(
    \instanceL2_row_sums[4] [7]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10197(.Y(instanceL2_n_10919), .AN(
    \instanceL2_row_sums[9] [11]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10198(.Y(instanceL2_n_10920), .AN(
    \instanceL2_row_sums[9] [9]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10199(.Y(instanceL2_n_10921), .AN(
    \instanceL2_row_sums[4] [9]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10200(.Y(instanceL2_n_10922), .AN(
    \instanceL2_row_sums[4] [10]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10201(.Y(instanceL2_n_10923), .AN(
    \instanceL2_row_sums[9] [3]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10202(.Y(instanceL2_n_10924), .AN(
    \instanceL2_row_sums[9] [1]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10203(.Y(instanceL2_n_10925), .AN(
    \instanceL2_row_sums[8] [13]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10204(.Y(instanceL2_n_10926), .AN(
    \instanceL2_row_sums[4] [11]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10205(.Y(instanceL2_n_10927), .AN(
    \instanceL2_row_sums[8] [9]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10206(.Y(instanceL2_n_10928), .AN(
    \instanceL2_row_sums[8] [7]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10207(.Y(instanceL2_n_10929), .AN(
    \instanceL2_row_sums[6] [12]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10208(.Y(instanceL2_n_10931), .AN(
    \instanceL2_row_sums[4] [13]), .B(\instanceL2_row_sums[4] [18]));
  NOR2BX1 instanceL2_g10209(.Y(instanceL2_n_10932), .AN(
    \instanceL2_row_sums[8] [1]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10210(.Y(instanceL2_n_10933), .AN(
    \instanceL2_row_sums[5] [0]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10211(.Y(instanceL2_n_10934), .AN(
    \instanceL2_row_sums[2] [10]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10212(.Y(instanceL2_n_10935), .AN(
    \instanceL2_row_sums[5] [2]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10213(.Y(instanceL2_n_10936), .AN(
    \instanceL2_row_sums[7] [9]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10214(.Y(instanceL2_n_10937), .AN(
    \instanceL2_row_sums[7] [7]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10215(.Y(instanceL2_n_10938), .AN(
    \instanceL2_row_sums[5] [4]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10216(.Y(instanceL2_n_10939), .AN(
    \instanceL2_row_sums[7] [2]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10217(.Y(instanceL2_n_10940), .AN(
    \instanceL2_row_sums[7] [1]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10218(.Y(instanceL2_n_10941), .AN(
    \instanceL2_row_sums[5] [6]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10219(.Y(instanceL2_n_10942), .AN(
    \instanceL2_row_sums[6] [13]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10220(.Y(instanceL2_n_10943), .AN(
    \instanceL2_row_sums[6] [11]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10221(.Y(instanceL2_n_10944), .AN(
    \instanceL2_row_sums[6] [9]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10222(.Y(instanceL2_n_10945), .AN(
    \instanceL2_row_sums[6] [7]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10223(.Y(instanceL2_n_10946), .AN(
    \instanceL2_row_sums[5] [8]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10224(.Y(instanceL2_n_10947), .AN(
    \instanceL2_row_sums[2] [8]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10225(.Y(instanceL2_n_10948), .AN(
    \instanceL2_row_sums[5] [10]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10226(.Y(instanceL2_n_10949), .AN(
    \instanceL2_row_sums[5] [11]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10227(.Y(instanceL2_n_10950), .AN(
    \instanceL2_row_sums[5] [12]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10228(.Y(instanceL2_n_10951), .AN(
    \instanceL2_row_sums[5] [14]), .B(\instanceL2_row_sums[5] [18]));
  NOR2BX1 instanceL2_g10229(.Y(instanceL2_n_10952), .AN(
    \instanceL2_row_sums[6] [1]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10230(.Y(instanceL2_n_10953), .AN(
    \instanceL2_row_sums[1] [14]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10231(.Y(instanceL2_n_10954), .AN(
    \instanceL2_row_sums[6] [3]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10232(.Y(instanceL2_n_10955), .AN(
    \instanceL2_row_sums[6] [4]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10233(.Y(instanceL2_n_10956), .AN(
    \instanceL2_row_sums[6] [5]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10234(.Y(instanceL2_n_10957), .AN(
    \instanceL2_row_sums[7] [0]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10235(.Y(instanceL2_n_10958), .AN(
    \instanceL2_row_sums[2] [4]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10236(.Y(instanceL2_n_10959), .AN(
    \instanceL2_row_sums[9] [6]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10237(.Y(instanceL2_n_10960), .AN(
    \instanceL2_row_sums[6] [15]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10238(.Y(instanceL2_n_10961), .AN(
    \instanceL2_row_sums[2] [2]), .B(\instanceL2_row_sums[2] [18]));
  NOR2BX1 instanceL2_g10239(.Y(instanceL2_n_10962), .AN(
    \instanceL2_row_sums[7] [3]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10240(.Y(instanceL2_n_10963), .AN(
    \instanceL2_row_sums[7] [5]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10241(.Y(instanceL2_n_10964), .AN(
    \instanceL2_row_sums[6] [14]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10242(.Y(instanceL2_n_10965), .AN(
    \instanceL2_row_sums[7] [11]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10243(.Y(instanceL2_n_10966), .AN(
    \instanceL2_row_sums[7] [13]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10244(.Y(instanceL2_n_10967), .AN(
    \instanceL2_row_sums[7] [15]), .B(\instanceL2_row_sums[7] [18]));
  NOR2BX1 instanceL2_g10245(.Y(instanceL2_n_10968), .AN(
    \instanceL2_row_sums[0] [5]), .B(\instanceL2_row_sums[0] [18]));
  NOR2BX1 instanceL2_g10246(.Y(instanceL2_n_10969), .AN(
    \instanceL2_row_sums[1] [6]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10247(.Y(instanceL2_n_10970), .AN(
    \instanceL2_row_sums[8] [3]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10248(.Y(instanceL2_n_10971), .AN(
    \instanceL2_row_sums[8] [5]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10249(.Y(instanceL2_n_10972), .AN(
    \instanceL2_row_sums[9] [2]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10250(.Y(instanceL2_n_10973), .AN(
    \instanceL2_row_sums[9] [4]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10251(.Y(instanceL2_n_10974), .AN(
    \instanceL2_row_sums[8] [11]), .B(\instanceL2_row_sums[8] [18]));
  NOR2BX1 instanceL2_g10252(.Y(instanceL2_n_10975), .AN(
    \instanceL2_row_sums[6] [0]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10253(.Y(instanceL2_n_10976), .AN(
    \instanceL2_row_sums[1] [10]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10254(.Y(instanceL2_n_10977), .AN(
    \instanceL2_row_sums[9] [5]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10255(.Y(instanceL2_n_10978), .AN(
    \instanceL2_row_sums[9] [7]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10256(.Y(instanceL2_n_10979), .AN(
    \instanceL2_row_sums[6] [10]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10257(.Y(instanceL2_n_10980), .AN(
    \instanceL2_row_sums[9] [13]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10258(.Y(instanceL2_n_10981), .AN(
    \instanceL2_row_sums[9] [15]), .B(\instanceL2_row_sums[9] [18]));
  NOR2BX1 instanceL2_g10259(.Y(instanceL2_n_10982), .AN(
    \instanceL2_row_sums[1] [2]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10260(.Y(instanceL2_n_10983), .AN(
    \instanceL2_row_sums[6] [8]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10261(.Y(instanceL2_n_10984), .AN(
    \instanceL2_row_sums[1] [4]), .B(\instanceL2_row_sums[1] [18]));
  NOR2BX1 instanceL2_g10262(.Y(instanceL2_n_10985), .AN(
    \instanceL2_row_sums[6] [2]), .B(\instanceL2_row_sums[6] [18]));
  NOR2BX1 instanceL2_g10263(.Y(instanceL2_n_10986), .AN(
    \instanceL2_row_sums[3] [10]), .B(\instanceL2_row_sums[3] [18]));
  OAI2BB1X1 instanceL2_g10488(.Y(\instanceL2_prod_terms[0][4][10] ), .A0N(
    instanceL2_n_11250), .A1N(instanceL2_n_11176), .B0(instanceL2_n_11171));
  OAI2BB1X1 instanceL2_g10489(.Y(\instanceL2_prod_terms[7][4] [10]), .A0N(
    instanceL2_n_11250), .A1N(instanceL2_n_11173), .B0(instanceL2_n_11171));
  OR2X1 instanceL2_g10490(.Y(instanceL2_n_11171), .A(instanceL2_n_11250), .B(
    instanceL2_n_11173));
  ADDFX1 instanceL2_g10491(.CO(instanceL2_n_11173), .S(
    \instanceL2_prod_terms[7][4] [9]), .A(instanceL2_n_11334), .B(
    instanceL2_n_11303), .CI(instanceL2_n_11181));
  ADDFX1 instanceL2_g10492(.CO(instanceL2_n_11176), .S(
    \instanceL2_prod_terms[0][4][9] ), .A(instanceL2_n_11303), .B(
    instanceL2_n_11283), .CI(instanceL2_n_11179));
  ADDFX1 instanceL2_g10493(.CO(instanceL2_n_11179), .S(
    \instanceL2_prod_terms[0][4][8] ), .A(instanceL2_n_11275), .B(
    instanceL2_n_11261), .CI(instanceL2_n_11192));
  ADDFX1 instanceL2_g10494(.CO(instanceL2_n_11181), .S(
    \instanceL2_prod_terms[7][4] [8]), .A(instanceL2_n_11311), .B(
    instanceL2_n_11271), .CI(instanceL2_n_11190));
  AOI21X1 instanceL2_g10495(.Y(\instanceL2_prod_terms[1][4] [9]), .A0(
    instanceL2_n_11347), .A1(instanceL2_n_11199), .B0(
    \instanceL2_prod_terms[1][4] [10]));
  NOR2X1 instanceL2_g10496(.Y(\instanceL2_prod_terms[1][4] [10]), .A(
    instanceL2_n_11347), .B(instanceL2_n_11199));
  AOI21X1 instanceL2_g10497(.Y(\instanceL2_prod_terms[5][4] [9]), .A0(
    layer1_out[43]), .A1(instanceL2_n_11203), .B0(instanceL2_n_11194));
  ADDFX1 instanceL2_g10498(.CO(instanceL2_n_11190), .S(
    \instanceL2_prod_terms[7][4] [7]), .A(instanceL2_n_11274), .B(
    instanceL2_n_11253), .CI(instanceL2_n_11207));
  ADDFX1 instanceL2_g10499(.CO(instanceL2_n_11192), .S(
    \instanceL2_prod_terms[0][4][7] ), .A(instanceL2_n_11279), .B(
    instanceL2_n_11258), .CI(instanceL2_n_11205));
  INVX1 instanceL2_g10500(.Y(\instanceL2_prod_terms[5][4] [13]), .A(
    instanceL2_n_11194));
  NOR2X1 instanceL2_g10501(.Y(instanceL2_n_11194), .A(layer1_out[43]), .B(
    instanceL2_n_11203));
  OA21X1 instanceL2_g10502(.Y(\instanceL2_prod_terms[1][4] [8]), .A0(
    layer1_out[42]), .A1(instanceL2_n_11210), .B0(instanceL2_n_11199));
  NAND2X1 instanceL2_g10503(.Y(instanceL2_n_11199), .A(layer1_out[42]), .B(
    instanceL2_n_11210));
  OA21X1 instanceL2_g10504(.Y(\instanceL2_prod_terms[5][4] [8]), .A0(
    instanceL2_n_11337), .A1(instanceL2_n_11222), .B0(instanceL2_n_11203));
  ADDFX1 instanceL2_g10505(.CO(instanceL2_n_11205), .S(
    \instanceL2_prod_terms[0][4][6] ), .A(instanceL2_n_11286), .B(
    instanceL2_n_11254), .CI(instanceL2_n_11218));
  ADDFX1 instanceL2_g10506(.CO(instanceL2_n_11207), .S(
    \instanceL2_prod_terms[7][4] [6]), .A(instanceL2_n_11272), .B(
    instanceL2_n_11256), .CI(instanceL2_n_11220));
  NAND2X1 instanceL2_g10507(.Y(instanceL2_n_11203), .A(instanceL2_n_11337), .B(
    instanceL2_n_11222));
  XNOR2X1 instanceL2_g10508(.Y(\instanceL2_prod_terms[1][4] [7]), .A(
    instanceL2_n_11294), .B(instanceL2_n_11215));
  OAI21X1 instanceL2_g10509(.Y(instanceL2_n_11210), .A0(instanceL2_n_11320), .A1(
    instanceL2_n_11214), .B0(instanceL2_n_11321));
  AOI21X1 instanceL2_g10510(.Y(\instanceL2_prod_terms[5][4] [7]), .A0(
    layer1_out[41]), .A1(instanceL2_n_11231), .B0(instanceL2_n_11222));
  INVX1 instanceL2_g10511(.Y(instanceL2_n_11214), .A(instanceL2_n_11215));
  XNOR2X1 instanceL2_g10512(.Y(\instanceL2_prod_terms[1][4] [6]), .A(
    instanceL2_n_11295), .B(instanceL2_n_11227));
  OAI21X1 instanceL2_g10513(.Y(instanceL2_n_11215), .A0(instanceL2_n_11329), .A1(
    instanceL2_n_11226), .B0(instanceL2_n_11319));
  ADDFX1 instanceL2_g10514(.CO(instanceL2_n_11218), .S(
    \instanceL2_prod_terms[0][4][5] ), .A(instanceL2_n_11333), .B(
    instanceL2_n_11252), .CI(instanceL2_n_11236));
  ADDFX1 instanceL2_g10515(.CO(instanceL2_n_11220), .S(
    \instanceL2_prod_terms[7][4] [5]), .A(instanceL2_n_11333), .B(
    instanceL2_n_11263), .CI(instanceL2_n_11233));
  NOR2X1 instanceL2_g10516(.Y(instanceL2_n_11222), .A(layer1_out[41]), .B(
    instanceL2_n_11231));
  INVX1 instanceL2_g10517(.Y(instanceL2_n_11226), .A(instanceL2_n_11227));
  OAI2BB1X1 instanceL2_g10518(.Y(instanceL2_n_11227), .A0N(instanceL2_n_11330),
     .A1N(instanceL2_n_11239), .B0(instanceL2_n_11331));
  XNOR2X1 instanceL2_g10519(.Y(\instanceL2_prod_terms[1][4] [5]), .A(
    instanceL2_n_11310), .B(instanceL2_n_11239));
  OA21X1 instanceL2_g10520(.Y(\instanceL2_prod_terms[5][4] [6]), .A0(
    instanceL2_n_11351), .A1(instanceL2_n_11248), .B0(instanceL2_n_11231));
  ADDFX1 instanceL2_g10521(.CO(instanceL2_n_11233), .S(
    \instanceL2_prod_terms[7][4] [4]), .A(layer1_out[40]), .B(
    instanceL2_n_11322), .CI(\instanceL2_prod_terms[5][4] [3]));
  ADDFX1 instanceL2_g10522(.CO(instanceL2_n_11236), .S(
    \instanceL2_prod_terms[0][4][4] ), .A(layer1_out[39]), .B(
    instanceL2_n_11266), .CI(\instanceL2_prod_terms[5][4] [3]));
  NAND2X1 instanceL2_g10523(.Y(instanceL2_n_11231), .A(instanceL2_n_11351), .B(
    instanceL2_n_11248));
  XNOR2X1 instanceL2_g10524(.Y(\instanceL2_prod_terms[1][4] [4]), .A(
    instanceL2_n_11293), .B(instanceL2_n_11244));
  OAI21X1 instanceL2_g10525(.Y(instanceL2_n_11239), .A0(instanceL2_n_11328), .A1(
    instanceL2_n_11244), .B0(instanceL2_n_11327));
  INVX1 instanceL2_g10526(.Y(\instanceL2_prod_terms[1][4] [3]), .A(
    instanceL2_n_11245));
  ADDFX1 instanceL2_g10527(.CO(instanceL2_n_11244), .S(instanceL2_n_11245), .A(
    instanceL2_n_11343), .B(instanceL2_n_11349), .CI(instanceL2_n_11323));
  AOI21X1 instanceL2_g10528(.Y(\instanceL2_prod_terms[5][4] [5]), .A0(
    layer1_out[39]), .A1(instanceL2_n_11289), .B0(instanceL2_n_11248));
  NOR2X1 instanceL2_g10529(.Y(instanceL2_n_11248), .A(layer1_out[39]), .B(
    instanceL2_n_11289));
  XNOR2X1 instanceL2_g10530(.Y(instanceL2_n_11250), .A(instanceL2_n_11332), .B(
    instanceL2_n_11309));
  XNOR2X1 instanceL2_g10531(.Y(instanceL2_n_11252), .A(layer1_out[38]), .B(
    instanceL2_n_11308));
  XNOR2X1 instanceL2_g10532(.Y(instanceL2_n_11253), .A(layer1_out[39]), .B(
    instanceL2_n_11292));
  MXI2XL instanceL2_g10533(.Y(instanceL2_n_11254), .A(layer1_out[39]), .B(
    instanceL2_n_11343), .S0(instanceL2_n_11291));
  XNOR2X1 instanceL2_g10534(.Y(instanceL2_n_11256), .A(layer1_out[38]), .B(
    instanceL2_n_11290));
  MXI2XL instanceL2_g10535(.Y(instanceL2_n_11258), .A(layer1_out[40]), .B(
    instanceL2_n_11351), .S0(instanceL2_n_11290));
  XNOR2X1 instanceL2_g10536(.Y(instanceL2_n_11261), .A(layer1_out[41]), .B(
    instanceL2_n_11292));
  MXI2XL instanceL2_g10537(.Y(instanceL2_n_11263), .A(layer1_out[37]), .B(
    instanceL2_n_11349), .S0(instanceL2_n_11291));
  INVX1 instanceL2_g10538(.Y(instanceL2_n_11266), .A(instanceL2_n_11323));
  OAI21X1 instanceL2_g10539(.Y(instanceL2_n_11271), .A0(layer1_out[39]), .A1(
    instanceL2_n_11314), .B0(instanceL2_n_11317));
  OAI21X1 instanceL2_g10540(.Y(instanceL2_n_11272), .A0(layer1_out[37]), .A1(
    instanceL2_n_11318), .B0(instanceL2_n_11315));
  OAI21X1 instanceL2_g10541(.Y(instanceL2_n_11274), .A0(layer1_out[38]), .A1(
    instanceL2_n_11325), .B0(instanceL2_n_11326));
  OAI21X1 instanceL2_g10542(.Y(instanceL2_n_11275), .A0(layer1_out[39]), .A1(
    instanceL2_n_11329), .B0(instanceL2_n_11319));
  OA21X1 instanceL2_g10543(.Y(\instanceL2_prod_terms[5][4] [4]), .A0(
    instanceL2_n_11339), .A1(instanceL2_n_11316), .B0(instanceL2_n_11289));
  OAI2BB1X1 instanceL2_g10544(.Y(instanceL2_n_11279), .A0N(instanceL2_n_11339),
     .A1N(instanceL2_n_11330), .B0(instanceL2_n_11331));
  OAI21X1 instanceL2_g10545(.Y(instanceL2_n_11283), .A0(layer1_out[40]), .A1(
    instanceL2_n_11320), .B0(instanceL2_n_11321));
  OAI21X1 instanceL2_g10546(.Y(instanceL2_n_11286), .A0(layer1_out[37]), .A1(
    instanceL2_n_11328), .B0(instanceL2_n_11327));
  NOR2BX1 instanceL2_g10547(.Y(instanceL2_n_11293), .AN(instanceL2_n_11327), .B(
    instanceL2_n_11328));
  NAND2BX1 instanceL2_g10548(.Y(instanceL2_n_11294), .AN(instanceL2_n_11320), .B(
    instanceL2_n_11321));
  NAND2BX1 instanceL2_g10549(.Y(instanceL2_n_11295), .AN(instanceL2_n_11329), .B(
    instanceL2_n_11319));
  NAND2X1 instanceL2_g10550(.Y(instanceL2_n_11289), .A(instanceL2_n_11339), .B(
    instanceL2_n_11316));
  NOR2BX1 instanceL2_g10551(.Y(instanceL2_n_11290), .AN(instanceL2_n_11326), .B(
    instanceL2_n_11325));
  NOR2BX1 instanceL2_g10552(.Y(instanceL2_n_11291), .AN(instanceL2_n_11315), .B(
    instanceL2_n_11318));
  NOR2BX1 instanceL2_g10553(.Y(instanceL2_n_11292), .AN(instanceL2_n_11317), .B(
    instanceL2_n_11314));
  AOI21X1 instanceL2_g10554(.Y(\instanceL2_prod_terms[7][4] [3]), .A0(
    instanceL2_n_11343), .A1(instanceL2_n_11345), .B0(instanceL2_n_11322));
  OA21X1 instanceL2_g10555(.Y(\instanceL2_prod_terms[1][4] [2]), .A0(
    layer1_out[36]), .A1(layer1_out[38]), .B0(instanceL2_n_11323));
  AOI22X1 instanceL2_g10556(.Y(instanceL2_n_11308), .A0(instanceL2_n_11351), .A1(
    instanceL2_n_11349), .B0(layer1_out[40]), .B1(layer1_out[37]));
  OAI22X1 instanceL2_g10557(.Y(instanceL2_n_11309), .A0(layer1_out[43]), .A1(
    layer1_out[42]), .B0(instanceL2_n_11347), .B1(instanceL2_n_11337));
  NAND2XL instanceL2_g10558(.Y(instanceL2_n_11310), .A(instanceL2_n_11331), .B(
    instanceL2_n_11330));
  OAI22X1 instanceL2_g10559(.Y(instanceL2_n_11311), .A0(layer1_out[41]), .A1(
    layer1_out[40]), .B0(instanceL2_n_11341), .B1(instanceL2_n_11351));
  AOI21X1 instanceL2_g10560(.Y(instanceL2_n_11303), .A0(instanceL2_n_11337), .A1(
    layer1_out[41]), .B0(instanceL2_n_11332));
  OAI21X1 instanceL2_g10561(.Y(\instanceL2_prod_terms[5][4] [3]), .A0(
    instanceL2_n_11349), .A1(layer1_out[36]), .B0(instanceL2_n_11333));
  NOR2X1 instanceL2_g10562(.Y(instanceL2_n_11314), .A(layer1_out[43]), .B(
    layer1_out[40]));
  NAND2XL instanceL2_g10563(.Y(instanceL2_n_11315), .A(layer1_out[38]), .B(
    layer1_out[41]));
  NOR2X1 instanceL2_g10564(.Y(instanceL2_n_11316), .A(layer1_out[36]), .B(
    layer1_out[37]));
  NAND2XL instanceL2_g10565(.Y(instanceL2_n_11317), .A(layer1_out[43]), .B(
    layer1_out[40]));
  NOR2X1 instanceL2_g10566(.Y(instanceL2_n_11318), .A(layer1_out[38]), .B(
    layer1_out[41]));
  NAND2X1 instanceL2_g10567(.Y(instanceL2_n_11319), .A(layer1_out[42]), .B(
    layer1_out[40]));
  NOR2X1 instanceL2_g10568(.Y(instanceL2_n_11320), .A(layer1_out[43]), .B(
    layer1_out[41]));
  NAND2X1 instanceL2_g10569(.Y(instanceL2_n_11321), .A(layer1_out[43]), .B(
    layer1_out[41]));
  NOR2X1 instanceL2_g10570(.Y(instanceL2_n_11322), .A(instanceL2_n_11343), .B(
    instanceL2_n_11345));
  NAND2X1 instanceL2_g10571(.Y(instanceL2_n_11323), .A(layer1_out[38]), .B(
    layer1_out[36]));
  NOR2X1 instanceL2_g10572(.Y(instanceL2_n_11325), .A(layer1_out[39]), .B(
    layer1_out[42]));
  NAND2XL instanceL2_g10573(.Y(instanceL2_n_11326), .A(layer1_out[42]), .B(
    layer1_out[39]));
  NOR2XL instanceL2_g10574(.Y(instanceL2_n_11334), .A(layer1_out[40]), .B(
    instanceL2_n_11341));
  NAND2X1 instanceL2_g10575(.Y(instanceL2_n_11327), .A(layer1_out[38]), .B(
    layer1_out[40]));
  NOR2X1 instanceL2_g10576(.Y(instanceL2_n_11328), .A(layer1_out[38]), .B(
    layer1_out[40]));
  NOR2X1 instanceL2_g10577(.Y(instanceL2_n_11329), .A(layer1_out[42]), .B(
    layer1_out[40]));
  NAND2X1 instanceL2_g10578(.Y(instanceL2_n_11330), .A(instanceL2_n_11341), .B(
    instanceL2_n_11343));
  NAND2X1 instanceL2_g10579(.Y(instanceL2_n_11331), .A(layer1_out[41]), .B(
    layer1_out[39]));
  NOR2X1 instanceL2_g10580(.Y(instanceL2_n_11332), .A(instanceL2_n_11337), .B(
    layer1_out[41]));
  NAND2X1 instanceL2_g10581(.Y(instanceL2_n_11333), .A(instanceL2_n_11349), .B(
    layer1_out[36]));
  INVX1 instanceL2_g10582(.Y(instanceL2_n_11337), .A(layer1_out[42]));
  INVX1 instanceL2_g10583(.Y(instanceL2_n_11339), .A(layer1_out[38]));
  INVX1 instanceL2_g10584(.Y(instanceL2_n_11341), .A(layer1_out[41]));
  INVX1 instanceL2_g10585(.Y(instanceL2_n_11343), .A(layer1_out[39]));
  INVX1 instanceL2_g10586(.Y(instanceL2_n_11345), .A(layer1_out[36]));
  INVX1 instanceL2_g10587(.Y(instanceL2_n_11347), .A(layer1_out[43]));
  INVX1 instanceL2_g10588(.Y(instanceL2_n_11349), .A(layer1_out[37]));
  INVX1 instanceL2_g10589(.Y(instanceL2_n_11351), .A(layer1_out[40]));
  AOI21X1 instanceL2_g10353(.Y(\instanceL2_prod_terms[2][16] [10]), .A0(
    instanceL2_n_11780), .A1(instanceL2_n_11114), .B0(
    \instanceL2_prod_terms[2][16] [11]));
  NOR2X1 instanceL2_g10354(.Y(\instanceL2_prod_terms[2][16] [11]), .A(
    instanceL2_n_11780), .B(instanceL2_n_11114));
  AOI21X1 instanceL2_g10355(.Y(instanceL2_n_11114), .A0(instanceL2_n_11221), .A1(
    instanceL2_n_11118), .B0(instanceL2_n_11216));
  XNOR2X1 instanceL2_g10356(.Y(\instanceL2_prod_terms[2][16] [9]), .A(
    instanceL2_n_11760), .B(instanceL2_n_11118));
  OAI21X1 instanceL2_g10357(.Y(\instanceL2_prod_terms[1][16] [9]), .A0(
    instanceL2_n_11284), .A1(instanceL2_n_11124), .B0(instanceL2_n_11129));
  ADDFX1 instanceL2_g10358(.CO(instanceL2_n_11118), .S(
    \instanceL2_prod_terms[2][16] [8]), .A(instanceL2_n_11769), .B(
    instanceL2_n_11235), .CI(instanceL2_n_11126));
  AND2XL instanceL2_g10359(.Y(\instanceL2_prod_terms[1][16] [10]), .A(
    layer1_out[151]), .B(instanceL2_n_11129));
  AO21XL instanceL2_g10360(.Y(\instanceL2_prod_terms[1][16] [8]), .A0(
    layer1_out[149]), .A1(instanceL2_n_11131), .B0(instanceL2_n_11124));
  ADDFX1 instanceL2_g10361(.CO(instanceL2_n_11126), .S(
    \instanceL2_prod_terms[2][16] [7]), .A(instanceL2_n_11238), .B(
    instanceL2_n_11224), .CI(instanceL2_n_11136));
  NOR2X1 instanceL2_g10362(.Y(instanceL2_n_11124), .A(layer1_out[149]), .B(
    instanceL2_n_11131));
  NAND3BXL instanceL2_g10363(.Y(instanceL2_n_11129), .AN(instanceL2_n_11131), .B(
    instanceL2_n_11284), .C(instanceL2_n_11777));
  ADDFX1 instanceL2_g10364(.CO(instanceL2_n_11131), .S(
    \instanceL2_prod_terms[1][16] [7]), .A(instanceL2_n_11780), .B(
    layer1_out[148]), .CI(instanceL2_n_11142));
  AOI21X1 instanceL2_g10365(.Y(\instanceL2_prod_terms[0][16][7] ), .A0(
    layer1_out[151]), .A1(instanceL2_n_11145), .B0(instanceL2_n_11137));
  ADDFX1 instanceL2_g10366(.CO(instanceL2_n_11136), .S(
    \instanceL2_prod_terms[2][16] [6]), .A(instanceL2_n_11242), .B(
    instanceL2_n_11763), .CI(instanceL2_n_11147));
  INVX1 instanceL2_g10367(.Y(instanceL2_n_11137), .A(
    \instanceL2_prod_terms[0][16][13] ));
  OR2X1 instanceL2_g10368(.Y(\instanceL2_prod_terms[0][16][13] ), .A(
    layer1_out[151]), .B(instanceL2_n_11145));
  ADDFX1 instanceL2_g10369(.CO(instanceL2_n_11142), .S(
    \instanceL2_prod_terms[1][16] [6]), .A(instanceL2_n_11284), .B(
    layer1_out[147]), .CI(instanceL2_n_11152));
  OA21X1 instanceL2_g10370(.Y(\instanceL2_prod_terms[0][16][6] ), .A0(
    instanceL2_n_11284), .A1(instanceL2_n_11164), .B0(instanceL2_n_11145));
  MXI2XL instanceL2_g10371(.Y(\instanceL2_prod_terms[9][16] [10]), .A(
    instanceL2_n_11780), .B(layer1_out[151]), .S0(instanceL2_n_11155));
  ADDFX1 instanceL2_g10372(.CO(instanceL2_n_11147), .S(
    \instanceL2_prod_terms[2][16] [5]), .A(instanceL2_n_11241), .B(
    instanceL2_n_11212), .CI(instanceL2_n_11166));
  NAND2X1 instanceL2_g10373(.Y(instanceL2_n_11145), .A(instanceL2_n_11284), .B(
    instanceL2_n_11164));
  MX2XL instanceL2_g10374(.Y(\instanceL2_prod_terms[9][16] [9]), .A(
    layer1_out[150]), .B(instanceL2_n_11284), .S0(instanceL2_n_11157));
  ADDFX1 instanceL2_g10375(.CO(instanceL2_n_11152), .S(
    \instanceL2_prod_terms[1][16] [5]), .A(instanceL2_n_11777), .B(
    layer1_out[146]), .CI(instanceL2_n_11758));
  NOR2X1 instanceL2_g10376(.Y(\instanceL2_prod_terms[9][16] [11]), .A(
    instanceL2_n_11780), .B(instanceL2_n_11159));
  OAI21X1 instanceL2_g10377(.Y(instanceL2_n_11155), .A0(instanceL2_n_11284), .A1(
    instanceL2_n_11168), .B0(instanceL2_n_11217));
  AOI21X1 instanceL2_g10378(.Y(\instanceL2_prod_terms[0][16][5] ), .A0(
    layer1_out[149]), .A1(instanceL2_n_11759), .B0(instanceL2_n_11164));
  NAND2X1 instanceL2_g10379(.Y(instanceL2_n_11157), .A(instanceL2_n_11776), .B(
    instanceL2_n_11168));
  AOI21X1 instanceL2_g10380(.Y(instanceL2_n_11159), .A0(layer1_out[150]), .A1(
    instanceL2_n_11757), .B0(instanceL2_n_11216));
  ADDFX1 instanceL2_g10382(.CO(instanceL2_n_11166), .S(
    \instanceL2_prod_terms[2][16] [4]), .A(instanceL2_n_11232), .B(
    instanceL2_n_11764), .CI(instanceL2_n_11184));
  NOR2X1 instanceL2_g10383(.Y(instanceL2_n_11164), .A(layer1_out[149]), .B(
    instanceL2_n_11759));
  OAI2BB1X1 instanceL2_g10384(.Y(instanceL2_n_11168), .A0N(instanceL2_n_11780),
     .A1N(instanceL2_n_11777), .B0(instanceL2_n_11757));
  OAI21X1 instanceL2_g10386(.Y(instanceL2_n_11758), .A0(instanceL2_n_11774), .A1(
    instanceL2_n_11189), .B0(instanceL2_n_11773));
  OAI2BB1X1 instanceL2_g10387(.Y(instanceL2_n_11757), .A0N(instanceL2_n_11273),
     .A1N(instanceL2_n_11182), .B0(instanceL2_n_11277));
  XNOR2X1 instanceL2_g10388(.Y(\instanceL2_prod_terms[1][16] [4]), .A(
    instanceL2_n_11768), .B(instanceL2_n_11189));
  XNOR2X1 instanceL2_g10389(.Y(\instanceL2_prod_terms[9][16] [7]), .A(
    instanceL2_n_11766), .B(instanceL2_n_11182));
  OA21X1 instanceL2_g10390(.Y(\instanceL2_prod_terms[0][16][4] ), .A0(
    instanceL2_n_11779), .A1(instanceL2_n_11201), .B0(instanceL2_n_11759));
  MXI2XL instanceL2_g10391(.Y(\instanceL2_prod_terms[1][16] [3]), .A(
    instanceL2_n_11288), .B(layer1_out[144]), .S0(
    \instanceL2_prod_terms[0][16][3] ));
  ADDFX1 instanceL2_g10392(.CO(instanceL2_n_11184), .S(
    \instanceL2_prod_terms[2][16] [3]), .A(layer1_out[147]), .B(
    \instanceL2_prod_terms[9][16] [3]), .CI(instanceL2_n_11762));
  NAND2X1 instanceL2_g10393(.Y(instanceL2_n_11759), .A(instanceL2_n_11779), .B(
    instanceL2_n_11201));
  OAI21X1 instanceL2_g10394(.Y(instanceL2_n_11182), .A0(instanceL2_n_11775), .A1(
    instanceL2_n_11196), .B0(instanceL2_n_11276));
  XNOR2X1 instanceL2_g10395(.Y(\instanceL2_prod_terms[9][16] [6]), .A(
    instanceL2_n_11246), .B(instanceL2_n_11196));
  AOI21X1 instanceL2_g10396(.Y(instanceL2_n_11189), .A0(layer1_out[144]), .A1(
    instanceL2_n_11282), .B0(instanceL2_n_11201));
  XNOR2X1 instanceL2_g10397(.Y(\instanceL2_prod_terms[9][16] [5]), .A(
    instanceL2_n_11767), .B(instanceL2_n_11202));
  AOI221X1 instanceL2_g10398(.Y(instanceL2_n_11196), .A0(instanceL2_n_11771),
     .A1(instanceL2_n_11269), .B0(layer1_out[148]), .B1(layer1_out[146]), .C0(
    instanceL2_n_11761));
  XNOR2X1 instanceL2_g10399(.Y(\instanceL2_prod_terms[0][16][3] ), .A(
    instanceL2_n_11282), .B(instanceL2_n_11765));
  NOR2X1 instanceL2_g10400(.Y(instanceL2_n_11202), .A(instanceL2_n_11771), .B(
    instanceL2_n_11761));
  NAND2X1 instanceL2_g10401(.Y(instanceL2_n_11760), .A(instanceL2_n_11221), .B(
    instanceL2_n_11217));
  NOR2X1 instanceL2_g10402(.Y(instanceL2_n_11201), .A(layer1_out[147]), .B(
    instanceL2_n_11765));
  XNOR2X1 instanceL2_g10403(.Y(\instanceL2_prod_terms[9][16] [4]), .A(
    instanceL2_n_11232), .B(instanceL2_n_11249));
  XOR2XL instanceL2_g10404(.Y(\instanceL2_prod_terms[2][16] [2]), .A(
    instanceL2_n_11265), .B(instanceL2_n_11255));
  MXI2XL instanceL2_g10405(.Y(instanceL2_n_11212), .A(instanceL2_n_11777), .B(
    layer1_out[149]), .S0(instanceL2_n_11767));
  INVX1 instanceL2_g10406(.Y(instanceL2_n_11217), .A(instanceL2_n_11216));
  NOR2X1 instanceL2_g10407(.Y(instanceL2_n_11761), .A(instanceL2_n_11770), .B(
    instanceL2_n_11772));
  NAND2XL instanceL2_g10408(.Y(instanceL2_n_11762), .A(instanceL2_n_11265), .B(
    instanceL2_n_11262));
  NOR2X1 instanceL2_g10409(.Y(instanceL2_n_11216), .A(instanceL2_n_11284), .B(
    instanceL2_n_11776));
  MXI2XL instanceL2_g10410(.Y(instanceL2_n_11763), .A(instanceL2_n_11284), .B(
    layer1_out[150]), .S0(instanceL2_n_11246));
  MX2XL instanceL2_g10411(.Y(instanceL2_n_11224), .A(instanceL2_n_11780), .B(
    layer1_out[151]), .S0(instanceL2_n_11766));
  NAND2X1 instanceL2_g10412(.Y(instanceL2_n_11221), .A(instanceL2_n_11284), .B(
    instanceL2_n_11776));
  MXI2XL instanceL2_g10413(.Y(instanceL2_n_11764), .A(layer1_out[147]), .B(
    instanceL2_n_11282), .S0(instanceL2_n_11768));
  INVX1 instanceL2_g10414(.Y(instanceL2_n_11232), .A(instanceL2_n_11772));
  OA21X1 instanceL2_g10415(.Y(\instanceL2_prod_terms[0][16][2] ), .A0(
    instanceL2_n_11280), .A1(instanceL2_n_11264), .B0(instanceL2_n_11765));
  OAI2BB1X1 instanceL2_g10416(.Y(instanceL2_n_11235), .A0N(layer1_out[151]),
     .A1N(instanceL2_n_11273), .B0(instanceL2_n_11277));
  OAI21X1 instanceL2_g10417(.Y(instanceL2_n_11238), .A0(instanceL2_n_11284), .A1(
    instanceL2_n_11775), .B0(instanceL2_n_11276));
  OAI22X1 instanceL2_g10418(.Y(instanceL2_n_11241), .A0(instanceL2_n_11778), .A1(
    instanceL2_n_11268), .B0(instanceL2_n_11779), .B1(instanceL2_n_11282));
  OAI22X1 instanceL2_g10419(.Y(instanceL2_n_11242), .A0(instanceL2_n_11280), .A1(
    instanceL2_n_11278), .B0(instanceL2_n_11777), .B1(instanceL2_n_11779));
  NOR2BX1 instanceL2_g10420(.Y(\instanceL2_prod_terms[0][16][1] ), .AN(
    instanceL2_n_11265), .B(instanceL2_n_11264));
  OR2XL instanceL2_g10421(.Y(instanceL2_n_11249), .A(instanceL2_n_11771), .B(
    instanceL2_n_11770));
  NAND2X1 instanceL2_g10422(.Y(instanceL2_n_11765), .A(instanceL2_n_11280), .B(
    instanceL2_n_11264));
  NAND2X1 instanceL2_g10423(.Y(instanceL2_n_11766), .A(instanceL2_n_11277), .B(
    instanceL2_n_11273));
  NOR2BX1 instanceL2_g10424(.Y(instanceL2_n_11246), .AN(instanceL2_n_11276), .B(
    instanceL2_n_11775));
  OAI2BB1X1 instanceL2_g10425(.Y(instanceL2_n_11255), .A0N(instanceL2_n_11778),
     .A1N(instanceL2_n_11280), .B0(instanceL2_n_11262));
  AOI21X1 instanceL2_g10426(.Y(\instanceL2_prod_terms[9][16] [3]), .A0(
    instanceL2_n_11280), .A1(instanceL2_n_11288), .B0(instanceL2_n_11232));
  OAI22X1 instanceL2_g10427(.Y(instanceL2_n_11767), .A0(instanceL2_n_11779), .A1(
    layer1_out[146]), .B0(layer1_out[148]), .B1(instanceL2_n_11280));
  NOR2BX1 instanceL2_g10428(.Y(instanceL2_n_11768), .AN(instanceL2_n_11773), .B(
    instanceL2_n_11774));
  OAI22X1 instanceL2_g10429(.Y(instanceL2_n_11769), .A0(instanceL2_n_11780), .A1(
    layer1_out[149]), .B0(layer1_out[151]), .B1(instanceL2_n_11777));
  NOR2XL instanceL2_g10431(.Y(instanceL2_n_11268), .A(layer1_out[148]), .B(
    layer1_out[147]));
  NAND2X1 instanceL2_g10432(.Y(instanceL2_n_11269), .A(instanceL2_n_11779), .B(
    instanceL2_n_11280));
  NOR2X1 instanceL2_g10433(.Y(instanceL2_n_11770), .A(layer1_out[147]), .B(
    layer1_out[145]));
  NAND2X1 instanceL2_g10434(.Y(instanceL2_n_11262), .A(layer1_out[145]), .B(
    layer1_out[146]));
  NOR2X1 instanceL2_g10435(.Y(instanceL2_n_11771), .A(instanceL2_n_11282), .B(
    instanceL2_n_11778));
  NOR2X1 instanceL2_g10436(.Y(instanceL2_n_11264), .A(layer1_out[144]), .B(
    layer1_out[145]));
  NAND2XL instanceL2_g10437(.Y(instanceL2_n_11265), .A(layer1_out[144]), .B(
    layer1_out[145]));
  NAND2X1 instanceL2_g10438(.Y(instanceL2_n_11772), .A(layer1_out[144]), .B(
    layer1_out[146]));
  NOR2XL instanceL2_g10439(.Y(instanceL2_n_11278), .A(layer1_out[149]), .B(
    layer1_out[148]));
  NAND2X1 instanceL2_g10440(.Y(instanceL2_n_11773), .A(layer1_out[145]), .B(
    instanceL2_n_11779));
  NOR2X1 instanceL2_g10441(.Y(instanceL2_n_11774), .A(layer1_out[145]), .B(
    instanceL2_n_11779));
  NAND2X1 instanceL2_g10442(.Y(instanceL2_n_11273), .A(instanceL2_n_11284), .B(
    instanceL2_n_11779));
  NOR2X1 instanceL2_g10443(.Y(instanceL2_n_11775), .A(layer1_out[149]), .B(
    layer1_out[147]));
  NAND2X1 instanceL2_g10444(.Y(instanceL2_n_11776), .A(layer1_out[149]), .B(
    layer1_out[151]));
  NAND2X1 instanceL2_g10445(.Y(instanceL2_n_11276), .A(layer1_out[149]), .B(
    layer1_out[147]));
  NAND2X1 instanceL2_g10446(.Y(instanceL2_n_11277), .A(layer1_out[150]), .B(
    layer1_out[148]));
  INVX1 instanceL2_g10447(.Y(instanceL2_n_11280), .A(layer1_out[146]));
  INVX1 instanceL2_g10448(.Y(instanceL2_n_11282), .A(layer1_out[147]));
  INVX1 instanceL2_g10449(.Y(instanceL2_n_11284), .A(layer1_out[150]));
  INVX1 instanceL2_g10450(.Y(instanceL2_n_11777), .A(layer1_out[149]));
  INVX1 instanceL2_g10451(.Y(instanceL2_n_11288), .A(layer1_out[144]));
  INVX1 instanceL2_g10452(.Y(instanceL2_n_11778), .A(layer1_out[145]));
  INVX1 instanceL2_g10453(.Y(instanceL2_n_11779), .A(layer1_out[148]));
  INVX1 instanceL2_g10454(.Y(instanceL2_n_11780), .A(layer1_out[151]));
  CLKXOR2X1 instanceL2_g2(.Y(\instanceL2_prod_terms[9][16] [8]), .A(
    instanceL2_n_11769), .B(instanceL2_n_11757));
  INVX1 instanceL2_g10309(.Y(\instanceL2_prod_terms[1][14] [11]), .A(
    instanceL2_n_11073));
  AOI31X1 instanceL2_g10310(.Y(instanceL2_n_11073), .A0(instanceL2_n_11832), .A1(
    layer1_out[133]), .A2(instanceL2_n_11077), .B0(instanceL2_n_11113));
  MXI2XL instanceL2_g10311(.Y(\instanceL2_prod_terms[1][14] [10]), .A(
    layer1_out[132]), .B(instanceL2_n_11832), .S0(instanceL2_n_11077));
  OAI2BB1X1 instanceL2_g10312(.Y(instanceL2_n_11077), .A0N(instanceL2_n_11174),
     .A1N(instanceL2_n_11080), .B0(instanceL2_n_11792));
  XNOR2X1 instanceL2_g10313(.Y(\instanceL2_prod_terms[1][14] [9]), .A(
    instanceL2_n_11167), .B(instanceL2_n_11080));
  ADDFX1 instanceL2_g10314(.CO(instanceL2_n_11080), .S(
    \instanceL2_prod_terms[1][14] [8]), .A(instanceL2_n_11800), .B(
    instanceL2_n_11789), .CI(instanceL2_n_11083));
  ADDFX1 instanceL2_g10315(.CO(instanceL2_n_11083), .S(
    \instanceL2_prod_terms[1][14] [7]), .A(instanceL2_n_11188), .B(
    instanceL2_n_11185), .CI(instanceL2_n_11091));
  XNOR2X1 instanceL2_g10316(.Y(\instanceL2_prod_terms[8][14] [8]), .A(
    instanceL2_n_11790), .B(instanceL2_n_11086));
  ADDFX1 instanceL2_g10317(.CO(instanceL2_n_11086), .S(
    \instanceL2_prod_terms[8][14] [7]), .A(instanceL2_n_11824), .B(
    instanceL2_n_11793), .CI(instanceL2_n_11104));
  AOI21X1 instanceL2_g10318(.Y(\instanceL2_prod_terms[3][14] [9]), .A0(
    instanceL2_n_11285), .A1(instanceL2_n_11109), .B0(
    \instanceL2_prod_terms[3][14] [10]));
  ADDFX1 instanceL2_g10319(.CO(instanceL2_n_11091), .S(
    \instanceL2_prod_terms[1][14] [6]), .A(instanceL2_n_11791), .B(
    instanceL2_n_11787), .CI(instanceL2_n_11111));
  NOR2X1 instanceL2_g10320(.Y(\instanceL2_prod_terms[3][14] [10]), .A(
    instanceL2_n_11285), .B(instanceL2_n_11109));
  OAI21X1 instanceL2_g10321(.Y(\instanceL2_prod_terms[8][14] [9]), .A0(
    instanceL2_n_11285), .A1(instanceL2_n_11781), .B0(instanceL2_n_11096));
  INVX1 instanceL2_g10322(.Y(instanceL2_n_11096), .A(instanceL2_n_11113));
  AOI2BB1X1 instanceL2_g10323(.Y(\instanceL2_prod_terms[0][14][8] ), .A0N(
    layer1_out[133]), .A1N(instanceL2_n_11781), .B0(
    \instanceL2_prod_terms[0][14][9] ));
  ADDFX1 instanceL2_g10324(.CO(instanceL2_n_11104), .S(
    \instanceL2_prod_terms[8][14] [6]), .A(instanceL2_n_11826), .B(
    instanceL2_n_11796), .CI(instanceL2_n_11127));
  OA21X1 instanceL2_g10325(.Y(\instanceL2_prod_terms[3][14] [8]), .A0(
    layer1_out[132]), .A1(instanceL2_n_11117), .B0(instanceL2_n_11109));
  AND2X1 instanceL2_g10326(.Y(\instanceL2_prod_terms[0][14][9] ), .A(
    instanceL2_n_11781), .B(layer1_out[133]));
  AO21X1 instanceL2_g10327(.Y(\instanceL2_prod_terms[4][14] [7]), .A0(
    layer1_out[133]), .A1(instanceL2_n_11783), .B0(instanceL2_n_11113));
  XNOR2X1 instanceL2_g10328(.Y(\instanceL2_prod_terms[0][14][7] ), .A(
    instanceL2_n_11801), .B(instanceL2_n_11782));
  ADDFX1 instanceL2_g10329(.CO(instanceL2_n_11111), .S(
    \instanceL2_prod_terms[1][14] [5]), .A(instanceL2_n_11810), .B(
    instanceL2_n_11178), .CI(instanceL2_n_11133));
  NAND2X1 instanceL2_g10330(.Y(instanceL2_n_11109), .A(layer1_out[132]), .B(
    instanceL2_n_11117));
  NOR2X1 instanceL2_g10331(.Y(instanceL2_n_11113), .A(layer1_out[133]), .B(
    instanceL2_n_11783));
  OAI211X1 instanceL2_g10332(.Y(instanceL2_n_11781), .A0(instanceL2_n_11823),
     .A1(instanceL2_n_11125), .B0(instanceL2_n_11822), .C0(instanceL2_n_11270));
  NAND2X1 instanceL2_g10333(.Y(instanceL2_n_11782), .A(instanceL2_n_11822), .B(
    instanceL2_n_11125));
  OAI21X1 instanceL2_g10334(.Y(instanceL2_n_11117), .A0(instanceL2_n_11807), .A1(
    instanceL2_n_11784), .B0(instanceL2_n_11251));
  XNOR2X1 instanceL2_g10335(.Y(\instanceL2_prod_terms[0][14][6] ), .A(
    instanceL2_n_11799), .B(instanceL2_n_11138));
  CLKXOR2X1 instanceL2_g10336(.Y(\instanceL2_prod_terms[3][14] [7]), .A(
    instanceL2_n_11793), .B(instanceL2_n_11784));
  ADDFX1 instanceL2_g10337(.CO(instanceL2_n_11127), .S(
    \instanceL2_prod_terms[8][14] [5]), .A(instanceL2_n_11825), .B(
    instanceL2_n_11211), .CI(instanceL2_n_11151));
  NAND2X1 instanceL2_g10338(.Y(instanceL2_n_11125), .A(instanceL2_n_11821), .B(
    instanceL2_n_11138));
  XNOR2X1 instanceL2_g10339(.Y(\instanceL2_prod_terms[0][14][5] ), .A(
    instanceL2_n_11209), .B(instanceL2_n_11144));
  MX2XL instanceL2_g10340(.Y(\instanceL2_prod_terms[4][14] [6]), .A(
    layer1_out[132]), .B(instanceL2_n_11832), .S0(instanceL2_n_11785));
  ADDFX1 instanceL2_g10341(.CO(instanceL2_n_11133), .S(
    \instanceL2_prod_terms[1][14] [4]), .A(layer1_out[130]), .B(
    instanceL2_n_11803), .CI(instanceL2_n_11158));
  NOR2X1 instanceL2_g10343(.Y(instanceL2_n_11783), .A(layer1_out[132]), .B(
    instanceL2_n_11785));
  XNOR2X1 instanceL2_g10344(.Y(\instanceL2_prod_terms[3][14] [6]), .A(
    instanceL2_n_11796), .B(instanceL2_n_11149));
  AOI21X1 instanceL2_g10345(.Y(instanceL2_n_11784), .A0(instanceL2_n_11819), .A1(
    instanceL2_n_11149), .B0(instanceL2_n_11820));
  OAI22X1 instanceL2_g10346(.Y(instanceL2_n_11138), .A0(instanceL2_n_11259), .A1(
    instanceL2_n_11148), .B0(instanceL2_n_11831), .B1(instanceL2_n_11811));
  NAND2X1 instanceL2_g10348(.Y(instanceL2_n_11144), .A(instanceL2_n_11818), .B(
    instanceL2_n_11148));
  XNOR2X1 instanceL2_g10349(.Y(\instanceL2_prod_terms[0][14][4] ), .A(
    instanceL2_n_11228), .B(instanceL2_n_11158));
  ADDFX1 instanceL2_g10350(.CO(instanceL2_n_11151), .S(
    \instanceL2_prod_terms[8][14] [4]), .A(instanceL2_n_11828), .B(
    instanceL2_n_11797), .CI(instanceL2_n_11788));
  NAND2X1 instanceL2_g10351(.Y(instanceL2_n_11148), .A(instanceL2_n_11817), .B(
    instanceL2_n_11158));
  OAI21X1 instanceL2_g10352(.Y(instanceL2_n_11149), .A0(instanceL2_n_11811), .A1(
    instanceL2_n_11786), .B0(instanceL2_n_11247));
  OA21X1 instanceL2_g10590(.Y(\instanceL2_prod_terms[4][14] [5]), .A0(
    instanceL2_n_11281), .A1(instanceL2_n_11187), .B0(instanceL2_n_11785));
  CLKXOR2X1 instanceL2_g10591(.Y(\instanceL2_prod_terms[3][14] [5]), .A(
    instanceL2_n_11211), .B(instanceL2_n_11786));
  NAND2X1 instanceL2_g10592(.Y(instanceL2_n_11785), .A(instanceL2_n_11281), .B(
    instanceL2_n_11187));
  OAI2BB1X1 instanceL2_g10593(.Y(instanceL2_n_11158), .A0N(instanceL2_n_11812),
     .A1N(instanceL2_n_11175), .B0(instanceL2_n_11267));
  XNOR2X1 instanceL2_g10594(.Y(\instanceL2_prod_terms[0][14][3] ), .A(
    instanceL2_n_11175), .B(instanceL2_n_11795));
  XNOR2X1 instanceL2_g10595(.Y(\instanceL2_prod_terms[8][14] [3]), .A(
    instanceL2_n_11814), .B(instanceL2_n_11296));
  MX2X1 instanceL2_g10596(.Y(\instanceL2_prod_terms[4][14] [3]), .A(
    layer1_out[129]), .B(instanceL2_n_11829), .S0(instanceL2_n_11208));
  NAND2X1 instanceL2_g10597(.Y(instanceL2_n_11167), .A(instanceL2_n_11174), .B(
    instanceL2_n_11792));
  AOI21X1 instanceL2_g10598(.Y(instanceL2_n_11786), .A0(instanceL2_n_11816), .A1(
    instanceL2_n_11186), .B0(instanceL2_n_11815));
  XNOR2X1 instanceL2_g10599(.Y(\instanceL2_prod_terms[3][14] [4]), .A(
    instanceL2_n_11797), .B(instanceL2_n_11186));
  CLKXOR2X1 instanceL2_g10600(.Y(\instanceL2_prod_terms[0][14][2] ), .A(
    instanceL2_n_11260), .B(instanceL2_n_11802));
  AOI21X1 instanceL2_g10601(.Y(\instanceL2_prod_terms[4][14] [4]), .A0(
    layer1_out[130]), .A1(instanceL2_n_11206), .B0(instanceL2_n_11187));
  OAI21XL instanceL2_g10602(.Y(instanceL2_n_11174), .A0(instanceL2_n_11285), .A1(
    layer1_out[130]), .B0(layer1_out[131]));
  MXI2XL instanceL2_g10603(.Y(instanceL2_n_11178), .A(instanceL2_n_11287), .B(
    layer1_out[127]), .S0(instanceL2_n_11209));
  NAND2XL instanceL2_g10604(.Y(instanceL2_n_11175), .A(instanceL2_n_11809), .B(
    instanceL2_n_11260));
  XNOR2X1 instanceL2_g10605(.Y(\instanceL2_prod_terms[3][14] [3]), .A(
    instanceL2_n_11813), .B(instanceL2_n_11794));
  MXI2XL instanceL2_g10606(.Y(instanceL2_n_11787), .A(instanceL2_n_11281), .B(
    layer1_out[131]), .S0(instanceL2_n_11798));
  MXI2XL instanceL2_g10607(.Y(instanceL2_n_11185), .A(layer1_out[132]), .B(
    instanceL2_n_11832), .S0(instanceL2_n_11804));
  OAI2BB1X1 instanceL2_g10608(.Y(instanceL2_n_11188), .A0N(instanceL2_n_11830),
     .A1N(instanceL2_n_11821), .B0(instanceL2_n_11822));
  AOI21X1 instanceL2_g10609(.Y(instanceL2_n_11186), .A0(instanceL2_n_11806), .A1(
    instanceL2_n_11813), .B0(instanceL2_n_11805));
  NOR2X1 instanceL2_g10610(.Y(instanceL2_n_11187), .A(layer1_out[130]), .B(
    instanceL2_n_11206));
  AOI2BB1X1 instanceL2_g10611(.Y(instanceL2_n_11788), .A0N(layer1_out[128]),
     .A1N(instanceL2_n_11814), .B0(instanceL2_n_11794));
  OA21X1 instanceL2_g10612(.Y(\instanceL2_prod_terms[4][14] [2]), .A0(
    instanceL2_n_11830), .A1(instanceL2_n_11257), .B0(instanceL2_n_11208));
  OAI21X1 instanceL2_g10613(.Y(instanceL2_n_11789), .A0(layer1_out[129]), .A1(
    instanceL2_n_11823), .B0(instanceL2_n_11270));
  MXI2XL instanceL2_g10614(.Y(instanceL2_n_11790), .A(instanceL2_n_11832), .B(
    layer1_out[132]), .S0(instanceL2_n_11827));
  OAI21X1 instanceL2_g10615(.Y(instanceL2_n_11791), .A0(layer1_out[127]), .A1(
    instanceL2_n_11259), .B0(instanceL2_n_11808));
  NOR2BX1 instanceL2_g10381(.Y(\instanceL2_prod_terms[4][14] [1]), .AN(
    instanceL2_n_11260), .B(instanceL2_n_11257));
  NOR2BX1 instanceL2_g10616(.Y(\instanceL2_prod_terms[3][14] [2]), .AN(
    instanceL2_n_11813), .B(instanceL2_n_11814));
  NAND2BX1 instanceL2_g10617(.Y(instanceL2_n_11206), .AN(instanceL2_n_11812), .B(
    instanceL2_n_11257));
  NAND2X1 instanceL2_g10618(.Y(instanceL2_n_11792), .A(layer1_out[133]), .B(
    instanceL2_n_11259));
  NAND2XL instanceL2_g10385(.Y(instanceL2_n_11795), .A(instanceL2_n_11267), .B(
    instanceL2_n_11812));
  NAND2X1 instanceL2_g10619(.Y(instanceL2_n_11208), .A(instanceL2_n_11830), .B(
    instanceL2_n_11257));
  NAND2BX1 instanceL2_g10620(.Y(instanceL2_n_11209), .AN(instanceL2_n_11259), .B(
    instanceL2_n_11808));
  NAND2BX1 instanceL2_g10621(.Y(instanceL2_n_11793), .AN(instanceL2_n_11807), .B(
    instanceL2_n_11251));
  NAND2BX1 instanceL2_g10622(.Y(instanceL2_n_11211), .AN(instanceL2_n_11811), .B(
    instanceL2_n_11247));
  NOR2BX1 instanceL2_g10623(.Y(instanceL2_n_11794), .AN(instanceL2_n_11806), .B(
    instanceL2_n_11805));
  NAND2XL instanceL2_g10624(.Y(instanceL2_n_11228), .A(instanceL2_n_11818), .B(
    instanceL2_n_11817));
  OAI22X1 instanceL2_g10625(.Y(instanceL2_n_11798), .A0(layer1_out[132]), .A1(
    layer1_out[128]), .B0(instanceL2_n_11832), .B1(instanceL2_n_11830));
  NAND2XL instanceL2_g10626(.Y(instanceL2_n_11799), .A(instanceL2_n_11822), .B(
    instanceL2_n_11821));
  OAI22X1 instanceL2_g10627(.Y(instanceL2_n_11800), .A0(layer1_out[133]), .A1(
    layer1_out[130]), .B0(instanceL2_n_11285), .B1(instanceL2_n_11831));
  NAND2BX1 instanceL2_g10628(.Y(instanceL2_n_11801), .AN(instanceL2_n_11823), .B(
    instanceL2_n_11270));
  OAI2BB1X1 instanceL2_g10629(.Y(instanceL2_n_11802), .A0N(instanceL2_n_11287),
     .A1N(instanceL2_n_11830), .B0(instanceL2_n_11809));
  OAI21X1 instanceL2_g10630(.Y(instanceL2_n_11803), .A0(layer1_out[126]), .A1(
    instanceL2_n_11829), .B0(instanceL2_n_11810));
  AOI22X1 instanceL2_g10631(.Y(instanceL2_n_11804), .A0(instanceL2_n_11285), .A1(
    instanceL2_n_11829), .B0(layer1_out[133]), .B1(layer1_out[129]));
  NAND2BX1 instanceL2_g10632(.Y(instanceL2_n_11796), .AN(instanceL2_n_11820), .B(
    instanceL2_n_11819));
  NAND2BX1 instanceL2_g10633(.Y(instanceL2_n_11797), .AN(instanceL2_n_11815), .B(
    instanceL2_n_11816));
  NAND2XL instanceL2_g10634(.Y(instanceL2_n_11247), .A(layer1_out[131]), .B(
    layer1_out[129]));
  NOR2X1 instanceL2_g10635(.Y(instanceL2_n_11805), .A(layer1_out[129]), .B(
    layer1_out[127]));
  NAND2X1 instanceL2_g10636(.Y(instanceL2_n_11806), .A(layer1_out[127]), .B(
    layer1_out[129]));
  NOR2XL instanceL2_g10637(.Y(instanceL2_n_11807), .A(layer1_out[133]), .B(
    layer1_out[131]));
  NAND2X1 instanceL2_g10638(.Y(instanceL2_n_11251), .A(layer1_out[133]), .B(
    layer1_out[131]));
  NAND2X1 instanceL2_g10639(.Y(instanceL2_n_11808), .A(layer1_out[130]), .B(
    layer1_out[131]));
  NAND2X1 instanceL2_g10640(.Y(instanceL2_n_11809), .A(layer1_out[127]), .B(
    layer1_out[128]));
  NAND2X1 instanceL2_g10641(.Y(instanceL2_n_11810), .A(layer1_out[126]), .B(
    instanceL2_n_11829));
  NOR2X1 instanceL2_g10642(.Y(instanceL2_n_11811), .A(layer1_out[131]), .B(
    layer1_out[129]));
  NAND2X1 instanceL2_g10643(.Y(instanceL2_n_11812), .A(instanceL2_n_11830), .B(
    instanceL2_n_11829));
  NOR2X1 instanceL2_g10644(.Y(instanceL2_n_11257), .A(layer1_out[126]), .B(
    layer1_out[127]));
  NAND2X1 instanceL2_g10645(.Y(instanceL2_n_11813), .A(layer1_out[128]), .B(
    layer1_out[126]));
  NOR2X1 instanceL2_g10646(.Y(instanceL2_n_11259), .A(layer1_out[130]), .B(
    layer1_out[131]));
  NAND2X1 instanceL2_g10647(.Y(instanceL2_n_11260), .A(layer1_out[126]), .B(
    layer1_out[127]));
  NOR2XL instanceL2_g10648(.Y(instanceL2_n_11814), .A(layer1_out[126]), .B(
    layer1_out[128]));
  NOR2XL instanceL2_g10649(.Y(instanceL2_n_11824), .A(layer1_out[130]), .B(
    instanceL2_n_11832));
  NOR2XL instanceL2_g10650(.Y(instanceL2_n_11815), .A(instanceL2_n_11831), .B(
    instanceL2_n_11830));
  NAND2X1 instanceL2_g10651(.Y(instanceL2_n_11816), .A(instanceL2_n_11831), .B(
    instanceL2_n_11830));
  NAND2X1 instanceL2_g10652(.Y(instanceL2_n_11817), .A(instanceL2_n_11831), .B(
    instanceL2_n_11829));
  NAND2XL instanceL2_g10653(.Y(instanceL2_n_11818), .A(layer1_out[130]), .B(
    layer1_out[129]));
  NAND2X1 instanceL2_g10654(.Y(instanceL2_n_11267), .A(layer1_out[128]), .B(
    layer1_out[129]));
  NOR2X1 instanceL2_g10655(.Y(instanceL2_n_11825), .A(instanceL2_n_11831), .B(
    layer1_out[128]));
  NAND2X1 instanceL2_g10656(.Y(instanceL2_n_11819), .A(instanceL2_n_11832), .B(
    instanceL2_n_11831));
  NOR2XL instanceL2_g10657(.Y(instanceL2_n_11820), .A(instanceL2_n_11832), .B(
    instanceL2_n_11831));
  NOR2XL instanceL2_g10658(.Y(instanceL2_n_11826), .A(layer1_out[129]), .B(
    instanceL2_n_11281));
  NOR2X1 instanceL2_g10659(.Y(instanceL2_n_11827), .A(instanceL2_n_11285), .B(
    layer1_out[131]));
  NOR2X1 instanceL2_g10660(.Y(instanceL2_n_11828), .A(layer1_out[127]), .B(
    instanceL2_n_11829));
  NAND2XL instanceL2_g10661(.Y(instanceL2_n_11270), .A(layer1_out[133]), .B(
    layer1_out[132]));
  NAND2X1 instanceL2_g10662(.Y(instanceL2_n_11821), .A(instanceL2_n_11832), .B(
    instanceL2_n_11281));
  NAND2X1 instanceL2_g10430(.Y(instanceL2_n_11822), .A(layer1_out[131]), .B(
    layer1_out[132]));
  NOR2X1 instanceL2_g10663(.Y(instanceL2_n_11823), .A(layer1_out[132]), .B(
    layer1_out[133]));
  INVX1 instanceL2_g10664(.Y(instanceL2_n_11281), .A(layer1_out[131]));
  INVX1 instanceL2_g10665(.Y(instanceL2_n_11829), .A(layer1_out[129]));
  INVX1 instanceL2_g10666(.Y(instanceL2_n_11285), .A(layer1_out[133]));
  INVX1 instanceL2_g10667(.Y(instanceL2_n_11287), .A(layer1_out[127]));
  INVX1 instanceL2_g10668(.Y(instanceL2_n_11830), .A(layer1_out[128]));
  INVX1 instanceL2_g10669(.Y(instanceL2_n_11831), .A(layer1_out[130]));
  INVX1 instanceL2_g10670(.Y(instanceL2_n_11832), .A(layer1_out[132]));
  NAND2BX2 instanceL2_g10671(.Y(\instanceL2_prod_terms[4][14] [13]), .AN(
    instanceL2_n_11785), .B(instanceL2_n_11823));
  XOR2XL instanceL2_g10672(.Y(instanceL2_n_11296), .A(layer1_out[128]), .B(
    instanceL2_n_11794));
  OAI2BB1X1 instanceL2_g10673(.Y(\instanceL2_prod_terms[2][11][11] ), .A0N(
    layer1_out[106]), .A1N(instanceL2_n_11833), .B0(instanceL2_n_11851));
  ADDFX1 instanceL2_g10674(.CO(instanceL2_n_11833), .S(
    \instanceL2_prod_terms[2][11][10] ), .A(instanceL2_n_11392), .B(
    instanceL2_n_11380), .CI(instanceL2_n_11191));
  ADDFX1 instanceL2_g10675(.CO(instanceL2_n_11191), .S(
    \instanceL2_prod_terms[2][11][9] ), .A(instanceL2_n_11382), .B(
    instanceL2_n_11868), .CI(instanceL2_n_11193));
  ADDFX1 instanceL2_g10676(.CO(instanceL2_n_11193), .S(
    \instanceL2_prod_terms[2][11][8] ), .A(instanceL2_n_11866), .B(
    instanceL2_n_11861), .CI(instanceL2_n_11195));
  ADDFX1 instanceL2_g10677(.CO(instanceL2_n_11195), .S(
    \instanceL2_prod_terms[2][11][7] ), .A(instanceL2_n_11324), .B(
    instanceL2_n_11403), .CI(instanceL2_n_11834));
  XNOR2X1 instanceL2_g10678(.Y(\instanceL2_prod_terms[4][11] [9]), .A(
    layer1_out[106]), .B(instanceL2_n_11837));
  XNOR2X1 instanceL2_g10679(.Y(\instanceL2_prod_terms[0][11][6] ), .A(
    layer1_out[105]), .B(instanceL2_n_11229));
  XNOR2X1 instanceL2_g10680(.Y(\instanceL2_prod_terms[8][11] [10]), .A(
    instanceL2_n_11392), .B(instanceL2_n_11835));
  ADDFX1 instanceL2_g10681(.CO(instanceL2_n_11834), .S(
    \instanceL2_prod_terms[2][11][6] ), .A(instanceL2_n_11864), .B(
    instanceL2_n_11859), .CI(instanceL2_n_11839));
  NAND2X1 instanceL2_g10682(.Y(\instanceL2_prod_terms[8][11] [11]), .A(
    instanceL2_n_11851), .B(instanceL2_n_11836));
  OAI21X1 instanceL2_g10683(.Y(\instanceL2_prod_terms[6][11] [9]), .A0(
    layer1_out[106]), .A1(instanceL2_n_11838), .B0(instanceL2_n_11836));
  NOR2X1 instanceL2_g10684(.Y(instanceL2_n_11835), .A(instanceL2_n_11380), .B(
    instanceL2_n_11223));
  OA21X1 instanceL2_g10685(.Y(\instanceL2_prod_terms[4][11] [8]), .A0(
    layer1_out[105]), .A1(instanceL2_n_11840), .B0(instanceL2_n_11837));
  OAI21X1 instanceL2_g10686(.Y(\instanceL2_prod_terms[6][11] [10]), .A0(
    instanceL2_n_11388), .A1(instanceL2_n_11838), .B0(instanceL2_n_11367));
  XNOR2X1 instanceL2_g10687(.Y(\instanceL2_prod_terms[8][11] [9]), .A(
    instanceL2_n_11868), .B(instanceL2_n_11230));
  NOR2BX1 instanceL2_g10688(.Y(\instanceL2_prod_terms[4][11] [10]), .AN(
    instanceL2_n_11840), .B(instanceL2_n_11367));
  NAND3X1 instanceL2_g10689(.Y(instanceL2_n_11836), .A(layer1_out[106]), .B(
    instanceL2_n_11367), .C(instanceL2_n_11838));
  NAND2X1 instanceL2_g10690(.Y(instanceL2_n_11837), .A(layer1_out[105]), .B(
    instanceL2_n_11840));
  AOI21X1 instanceL2_g10691(.Y(\instanceL2_prod_terms[0][11][5] ), .A0(
    layer1_out[104]), .A1(instanceL2_n_11847), .B0(instanceL2_n_11229));
  AOI21X1 instanceL2_g10692(.Y(instanceL2_n_11223), .A0(instanceL2_n_11388), .A1(
    layer1_out[104]), .B0(instanceL2_n_11230));
  XNOR2X1 instanceL2_g10693(.Y(\instanceL2_prod_terms[6][11] [8]), .A(
    instanceL2_n_11338), .B(instanceL2_n_11841));
  ADDFX1 instanceL2_g10694(.CO(instanceL2_n_11839), .S(
    \instanceL2_prod_terms[2][11][5] ), .A(instanceL2_n_11368), .B(
    instanceL2_n_11860), .CI(instanceL2_n_11846));
  NAND2X1 instanceL2_g10695(.Y(instanceL2_n_11838), .A(instanceL2_n_11359), .B(
    instanceL2_n_11841));
  NOR2X1 instanceL2_g10696(.Y(instanceL2_n_11229), .A(layer1_out[104]), .B(
    instanceL2_n_11847));
  AOI21X1 instanceL2_g10697(.Y(instanceL2_n_11230), .A0(instanceL2_n_11386), .A1(
    instanceL2_n_11844), .B0(instanceL2_n_11382));
  MXI2XL instanceL2_g10698(.Y(\instanceL2_prod_terms[8][11] [8]), .A(
    instanceL2_n_11867), .B(instanceL2_n_11866), .S0(instanceL2_n_11844));
  XNOR2X1 instanceL2_g10699(.Y(\instanceL2_prod_terms[4][11] [7]), .A(
    instanceL2_n_11868), .B(instanceL2_n_11842));
  XNOR2X1 instanceL2_g10700(.Y(\instanceL2_prod_terms[6][11] [7]), .A(
    instanceL2_n_11340), .B(instanceL2_n_11843));
  OAI2BB1X1 instanceL2_g10701(.Y(instanceL2_n_11840), .A0N(instanceL2_n_11360),
     .A1N(instanceL2_n_11842), .B0(instanceL2_n_11363));
  OAI211X1 instanceL2_g10702(.Y(instanceL2_n_11841), .A0(instanceL2_n_11364),
     .A1(instanceL2_n_11845), .B0(instanceL2_n_11362), .C0(instanceL2_n_11357));
  OA21X1 instanceL2_g10703(.Y(\instanceL2_prod_terms[0][11][4] ), .A0(
    instanceL2_n_11390), .A1(instanceL2_n_11855), .B0(instanceL2_n_11847));
  NAND2X1 instanceL2_g10704(.Y(instanceL2_n_11843), .A(instanceL2_n_11362), .B(
    instanceL2_n_11845));
  OAI21X1 instanceL2_g10705(.Y(instanceL2_n_11842), .A0(instanceL2_n_11377), .A1(
    instanceL2_n_11848), .B0(instanceL2_n_11373));
  XNOR2X1 instanceL2_g10706(.Y(\instanceL2_prod_terms[8][11] [7]), .A(
    instanceL2_n_11870), .B(instanceL2_n_11849));
  MXI2XL instanceL2_g10707(.Y(\instanceL2_prod_terms[4][11] [6]), .A(
    instanceL2_n_11867), .B(instanceL2_n_11866), .S0(instanceL2_n_11848));
  XNOR2X1 instanceL2_g10708(.Y(\instanceL2_prod_terms[6][11] [6]), .A(
    instanceL2_n_11336), .B(instanceL2_n_11850));
  OAI2BB1X1 instanceL2_g10709(.Y(instanceL2_n_11844), .A0N(instanceL2_n_11375),
     .A1N(instanceL2_n_11849), .B0(instanceL2_n_11374));
  ADDFX1 instanceL2_g10710(.CO(instanceL2_n_11846), .S(
    \instanceL2_prod_terms[2][11][4] ), .A(layer1_out[103]), .B(
    \instanceL2_prod_terms[2][11][2] ), .CI(instanceL2_n_11862));
  NAND2X1 instanceL2_g10711(.Y(instanceL2_n_11845), .A(instanceL2_n_11358), .B(
    instanceL2_n_11850));
  XNOR2X1 instanceL2_g10712(.Y(\instanceL2_prod_terms[6][11] [5]), .A(
    instanceL2_n_11871), .B(instanceL2_n_11852));
  NAND2X1 instanceL2_g10713(.Y(instanceL2_n_11847), .A(instanceL2_n_11390), .B(
    instanceL2_n_11855));
  OAI21X1 instanceL2_g10714(.Y(\instanceL2_prod_terms[0][11][7] ), .A0(
    instanceL2_n_11388), .A1(instanceL2_n_11854), .B0(instanceL2_n_11851));
  AOI22X1 instanceL2_g10715(.Y(instanceL2_n_11848), .A0(instanceL2_n_11385), .A1(
    instanceL2_n_11857), .B0(layer1_out[102]), .B1(layer1_out[104]));
  OAI21X1 instanceL2_g10716(.Y(instanceL2_n_11849), .A0(instanceL2_n_11381), .A1(
    instanceL2_n_11856), .B0(instanceL2_n_11378));
  XOR2XL instanceL2_g10717(.Y(\instanceL2_prod_terms[4][11] [5]), .A(
    instanceL2_n_11870), .B(instanceL2_n_11857));
  XNOR2X1 instanceL2_g10718(.Y(\instanceL2_prod_terms[8][11] [6]), .A(
    instanceL2_n_11869), .B(instanceL2_n_11856));
  OAI22X1 instanceL2_g10719(.Y(instanceL2_n_11850), .A0(instanceL2_n_11379), .A1(
    instanceL2_n_11853), .B0(instanceL2_n_11394), .B1(instanceL2_n_11376));
  OR2X1 instanceL2_g10720(.Y(\instanceL2_prod_terms[0][11][13] ), .A(
    layer1_out[106]), .B(instanceL2_n_11854));
  NAND2X1 instanceL2_g10721(.Y(instanceL2_n_11851), .A(instanceL2_n_11388), .B(
    instanceL2_n_11854));
  AOI21X1 instanceL2_g10722(.Y(\instanceL2_prod_terms[0][11][3] ), .A0(
    layer1_out[102]), .A1(instanceL2_n_11865), .B0(instanceL2_n_11855));
  XNOR2X1 instanceL2_g10723(.Y(\instanceL2_prod_terms[6][11] [4]), .A(
    instanceL2_n_11858), .B(instanceL2_n_11348));
  OAI2BB1X1 instanceL2_g10724(.Y(instanceL2_n_11852), .A0N(layer1_out[101]),
     .A1N(layer1_out[102]), .B0(instanceL2_n_11853));
  OAI21X1 instanceL2_g10725(.Y(instanceL2_n_11853), .A0(layer1_out[101]), .A1(
    layer1_out[102]), .B0(instanceL2_n_11858));
  NAND3BXL instanceL2_g10726(.Y(instanceL2_n_11854), .AN(instanceL2_n_11865), .B(
    instanceL2_n_11364), .C(instanceL2_n_11379));
  NOR2X1 instanceL2_g10727(.Y(instanceL2_n_11855), .A(layer1_out[102]), .B(
    instanceL2_n_11865));
  AOI21X1 instanceL2_g10728(.Y(instanceL2_n_11856), .A0(instanceL2_n_11383), .A1(
    instanceL2_n_11368), .B0(instanceL2_n_11384));
  XNOR2X1 instanceL2_g10729(.Y(\instanceL2_prod_terms[8][11] [5]), .A(
    instanceL2_n_11368), .B(instanceL2_n_11346));
  XNOR2X1 instanceL2_g10730(.Y(\instanceL2_prod_terms[4][11] [4]), .A(
    instanceL2_n_11869), .B(instanceL2_n_11862));
  XOR2XL instanceL2_g10731(.Y(\instanceL2_prod_terms[6][11] [3]), .A(
    instanceL2_n_11366), .B(instanceL2_n_11872));
  OAI22X1 instanceL2_g10732(.Y(instanceL2_n_11857), .A0(instanceL2_n_11376), .A1(
    instanceL2_n_11863), .B0(instanceL2_n_11390), .B1(instanceL2_n_11402));
  XNOR2X1 instanceL2_g10733(.Y(\instanceL2_prod_terms[4][11] [3]), .A(
    instanceL2_n_11365), .B(instanceL2_n_11346));
  NAND2XL instanceL2_g10734(.Y(instanceL2_n_11858), .A(instanceL2_n_11356), .B(
    instanceL2_n_11366));
  OAI22X1 instanceL2_g10735(.Y(instanceL2_n_11859), .A0(instanceL2_n_11402), .A1(
    instanceL2_n_11866), .B0(layer1_out[101]), .B1(instanceL2_n_11867));
  XNOR2X1 instanceL2_g10736(.Y(instanceL2_n_11860), .A(layer1_out[100]), .B(
    instanceL2_n_11870));
  OA21X1 instanceL2_g10737(.Y(\instanceL2_prod_terms[0][11][2] ), .A0(
    instanceL2_n_11402), .A1(instanceL2_n_11361), .B0(instanceL2_n_11865));
  OAI2BB1X1 instanceL2_g10738(.Y(instanceL2_n_11861), .A0N(instanceL2_n_11394),
     .A1N(instanceL2_n_11360), .B0(instanceL2_n_11363));
  INVX1 instanceL2_g10739(.Y(instanceL2_n_11863), .A(instanceL2_n_11862));
  AO21XL instanceL2_g10740(.Y(instanceL2_n_11864), .A0(layer1_out[104]), .A1(
    instanceL2_n_11383), .B0(instanceL2_n_11384));
  OAI21X1 instanceL2_g10741(.Y(instanceL2_n_11324), .A0(instanceL2_n_11392), .A1(
    instanceL2_n_11381), .B0(instanceL2_n_11378));
  AOI22X1 instanceL2_g10742(.Y(instanceL2_n_11862), .A0(instanceL2_n_11369), .A1(
    instanceL2_n_11365), .B0(instanceL2_n_11398), .B1(instanceL2_n_11394));
  INVX1 instanceL2_g10743(.Y(instanceL2_n_11867), .A(instanceL2_n_11866));
  NOR2BX1 instanceL2_g10744(.Y(\instanceL2_prod_terms[0][11][1] ), .AN(
    instanceL2_n_11366), .B(instanceL2_n_11361));
  NAND2XL instanceL2_g10745(.Y(instanceL2_n_11336), .A(instanceL2_n_11362), .B(
    instanceL2_n_11358));
  NAND2XL instanceL2_g10746(.Y(instanceL2_n_11338), .A(instanceL2_n_11367), .B(
    instanceL2_n_11359));
  NAND2BXL instanceL2_g10747(.Y(instanceL2_n_11340), .AN(instanceL2_n_11364), .B(
    instanceL2_n_11357));
  NAND2X1 instanceL2_g10748(.Y(instanceL2_n_11865), .A(instanceL2_n_11402), .B(
    instanceL2_n_11361));
  NAND2BX1 instanceL2_g10749(.Y(instanceL2_n_11866), .AN(instanceL2_n_11377), .B(
    instanceL2_n_11373));
  NAND2X1 instanceL2_g10750(.Y(instanceL2_n_11868), .A(instanceL2_n_11363), .B(
    instanceL2_n_11360));
  OAI22X1 instanceL2_g10751(.Y(instanceL2_n_11348), .A0(layer1_out[101]), .A1(
    layer1_out[102]), .B0(instanceL2_n_11402), .B1(instanceL2_n_11394));
  AO21XL instanceL2_g10752(.Y(instanceL2_n_11871), .A0(layer1_out[103]), .A1(
    layer1_out[102]), .B0(instanceL2_n_11379));
  OAI2BB1X1 instanceL2_g10753(.Y(instanceL2_n_11872), .A0N(instanceL2_n_11398),
     .A1N(instanceL2_n_11402), .B0(instanceL2_n_11356));
  OAI21X1 instanceL2_g10754(.Y(\instanceL2_prod_terms[2][11][2] ), .A0(
    layer1_out[99]), .A1(instanceL2_n_11402), .B0(instanceL2_n_11368));
  NOR2BX1 instanceL2_g10755(.Y(instanceL2_n_11869), .AN(instanceL2_n_11378), .B(
    instanceL2_n_11381));
  NAND2BX1 instanceL2_g10756(.Y(instanceL2_n_11346), .AN(instanceL2_n_11384), .B(
    instanceL2_n_11383));
  NAND2X1 instanceL2_g10757(.Y(instanceL2_n_11870), .A(instanceL2_n_11374), .B(
    instanceL2_n_11375));
  NAND2XL instanceL2_g10758(.Y(instanceL2_n_11369), .A(layer1_out[100]), .B(
    layer1_out[102]));
  NAND2XL instanceL2_g10759(.Y(instanceL2_n_11356), .A(layer1_out[101]), .B(
    layer1_out[100]));
  NAND2XL instanceL2_g10760(.Y(instanceL2_n_11357), .A(layer1_out[105]), .B(
    layer1_out[104]));
  NAND2X1 instanceL2_g10761(.Y(instanceL2_n_11358), .A(instanceL2_n_11390), .B(
    instanceL2_n_11400));
  NAND2X1 instanceL2_g10762(.Y(instanceL2_n_11359), .A(instanceL2_n_11392), .B(
    instanceL2_n_11388));
  NAND2X1 instanceL2_g10763(.Y(instanceL2_n_11360), .A(instanceL2_n_11388), .B(
    instanceL2_n_11400));
  NOR2X1 instanceL2_g10764(.Y(instanceL2_n_11361), .A(layer1_out[99]), .B(
    layer1_out[100]));
  NAND2X1 instanceL2_g10765(.Y(instanceL2_n_11362), .A(layer1_out[103]), .B(
    layer1_out[104]));
  NAND2X1 instanceL2_g10766(.Y(instanceL2_n_11363), .A(layer1_out[106]), .B(
    layer1_out[104]));
  NOR2X1 instanceL2_g10767(.Y(instanceL2_n_11364), .A(layer1_out[105]), .B(
    layer1_out[104]));
  NAND2X1 instanceL2_g10768(.Y(instanceL2_n_11365), .A(layer1_out[99]), .B(
    layer1_out[101]));
  NAND2XL instanceL2_g10769(.Y(instanceL2_n_11366), .A(layer1_out[100]), .B(
    layer1_out[99]));
  NAND2X1 instanceL2_g10770(.Y(instanceL2_n_11367), .A(layer1_out[105]), .B(
    layer1_out[106]));
  NAND2X1 instanceL2_g10771(.Y(instanceL2_n_11368), .A(instanceL2_n_11402), .B(
    layer1_out[99]));
  NAND2X1 instanceL2_g10772(.Y(instanceL2_n_11385), .A(instanceL2_n_11400), .B(
    instanceL2_n_11394));
  NAND2X1 instanceL2_g10773(.Y(instanceL2_n_11386), .A(instanceL2_n_11392), .B(
    layer1_out[103]));
  NAND2X1 instanceL2_g10774(.Y(instanceL2_n_11373), .A(layer1_out[105]), .B(
    layer1_out[103]));
  NAND2X1 instanceL2_g10775(.Y(instanceL2_n_11374), .A(layer1_out[104]), .B(
    instanceL2_n_11394));
  NAND2XL instanceL2_g10776(.Y(instanceL2_n_11375), .A(instanceL2_n_11400), .B(
    layer1_out[102]));
  NOR2X1 instanceL2_g10777(.Y(instanceL2_n_11376), .A(layer1_out[103]), .B(
    layer1_out[101]));
  NOR2XL instanceL2_g10778(.Y(instanceL2_n_11377), .A(layer1_out[105]), .B(
    layer1_out[103]));
  NAND2X1 instanceL2_g10779(.Y(instanceL2_n_11378), .A(instanceL2_n_11402), .B(
    layer1_out[103]));
  NOR2X1 instanceL2_g10780(.Y(instanceL2_n_11379), .A(layer1_out[103]), .B(
    layer1_out[102]));
  NOR2X1 instanceL2_g10781(.Y(instanceL2_n_11380), .A(instanceL2_n_11388), .B(
    layer1_out[104]));
  NOR2X1 instanceL2_g10782(.Y(instanceL2_n_11381), .A(layer1_out[103]), .B(
    instanceL2_n_11402));
  NOR2X1 instanceL2_g10783(.Y(instanceL2_n_11382), .A(instanceL2_n_11392), .B(
    layer1_out[103]));
  NAND2X1 instanceL2_g10784(.Y(instanceL2_n_11383), .A(instanceL2_n_11394), .B(
    layer1_out[100]));
  NOR2X1 instanceL2_g10785(.Y(instanceL2_n_11384), .A(layer1_out[100]), .B(
    instanceL2_n_11394));
  INVX1 instanceL2_g10786(.Y(instanceL2_n_11388), .A(layer1_out[106]));
  INVX1 instanceL2_g10787(.Y(instanceL2_n_11390), .A(layer1_out[103]));
  INVX1 instanceL2_g10788(.Y(instanceL2_n_11392), .A(layer1_out[105]));
  INVX1 instanceL2_g10789(.Y(instanceL2_n_11394), .A(layer1_out[102]));
  INVX1 instanceL2_g10790(.Y(instanceL2_n_11398), .A(layer1_out[100]));
  INVX1 instanceL2_g10791(.Y(instanceL2_n_11400), .A(layer1_out[104]));
  INVX1 instanceL2_g10792(.Y(instanceL2_n_11402), .A(layer1_out[101]));
  MXI2XL instanceL2_g10793(.Y(instanceL2_n_11403), .A(instanceL2_n_11394), .B(
    layer1_out[102]), .S0(instanceL2_n_11868));
  XNOR2X1 instanceL2_g10794(.Y(\instanceL2_prod_terms[4][12] [10]), .A(
    instanceL2_n_11893), .B(instanceL2_n_11143));
  AOI21X1 instanceL2_g10795(.Y(instanceL2_n_11143), .A0(instanceL2_n_11896), .A1(
    instanceL2_n_11146), .B0(instanceL2_n_11897));
  CLKXOR2X1 instanceL2_g10796(.Y(\instanceL2_prod_terms[4][12] [9]), .A(
    instanceL2_n_11895), .B(instanceL2_n_11146));
  ADDFX1 instanceL2_g10797(.CO(instanceL2_n_11146), .S(
    \instanceL2_prod_terms[4][12] [8]), .A(instanceL2_n_11900), .B(
    instanceL2_n_11890), .CI(instanceL2_n_11153));
  NAND2X1 instanceL2_g10798(.Y(\instanceL2_prod_terms[5][12] [9]), .A(
    instanceL2_n_11156), .B(instanceL2_n_11169));
  XOR2XL instanceL2_g10799(.Y(\instanceL2_prod_terms[5][12] [8]), .A(
    instanceL2_n_11234), .B(instanceL2_n_11873));
  OAI2BB1X1 instanceL2_g10800(.Y(\instanceL2_prod_terms[3][12] [9]), .A0N(
    layer1_out[115]), .A1N(instanceL2_n_11170), .B0(instanceL2_n_11156));
  ADDFX1 instanceL2_g10801(.CO(instanceL2_n_11153), .S(
    \instanceL2_prod_terms[4][12] [7]), .A(instanceL2_n_11219), .B(
    instanceL2_n_11889), .CI(instanceL2_n_11875));
  ADDFX1 instanceL2_g10802(.CO(instanceL2_n_11873), .S(
    \instanceL2_prod_terms[5][12] [7]), .A(instanceL2_n_11304), .B(
    instanceL2_n_11905), .CI(instanceL2_n_11874));
  OR2X1 instanceL2_g10803(.Y(instanceL2_n_11156), .A(layer1_out[115]), .B(
    instanceL2_n_11170));
  OAI2BB1X1 instanceL2_g10804(.Y(\instanceL2_prod_terms[7][12] [9]), .A0N(
    instanceL2_n_11927), .A1N(instanceL2_n_11876), .B0(instanceL2_n_11169));
  XNOR2X1 instanceL2_g10805(.Y(\instanceL2_prod_terms[3][12] [8]), .A(
    layer1_out[114]), .B(instanceL2_n_11877));
  ADDFX1 instanceL2_g10806(.CO(instanceL2_n_11874), .S(
    \instanceL2_prod_terms[5][12] [6]), .A(instanceL2_n_11923), .B(
    instanceL2_n_11907), .CI(instanceL2_n_11183));
  ADDFX1 instanceL2_g10807(.CO(instanceL2_n_11875), .S(
    \instanceL2_prod_terms[4][12] [6]), .A(instanceL2_n_11225), .B(
    instanceL2_n_11888), .CI(instanceL2_n_11878));
  NAND2X2 instanceL2_g10808(.Y(\instanceL2_prod_terms[3][12] [13]), .A(
    instanceL2_n_11913), .B(instanceL2_n_11877));
  OR2XL instanceL2_g10809(.Y(instanceL2_n_11169), .A(instanceL2_n_11927), .B(
    instanceL2_n_11876));
  NOR2BX1 instanceL2_g10810(.Y(instanceL2_n_11170), .AN(instanceL2_n_11877), .B(
    layer1_out[114]));
  OAI2BB1X1 instanceL2_g10811(.Y(instanceL2_n_11876), .A0N(layer1_out[114]),
     .A1N(instanceL2_n_11879), .B0(instanceL2_n_11177));
  INVX1 instanceL2_g10812(.Y(\instanceL2_prod_terms[7][12] [10]), .A(
    instanceL2_n_11177));
  OAI21X1 instanceL2_g10813(.Y(instanceL2_n_11177), .A0(layer1_out[114]), .A1(
    instanceL2_n_11879), .B0(layer1_out[115]));
  AOI21X1 instanceL2_g10814(.Y(\instanceL2_prod_terms[3][12] [7]), .A0(
    layer1_out[113]), .A1(instanceL2_n_11197), .B0(instanceL2_n_11877));
  XNOR2X1 instanceL2_g10815(.Y(\instanceL2_prod_terms[7][12] [8]), .A(
    instanceL2_n_11904), .B(instanceL2_n_11879));
  ADDFX1 instanceL2_g10816(.CO(instanceL2_n_11183), .S(
    \instanceL2_prod_terms[5][12] [5]), .A(instanceL2_n_11300), .B(
    instanceL2_n_11908), .CI(instanceL2_n_11882));
  ADDFX1 instanceL2_g10817(.CO(instanceL2_n_11878), .S(
    \instanceL2_prod_terms[4][12] [5]), .A(instanceL2_n_11914), .B(
    instanceL2_n_11891), .CI(instanceL2_n_11881));
  NOR2X1 instanceL2_g10818(.Y(instanceL2_n_11877), .A(layer1_out[113]), .B(
    instanceL2_n_11197));
  XNOR2X1 instanceL2_g10819(.Y(\instanceL2_prod_terms[7][12] [7]), .A(
    instanceL2_n_11899), .B(instanceL2_n_11880));
  OAI211X1 instanceL2_g10820(.Y(instanceL2_n_11879), .A0(instanceL2_n_11917),
     .A1(instanceL2_n_11883), .B0(instanceL2_n_11297), .C0(instanceL2_n_11916));
  NAND2X1 instanceL2_g10821(.Y(instanceL2_n_11880), .A(instanceL2_n_11297), .B(
    instanceL2_n_11883));
  OA21X1 instanceL2_g10822(.Y(\instanceL2_prod_terms[3][12] [6]), .A0(
    instanceL2_n_11929), .A1(instanceL2_n_11887), .B0(instanceL2_n_11197));
  XNOR2X1 instanceL2_g10823(.Y(\instanceL2_prod_terms[7][12] [6]), .A(
    instanceL2_n_11900), .B(instanceL2_n_11884));
  ADDFX1 instanceL2_g10824(.CO(instanceL2_n_11881), .S(
    \instanceL2_prod_terms[4][12] [4]), .A(layer1_out[112]), .B(
    instanceL2_n_11919), .CI(\instanceL2_prod_terms[3][12] [3]));
  ADDFX1 instanceL2_g10825(.CO(instanceL2_n_11882), .S(
    \instanceL2_prod_terms[5][12] [4]), .A(instanceL2_n_11302), .B(
    instanceL2_n_11906), .CI(instanceL2_n_11892));
  NAND2X1 instanceL2_g10826(.Y(instanceL2_n_11197), .A(instanceL2_n_11929), .B(
    instanceL2_n_11887));
  XNOR2X1 instanceL2_g10827(.Y(\instanceL2_prod_terms[7][12] [5]), .A(
    instanceL2_n_11902), .B(instanceL2_n_11885));
  NAND2X1 instanceL2_g10828(.Y(instanceL2_n_11883), .A(instanceL2_n_11912), .B(
    instanceL2_n_11884));
  OAI211X1 instanceL2_g10829(.Y(instanceL2_n_11884), .A0(instanceL2_n_11922),
     .A1(instanceL2_n_11886), .B0(instanceL2_n_11298), .C0(instanceL2_n_11921));
  XNOR2X1 instanceL2_g10830(.Y(\instanceL2_prod_terms[5][12] [3]), .A(
    instanceL2_n_11918), .B(instanceL2_n_11894));
  NAND2X1 instanceL2_g10831(.Y(instanceL2_n_11885), .A(instanceL2_n_11298), .B(
    instanceL2_n_11886));
  AOI21X1 instanceL2_g10832(.Y(\instanceL2_prod_terms[3][12] [5]), .A0(
    layer1_out[111]), .A1(instanceL2_n_11898), .B0(instanceL2_n_11887));
  XNOR2X1 instanceL2_g10833(.Y(\instanceL2_prod_terms[7][12] [4]), .A(
    instanceL2_n_11240), .B(instanceL2_n_11901));
  ADDFX1 instanceL2_g10834(.CO(instanceL2_n_11219), .S(instanceL2_n_11888), .A(
    layer1_out[114]), .B(instanceL2_n_11925), .CI(layer1_out[111]));
  ADDFX1 instanceL2_g10835(.CO(instanceL2_n_11890), .S(instanceL2_n_11889), .A(
    layer1_out[115]), .B(layer1_out[112]), .CI(instanceL2_n_11313));
  ADDFX1 instanceL2_g10836(.CO(instanceL2_n_11225), .S(instanceL2_n_11891), .A(
    layer1_out[113]), .B(layer1_out[110]), .CI(instanceL2_n_11926));
  NAND2X1 instanceL2_g10837(.Y(instanceL2_n_11886), .A(instanceL2_n_11920), .B(
    instanceL2_n_11240));
  AOI2BB1X1 instanceL2_g10838(.Y(instanceL2_n_11892), .A0N(layer1_out[110]),
     .A1N(instanceL2_n_11918), .B0(instanceL2_n_11903));
  NOR2X1 instanceL2_g10839(.Y(instanceL2_n_11887), .A(layer1_out[111]), .B(
    instanceL2_n_11898));
  XOR2XL instanceL2_g10840(.Y(\instanceL2_prod_terms[7][12] [3]), .A(
    instanceL2_n_11915), .B(instanceL2_n_11909));
  XNOR2X1 instanceL2_g10841(.Y(instanceL2_n_11893), .A(instanceL2_n_11301), .B(
    instanceL2_n_11904));
  AOI22X1 instanceL2_g10842(.Y(instanceL2_n_11234), .A0(layer1_out[115]), .A1(
    instanceL2_n_11917), .B0(layer1_out[114]), .B1(instanceL2_n_11299));
  MXI2XL instanceL2_g10843(.Y(instanceL2_n_11894), .A(instanceL2_n_11925), .B(
    layer1_out[110]), .S0(instanceL2_n_11903));
  NAND2X1 instanceL2_g10844(.Y(instanceL2_n_11240), .A(instanceL2_n_11915), .B(
    instanceL2_n_11910));
  NOR2BX1 instanceL2_g10845(.Y(instanceL2_n_11895), .AN(instanceL2_n_11896), .B(
    instanceL2_n_11897));
  OA21X1 instanceL2_g10846(.Y(\instanceL2_prod_terms[3][12] [4]), .A0(
    instanceL2_n_11925), .A1(instanceL2_n_11911), .B0(instanceL2_n_11898));
  AO21XL instanceL2_g10455(.Y(instanceL2_n_11896), .A0(layer1_out[113]), .A1(
    instanceL2_n_11929), .B0(instanceL2_n_11899));
  AOI21X1 instanceL2_g10456(.Y(\instanceL2_prod_terms[4][12] [3]), .A0(
    instanceL2_n_11307), .A1(instanceL2_n_11313), .B0(instanceL2_n_11919));
  AOI21X1 instanceL2_g10457(.Y(\instanceL2_prod_terms[5][12] [2]), .A0(
    layer1_out[108]), .A1(layer1_out[110]), .B0(instanceL2_n_11918));
  NAND2X1 instanceL2_g10458(.Y(instanceL2_n_11901), .A(instanceL2_n_11298), .B(
    instanceL2_n_11920));
  NOR2X1 instanceL2_g10459(.Y(instanceL2_n_11897), .A(layer1_out[112]), .B(
    instanceL2_n_11916));
  NAND2BXL instanceL2_g10460(.Y(instanceL2_n_11902), .AN(instanceL2_n_11922), .B(
    instanceL2_n_11921));
  NAND2X1 instanceL2_g10461(.Y(instanceL2_n_11898), .A(instanceL2_n_11925), .B(
    instanceL2_n_11911));
  NAND2BX1 instanceL2_g10462(.Y(instanceL2_n_11899), .AN(instanceL2_n_11917), .B(
    instanceL2_n_11916));
  NAND2X1 instanceL2_g10463(.Y(instanceL2_n_11900), .A(instanceL2_n_11297), .B(
    instanceL2_n_11912));
  OAI22X1 instanceL2_g10464(.Y(instanceL2_n_11905), .A0(layer1_out[115]), .A1(
    layer1_out[113]), .B0(instanceL2_n_11927), .B1(instanceL2_n_11928));
  OAI22X1 instanceL2_g10465(.Y(instanceL2_n_11906), .A0(layer1_out[112]), .A1(
    layer1_out[110]), .B0(instanceL2_n_11929), .B1(instanceL2_n_11925));
  OAI22X1 instanceL2_g10466(.Y(instanceL2_n_11907), .A0(layer1_out[114]), .A1(
    layer1_out[112]), .B0(instanceL2_n_11924), .B1(instanceL2_n_11929));
  OAI22X1 instanceL2_g10467(.Y(instanceL2_n_11908), .A0(layer1_out[113]), .A1(
    layer1_out[111]), .B0(instanceL2_n_11928), .B1(instanceL2_n_11313));
  OAI2BB1X1 instanceL2_g10468(.Y(instanceL2_n_11909), .A0N(instanceL2_n_11925),
     .A1N(instanceL2_n_11926), .B0(instanceL2_n_11910));
  AOI22X1 instanceL2_g10469(.Y(instanceL2_n_11903), .A0(instanceL2_n_11313), .A1(
    instanceL2_n_11926), .B0(layer1_out[109]), .B1(layer1_out[111]));
  AO21XL instanceL2_g10470(.Y(instanceL2_n_11904), .A0(layer1_out[115]), .A1(
    layer1_out[114]), .B0(instanceL2_n_11913));
  OAI2BB1X1 instanceL2_g10471(.Y(\instanceL2_prod_terms[3][12] [3]), .A0N(
    layer1_out[109]), .A1N(instanceL2_n_11307), .B0(instanceL2_n_11914));
  NAND2XL instanceL2_g10472(.Y(instanceL2_n_11910), .A(layer1_out[110]), .B(
    layer1_out[109]));
  NOR2X1 instanceL2_g10473(.Y(instanceL2_n_11911), .A(layer1_out[108]), .B(
    layer1_out[109]));
  NAND2X1 instanceL2_g10474(.Y(instanceL2_n_11912), .A(instanceL2_n_11928), .B(
    instanceL2_n_11929));
  NOR2X1 instanceL2_g10475(.Y(instanceL2_n_11913), .A(layer1_out[114]), .B(
    layer1_out[115]));
  NAND2X1 instanceL2_g10476(.Y(instanceL2_n_11914), .A(instanceL2_n_11926), .B(
    layer1_out[108]));
  NAND2XL instanceL2_g10477(.Y(instanceL2_n_11915), .A(layer1_out[108]), .B(
    layer1_out[109]));
  NAND2XL instanceL2_g10478(.Y(instanceL2_n_11916), .A(layer1_out[114]), .B(
    layer1_out[113]));
  NOR2X1 instanceL2_g10479(.Y(instanceL2_n_11917), .A(layer1_out[113]), .B(
    layer1_out[114]));
  NOR2X1 instanceL2_g10480(.Y(instanceL2_n_11918), .A(layer1_out[108]), .B(
    layer1_out[110]));
  NOR2X1 instanceL2_g10481(.Y(instanceL2_n_11919), .A(instanceL2_n_11313), .B(
    instanceL2_n_11307));
  NAND2XL instanceL2_g10482(.Y(instanceL2_n_11299), .A(layer1_out[115]), .B(
    instanceL2_n_11928));
  NAND2X1 instanceL2_g10483(.Y(instanceL2_n_11920), .A(instanceL2_n_11925), .B(
    instanceL2_n_11313));
  NOR2X1 instanceL2_g10484(.Y(instanceL2_n_11300), .A(layer1_out[110]), .B(
    instanceL2_n_11929));
  NAND2XL instanceL2_g10485(.Y(instanceL2_n_11921), .A(layer1_out[112]), .B(
    layer1_out[111]));
  NOR2XL instanceL2_g10486(.Y(instanceL2_n_11922), .A(layer1_out[112]), .B(
    layer1_out[111]));
  NAND2XL instanceL2_g10487(.Y(instanceL2_n_11301), .A(instanceL2_n_11928), .B(
    layer1_out[114]));
  NOR2X1 instanceL2_g10847(.Y(instanceL2_n_11302), .A(layer1_out[109]), .B(
    instanceL2_n_11313));
  NOR2X1 instanceL2_g10848(.Y(instanceL2_n_11923), .A(instanceL2_n_11928), .B(
    layer1_out[111]));
  NOR2X1 instanceL2_g10849(.Y(instanceL2_n_11304), .A(instanceL2_n_11924), .B(
    layer1_out[112]));
  NAND2X1 instanceL2_g10850(.Y(instanceL2_n_11297), .A(layer1_out[112]), .B(
    layer1_out[113]));
  NAND2X1 instanceL2_g10851(.Y(instanceL2_n_11298), .A(layer1_out[111]), .B(
    layer1_out[110]));
  INVX1 instanceL2_g10852(.Y(instanceL2_n_11307), .A(layer1_out[108]));
  INVX1 instanceL2_g10853(.Y(instanceL2_n_11924), .A(layer1_out[114]));
  INVX1 instanceL2_g10854(.Y(instanceL2_n_11925), .A(layer1_out[110]));
  INVX1 instanceL2_g10855(.Y(instanceL2_n_11313), .A(layer1_out[111]));
  INVX1 instanceL2_g10856(.Y(instanceL2_n_11926), .A(layer1_out[109]));
  INVX1 instanceL2_g10857(.Y(instanceL2_n_11927), .A(layer1_out[115]));
  INVX1 instanceL2_g10858(.Y(instanceL2_n_11928), .A(layer1_out[113]));
  INVX1 instanceL2_g10859(.Y(instanceL2_n_11929), .A(layer1_out[112]));
  XNOR2X1 instanceL2_g10860(.Y(\instanceL2_prod_terms[2][6] [11]), .A(
    instanceL2_n_11935), .B(instanceL2_n_11039));
  ADDFX1 instanceL2_g10861(.CO(instanceL2_n_11039), .S(
    \instanceL2_prod_terms[2][6] [10]), .A(instanceL2_n_11949), .B(
    instanceL2_n_11941), .CI(instanceL2_n_11041));
  ADDFX1 instanceL2_g10862(.CO(instanceL2_n_11041), .S(
    \instanceL2_prod_terms[2][6] [9]), .A(instanceL2_n_11123), .B(
    instanceL2_n_11115), .CI(instanceL2_n_11045));
  OA21X1 instanceL2_g10863(.Y(\instanceL2_prod_terms[3][6] [10]), .A0(
    instanceL2_n_11969), .A1(instanceL2_n_11055), .B0(
    \instanceL2_prod_terms[2][6] [13]));
  ADDFX1 instanceL2_g10864(.CO(instanceL2_n_11045), .S(
    \instanceL2_prod_terms[2][6] [8]), .A(instanceL2_n_11942), .B(
    instanceL2_n_11936), .CI(instanceL2_n_11057));
  NAND2X1 instanceL2_g10865(.Y(\instanceL2_prod_terms[2][6] [13]), .A(
    instanceL2_n_11969), .B(instanceL2_n_11055));
  MXI2XL instanceL2_g10866(.Y(\instanceL2_prod_terms[4][6] [10]), .A(
    layer1_out[62]), .B(instanceL2_n_11969), .S0(instanceL2_n_11059));
  AOI21X1 instanceL2_g10867(.Y(\instanceL2_prod_terms[3][6] [9]), .A0(
    layer1_out[61]), .A1(instanceL2_n_11071), .B0(instanceL2_n_11055));
  OAI21X1 instanceL2_g10868(.Y(\instanceL2_prod_terms[4][6] [11]), .A0(
    instanceL2_n_11969), .A1(instanceL2_n_11064), .B0(instanceL2_n_11139));
  MX2XL instanceL2_g10869(.Y(\instanceL2_prod_terms[4][6] [9]), .A(
    layer1_out[61]), .B(instanceL2_n_11966), .S0(instanceL2_n_11063));
  ADDFX1 instanceL2_g10870(.CO(instanceL2_n_11057), .S(
    \instanceL2_prod_terms[2][6] [7]), .A(instanceL2_n_11940), .B(
    instanceL2_n_11937), .CI(instanceL2_n_11930));
  NOR2X1 instanceL2_g10871(.Y(instanceL2_n_11055), .A(layer1_out[61]), .B(
    instanceL2_n_11071));
  AND2XL instanceL2_g10872(.Y(instanceL2_n_11059), .A(instanceL2_n_11139), .B(
    instanceL2_n_11064));
  NAND2X1 instanceL2_g10873(.Y(instanceL2_n_11063), .A(instanceL2_n_11957), .B(
    instanceL2_n_11068));
  XNOR2X1 instanceL2_g10874(.Y(\instanceL2_prod_terms[4][6] [8]), .A(
    instanceL2_n_11943), .B(instanceL2_n_11076));
  OR2XL instanceL2_g10875(.Y(instanceL2_n_11064), .A(instanceL2_n_11966), .B(
    instanceL2_n_11068));
  NAND2BX1 instanceL2_g10876(.Y(instanceL2_n_11068), .AN(instanceL2_n_11959), .B(
    instanceL2_n_11076));
  OA21X1 instanceL2_g10877(.Y(\instanceL2_prod_terms[3][6] [8]), .A0(
    instanceL2_n_11965), .A1(instanceL2_n_11932), .B0(instanceL2_n_11071));
  ADDFX1 instanceL2_g10878(.CO(instanceL2_n_11930), .S(
    \instanceL2_prod_terms[2][6] [6]), .A(instanceL2_n_11939), .B(
    instanceL2_n_11938), .CI(instanceL2_n_11085));
  NAND2X1 instanceL2_g10879(.Y(instanceL2_n_11071), .A(instanceL2_n_11965), .B(
    instanceL2_n_11932));
  XNOR2X1 instanceL2_g10880(.Y(\instanceL2_prod_terms[4][6] [7]), .A(
    instanceL2_n_11946), .B(instanceL2_n_11931));
  OAI2BB1X1 instanceL2_g10881(.Y(instanceL2_n_11076), .A0N(instanceL2_n_11961),
     .A1N(instanceL2_n_11931), .B0(instanceL2_n_11960));
  OAI21X1 instanceL2_g10882(.Y(instanceL2_n_11931), .A0(instanceL2_n_11955), .A1(
    instanceL2_n_11090), .B0(instanceL2_n_11954));
  AOI21X1 instanceL2_g10883(.Y(\instanceL2_prod_terms[3][6] [7]), .A0(
    layer1_out[59]), .A1(instanceL2_n_11094), .B0(instanceL2_n_11932));
  XNOR2X1 instanceL2_g10884(.Y(\instanceL2_prod_terms[4][6] [6]), .A(
    instanceL2_n_11944), .B(instanceL2_n_11090));
  ADDFX1 instanceL2_g10885(.CO(instanceL2_n_11085), .S(
    \instanceL2_prod_terms[2][6] [5]), .A(instanceL2_n_11953), .B(
    instanceL2_n_11119), .CI(instanceL2_n_11933));
  NOR2X1 instanceL2_g10886(.Y(instanceL2_n_11932), .A(layer1_out[59]), .B(
    instanceL2_n_11094));
  AOI21X1 instanceL2_g10887(.Y(instanceL2_n_11090), .A0(instanceL2_n_11962), .A1(
    instanceL2_n_11100), .B0(instanceL2_n_11964));
  XNOR2X1 instanceL2_g10888(.Y(\instanceL2_prod_terms[4][6] [5]), .A(
    instanceL2_n_11947), .B(instanceL2_n_11100));
  OA21X1 instanceL2_g10889(.Y(\instanceL2_prod_terms[3][6] [6]), .A0(
    instanceL2_n_11971), .A1(instanceL2_n_11934), .B0(instanceL2_n_11094));
  ADDFX1 instanceL2_g10890(.CO(instanceL2_n_11933), .S(
    \instanceL2_prod_terms[2][6] [4]), .A(layer1_out[57]), .B(
    instanceL2_n_11120), .CI(\instanceL2_prod_terms[3][6] [3]));
  NAND2X1 instanceL2_g10891(.Y(instanceL2_n_11094), .A(instanceL2_n_11971), .B(
    instanceL2_n_11934));
  XNOR2X1 instanceL2_g10892(.Y(\instanceL2_prod_terms[4][6] [4]), .A(
    instanceL2_n_11945), .B(instanceL2_n_11105));
  OAI21X1 instanceL2_g10893(.Y(instanceL2_n_11100), .A0(instanceL2_n_11180), .A1(
    instanceL2_n_11105), .B0(instanceL2_n_11956));
  INVX1 instanceL2_g10894(.Y(\instanceL2_prod_terms[4][6] [3]), .A(
    instanceL2_n_11106));
  ADDFX1 instanceL2_g10895(.CO(instanceL2_n_11105), .S(instanceL2_n_11106), .A(
    instanceL2_n_11968), .B(instanceL2_n_11967), .CI(instanceL2_n_11172));
  AOI21X1 instanceL2_g10896(.Y(\instanceL2_prod_terms[3][6] [5]), .A0(
    layer1_out[57]), .A1(instanceL2_n_11140), .B0(instanceL2_n_11934));
  NOR2X1 instanceL2_g10897(.Y(instanceL2_n_11934), .A(layer1_out[57]), .B(
    instanceL2_n_11140));
  XNOR2X1 instanceL2_g10898(.Y(instanceL2_n_11935), .A(instanceL2_n_11958), .B(
    instanceL2_n_11948));
  XNOR2X1 instanceL2_g10899(.Y(instanceL2_n_11936), .A(layer1_out[59]), .B(
    instanceL2_n_11951));
  MXI2XL instanceL2_g10900(.Y(instanceL2_n_11937), .A(instanceL2_n_11971), .B(
    layer1_out[58]), .S0(instanceL2_n_11163));
  MXI2XL instanceL2_g10901(.Y(instanceL2_n_11115), .A(instanceL2_n_11969), .B(
    layer1_out[62]), .S0(instanceL2_n_11160));
  MXI2XL instanceL2_g10902(.Y(instanceL2_n_11938), .A(instanceL2_n_11967), .B(
    layer1_out[57]), .S0(instanceL2_n_11950));
  XNOR2X1 instanceL2_g10903(.Y(instanceL2_n_11119), .A(layer1_out[56]), .B(
    instanceL2_n_11154));
  INVX1 instanceL2_g10904(.Y(instanceL2_n_11120), .A(instanceL2_n_11172));
  OAI2BB1X1 instanceL2_g10905(.Y(instanceL2_n_11123), .A0N(instanceL2_n_11971),
     .A1N(instanceL2_n_11961), .B0(instanceL2_n_11960));
  OAI21X1 instanceL2_g10906(.Y(instanceL2_n_11939), .A0(layer1_out[55]), .A1(
    instanceL2_n_11180), .B0(instanceL2_n_11956));
  OAI2BB1X1 instanceL2_g10907(.Y(instanceL2_n_11940), .A0N(instanceL2_n_11970),
     .A1N(instanceL2_n_11962), .B0(instanceL2_n_11963));
  OA21X1 instanceL2_g10908(.Y(\instanceL2_prod_terms[3][6] [4]), .A0(
    instanceL2_n_11970), .A1(instanceL2_n_11952), .B0(instanceL2_n_11140));
  OAI21X1 instanceL2_g10909(.Y(instanceL2_n_11941), .A0(layer1_out[59]), .A1(
    instanceL2_n_11959), .B0(instanceL2_n_11957));
  OAI21X1 instanceL2_g10910(.Y(instanceL2_n_11942), .A0(layer1_out[57]), .A1(
    instanceL2_n_11955), .B0(instanceL2_n_11954));
  OA21X1 instanceL2_g10911(.Y(\instanceL2_prod_terms[2][6] [3]), .A0(
    layer1_out[56]), .A1(layer1_out[54]), .B0(instanceL2_n_11172));
  NAND2BX1 instanceL2_g10912(.Y(instanceL2_n_11943), .AN(instanceL2_n_11959), .B(
    instanceL2_n_11957));
  OR2XL instanceL2_g10913(.Y(instanceL2_n_11139), .A(instanceL2_n_11966), .B(
    instanceL2_n_11957));
  NOR2BX1 instanceL2_g10914(.Y(instanceL2_n_11944), .AN(instanceL2_n_11954), .B(
    instanceL2_n_11955));
  NOR2BX1 instanceL2_g10915(.Y(instanceL2_n_11945), .AN(instanceL2_n_11956), .B(
    instanceL2_n_11180));
  NAND2XL instanceL2_g10916(.Y(instanceL2_n_11946), .A(instanceL2_n_11960), .B(
    instanceL2_n_11961));
  NAND2XL instanceL2_g10917(.Y(instanceL2_n_11947), .A(instanceL2_n_11963), .B(
    instanceL2_n_11962));
  NAND2X1 instanceL2_g10918(.Y(instanceL2_n_11140), .A(instanceL2_n_11970), .B(
    instanceL2_n_11952));
  OAI22X1 instanceL2_g10919(.Y(instanceL2_n_11948), .A0(layer1_out[62]), .A1(
    layer1_out[61]), .B0(instanceL2_n_11969), .B1(instanceL2_n_11966));
  AOI21X1 instanceL2_g10920(.Y(instanceL2_n_11949), .A0(instanceL2_n_11966), .A1(
    layer1_out[60]), .B0(instanceL2_n_11958));
  AOI22X1 instanceL2_g10921(.Y(instanceL2_n_11154), .A0(instanceL2_n_11971), .A1(
    instanceL2_n_11968), .B0(layer1_out[58]), .B1(layer1_out[55]));
  OAI22X1 instanceL2_g10922(.Y(instanceL2_n_11950), .A0(layer1_out[59]), .A1(
    layer1_out[56]), .B0(instanceL2_n_11972), .B1(instanceL2_n_11970));
  AOI22X1 instanceL2_g10923(.Y(instanceL2_n_11951), .A0(instanceL2_n_11966), .A1(
    instanceL2_n_11971), .B0(layer1_out[61]), .B1(layer1_out[58]));
  OAI22X1 instanceL2_g10924(.Y(instanceL2_n_11160), .A0(layer1_out[60]), .A1(
    layer1_out[59]), .B0(instanceL2_n_11965), .B1(instanceL2_n_11972));
  OAI22X1 instanceL2_g10925(.Y(instanceL2_n_11163), .A0(layer1_out[60]), .A1(
    layer1_out[57]), .B0(instanceL2_n_11965), .B1(instanceL2_n_11967));
  OAI21X1 instanceL2_g10926(.Y(\instanceL2_prod_terms[3][6] [3]), .A0(
    instanceL2_n_11968), .A1(layer1_out[54]), .B0(instanceL2_n_11953));
  NOR2XL instanceL2_g10927(.Y(instanceL2_n_11952), .A(layer1_out[55]), .B(
    layer1_out[54]));
  NAND2X1 instanceL2_g10928(.Y(instanceL2_n_11953), .A(instanceL2_n_11968), .B(
    layer1_out[54]));
  NAND2X1 instanceL2_g10929(.Y(instanceL2_n_11954), .A(layer1_out[58]), .B(
    layer1_out[60]));
  NOR2X1 instanceL2_g10930(.Y(instanceL2_n_11955), .A(layer1_out[60]), .B(
    layer1_out[58]));
  NAND2X1 instanceL2_g10931(.Y(instanceL2_n_11956), .A(layer1_out[56]), .B(
    layer1_out[58]));
  NAND2X1 instanceL2_g10932(.Y(instanceL2_n_11957), .A(layer1_out[62]), .B(
    layer1_out[60]));
  NAND2X1 instanceL2_g10933(.Y(instanceL2_n_11172), .A(layer1_out[54]), .B(
    layer1_out[56]));
  INVX1 instanceL2_g10934(.Y(instanceL2_n_11964), .A(instanceL2_n_11963));
  NOR2X1 instanceL2_g10935(.Y(instanceL2_n_11958), .A(instanceL2_n_11966), .B(
    layer1_out[60]));
  NOR2X1 instanceL2_g10936(.Y(instanceL2_n_11959), .A(layer1_out[62]), .B(
    layer1_out[60]));
  NAND2X1 instanceL2_g10264(.Y(instanceL2_n_11960), .A(layer1_out[61]), .B(
    layer1_out[59]));
  NAND2X1 instanceL2_g10265(.Y(instanceL2_n_11961), .A(instanceL2_n_11966), .B(
    instanceL2_n_11972));
  NAND2X1 instanceL2_g10266(.Y(instanceL2_n_11962), .A(instanceL2_n_11972), .B(
    instanceL2_n_11967));
  NAND2X1 instanceL2_g10267(.Y(instanceL2_n_11963), .A(layer1_out[59]), .B(
    layer1_out[57]));
  NOR2X1 instanceL2_g10268(.Y(instanceL2_n_11180), .A(layer1_out[58]), .B(
    layer1_out[56]));
  INVX1 instanceL2_g10269(.Y(instanceL2_n_11965), .A(layer1_out[60]));
  INVX1 instanceL2_g10270(.Y(instanceL2_n_11966), .A(layer1_out[61]));
  INVX1 instanceL2_g10271(.Y(instanceL2_n_11967), .A(layer1_out[57]));
  INVX1 instanceL2_g10272(.Y(instanceL2_n_11968), .A(layer1_out[55]));
  INVX1 instanceL2_g10273(.Y(instanceL2_n_11969), .A(layer1_out[62]));
  INVX1 instanceL2_g10274(.Y(instanceL2_n_11970), .A(layer1_out[56]));
  INVX1 instanceL2_g10275(.Y(instanceL2_n_11971), .A(layer1_out[58]));
  INVX1 instanceL2_g10276(.Y(instanceL2_n_11972), .A(layer1_out[59]));
  INVX1 instanceL2_g10013(.Y(\instanceL2_prod_terms[8][19] [11]), .A(
    instanceL2_n_11973));
  AOI31X1 instanceL2_g10014(.Y(instanceL2_n_11973), .A0(instanceL2_n_11107), .A1(
    layer1_out[178]), .A2(instanceL2_n_11974), .B0(instanceL2_n_11013));
  MX2XL instanceL2_g10015(.Y(\instanceL2_prod_terms[8][19] [10]), .A(
    instanceL2_n_11107), .B(layer1_out[177]), .S0(instanceL2_n_11974));
  ADDFX1 instanceL2_g10016(.CO(instanceL2_n_11974), .S(
    \instanceL2_prod_terms[8][19] [9]), .A(instanceL2_n_11988), .B(
    instanceL2_n_11979), .CI(instanceL2_n_10989));
  ADDFX1 instanceL2_g10017(.CO(instanceL2_n_10989), .S(
    \instanceL2_prod_terms[8][19] [8]), .A(instanceL2_n_11981), .B(
    instanceL2_n_11067), .CI(instanceL2_n_10993));
  OAI2BB1X1 instanceL2_g10018(.Y(\instanceL2_prod_terms[5][19] [9]), .A0N(
    layer1_out[177]), .A1N(instanceL2_n_11000), .B0(instanceL2_n_11002));
  ADDFX1 instanceL2_g10019(.CO(instanceL2_n_10993), .S(
    \instanceL2_prod_terms[8][19] [7]), .A(instanceL2_n_11070), .B(
    instanceL2_n_11060), .CI(instanceL2_n_11008));
  AND2XL instanceL2_g10020(.Y(\instanceL2_prod_terms[5][19] [10]), .A(
    layer1_out[178]), .B(instanceL2_n_11002));
  OAI21X1 instanceL2_g10021(.Y(\instanceL2_prod_terms[5][19] [8]), .A0(
    instanceL2_n_11988), .A1(instanceL2_n_11003), .B0(instanceL2_n_11000));
  NAND2X1 instanceL2_g10022(.Y(instanceL2_n_11000), .A(instanceL2_n_11988), .B(
    instanceL2_n_11003));
  NAND2X1 instanceL2_g10023(.Y(instanceL2_n_11002), .A(instanceL2_n_11089), .B(
    instanceL2_n_11003));
  AOI22X1 instanceL2_g10024(.Y(instanceL2_n_11003), .A0(instanceL2_n_11092), .A1(
    instanceL2_n_11011), .B0(instanceL2_n_11103), .B1(layer1_out[175]));
  XOR2XL instanceL2_g10025(.Y(\instanceL2_prod_terms[5][19] [7]), .A(
    instanceL2_n_11981), .B(instanceL2_n_11011));
  ADDFX1 instanceL2_g10026(.CO(instanceL2_n_11008), .S(
    \instanceL2_prod_terms[8][19] [6]), .A(instanceL2_n_11052), .B(
    instanceL2_n_11978), .CI(instanceL2_n_11017));
  AO21X1 instanceL2_g10027(.Y(\instanceL2_prod_terms[1][19] [9]), .A0(
    layer1_out[178]), .A1(instanceL2_n_11023), .B0(instanceL2_n_11013));
  ADDFX1 instanceL2_g10028(.CO(instanceL2_n_11011), .S(
    \instanceL2_prod_terms[5][19] [6]), .A(instanceL2_n_11107), .B(
    layer1_out[174]), .CI(instanceL2_n_11020));
  NOR2X1 instanceL2_g10029(.Y(instanceL2_n_11013), .A(layer1_out[178]), .B(
    instanceL2_n_11023));
  ADDFX1 instanceL2_g10030(.CO(instanceL2_n_11017), .S(
    \instanceL2_prod_terms[8][19] [5]), .A(instanceL2_n_11985), .B(
    instanceL2_n_11051), .CI(instanceL2_n_11026));
  XNOR2X1 instanceL2_g10031(.Y(\instanceL2_prod_terms[1][19] [8]), .A(
    layer1_out[177]), .B(instanceL2_n_11031));
  ADDFX1 instanceL2_g10032(.CO(instanceL2_n_11020), .S(
    \instanceL2_prod_terms[5][19] [5]), .A(instanceL2_n_11988), .B(
    layer1_out[173]), .CI(instanceL2_n_11030));
  NAND2X1 instanceL2_g10033(.Y(\instanceL2_prod_terms[1][19] [13]), .A(
    instanceL2_n_11986), .B(instanceL2_n_11031));
  AND2XL instanceL2_g10034(.Y(instanceL2_n_11023), .A(instanceL2_n_11107), .B(
    instanceL2_n_11031));
  ADDFX1 instanceL2_g10035(.CO(instanceL2_n_11026), .S(
    \instanceL2_prod_terms[8][19] [4]), .A(layer1_out[175]), .B(
    instanceL2_n_11072), .CI(instanceL2_n_11038));
  AOI21X1 instanceL2_g10036(.Y(\instanceL2_prod_terms[1][19] [7]), .A0(
    layer1_out[176]), .A1(instanceL2_n_11975), .B0(instanceL2_n_11031));
  ADDFX1 instanceL2_g10037(.CO(instanceL2_n_11030), .S(
    \instanceL2_prod_terms[5][19] [4]), .A(layer1_out[172]), .B(
    instanceL2_n_11099), .CI(instanceL2_n_11042));
  NOR2X1 instanceL2_g10038(.Y(instanceL2_n_11031), .A(layer1_out[176]), .B(
    instanceL2_n_11975));
  OAI21X1 instanceL2_g10039(.Y(\instanceL2_prod_terms[1][19] [5]), .A0(
    layer1_out[174]), .A1(instanceL2_n_11976), .B0(instanceL2_n_11050));
  ADDFX1 instanceL2_g10040(.CO(instanceL2_n_11038), .S(
    \instanceL2_prod_terms[8][19] [3]), .A(layer1_out[174]), .B(layer1_out[173]),
     .CI(instanceL2_n_11977));
  OA21X1 instanceL2_g10041(.Y(\instanceL2_prod_terms[1][19] [6]), .A0(
    instanceL2_n_11099), .A1(instanceL2_n_11053), .B0(instanceL2_n_11975));
  NAND2BXL instanceL2_g10042(.Y(instanceL2_n_11042), .AN(instanceL2_n_11053), .B(
    instanceL2_n_11985));
  OAI21X1 instanceL2_g10043(.Y(\instanceL2_prod_terms[5][19] [3]), .A0(
    instanceL2_n_11976), .A1(instanceL2_n_11072), .B0(instanceL2_n_11050));
  NAND2X1 instanceL2_g10044(.Y(instanceL2_n_11975), .A(instanceL2_n_11099), .B(
    instanceL2_n_11053));
  ADDFX1 instanceL2_g10045(.CO(instanceL2_n_11052), .S(instanceL2_n_11051), .A(
    instanceL2_n_11095), .B(layer1_out[175]), .CI(layer1_out[176]));
  NAND2X1 instanceL2_g10046(.Y(instanceL2_n_11050), .A(instanceL2_n_11976), .B(
    instanceL2_n_11072));
  XOR2XL instanceL2_g10047(.Y(\instanceL2_prod_terms[8][19] [2]), .A(
    instanceL2_n_11984), .B(instanceL2_n_11982));
  NOR2X1 instanceL2_g10048(.Y(instanceL2_n_11053), .A(layer1_out[174]), .B(
    instanceL2_n_11980));
  INVX1 instanceL2_g10049(.Y(instanceL2_n_11976), .A(instanceL2_n_11980));
  NAND2XL instanceL2_g10050(.Y(instanceL2_n_11977), .A(instanceL2_n_11984), .B(
    instanceL2_n_11987));
  MX2XL instanceL2_g10051(.Y(instanceL2_n_11978), .A(layer1_out[176]), .B(
    instanceL2_n_11988), .S0(instanceL2_n_11983));
  XNOR2X1 instanceL2_g10052(.Y(instanceL2_n_11060), .A(instanceL2_n_11107), .B(
    instanceL2_n_11078));
  INVX1 instanceL2_g10053(.Y(instanceL2_n_11979), .A(instanceL2_n_11092));
  OA21X1 instanceL2_g10054(.Y(\instanceL2_prod_terms[1][19] [4]), .A0(
    instanceL2_n_11097), .A1(instanceL2_n_11084), .B0(instanceL2_n_11980));
  OAI22X1 instanceL2_g10055(.Y(instanceL2_n_11067), .A0(layer1_out[174]), .A1(
    instanceL2_n_11986), .B0(instanceL2_n_11103), .B1(instanceL2_n_11107));
  OAI22X1 instanceL2_g10056(.Y(instanceL2_n_11070), .A0(layer1_out[173]), .A1(
    instanceL2_n_11089), .B0(instanceL2_n_11107), .B1(instanceL2_n_11988));
  NOR2BX1 instanceL2_g10057(.Y(\instanceL2_prod_terms[1][19] [3]), .AN(
    instanceL2_n_11984), .B(instanceL2_n_11084));
  OAI21X1 instanceL2_g10058(.Y(instanceL2_n_11072), .A0(layer1_out[171]), .A1(
    instanceL2_n_11101), .B0(instanceL2_n_11985));
  NAND2X1 instanceL2_g10059(.Y(instanceL2_n_11980), .A(instanceL2_n_11097), .B(
    instanceL2_n_11084));
  OAI22X1 instanceL2_g10060(.Y(instanceL2_n_11078), .A0(layer1_out[178]), .A1(
    layer1_out[174]), .B0(instanceL2_n_11103), .B1(instanceL2_n_11101));
  OAI2BB1X1 instanceL2_g10061(.Y(instanceL2_n_11982), .A0N(instanceL2_n_11095),
     .A1N(instanceL2_n_11097), .B0(instanceL2_n_11987));
  OAI22X1 instanceL2_g10062(.Y(instanceL2_n_11983), .A0(layer1_out[177]), .A1(
    layer1_out[173]), .B0(instanceL2_n_11107), .B1(instanceL2_n_11097));
  OAI22X1 instanceL2_g10063(.Y(instanceL2_n_11981), .A0(layer1_out[178]), .A1(
    layer1_out[175]), .B0(instanceL2_n_11103), .B1(instanceL2_n_11099));
  NOR2X1 instanceL2_g10064(.Y(instanceL2_n_11084), .A(layer1_out[172]), .B(
    layer1_out[171]));
  NAND2XL instanceL2_g10065(.Y(instanceL2_n_11984), .A(layer1_out[172]), .B(
    layer1_out[171]));
  NAND2X1 instanceL2_g10066(.Y(instanceL2_n_11985), .A(layer1_out[171]), .B(
    instanceL2_n_11101));
  NOR2X1 instanceL2_g10067(.Y(instanceL2_n_11089), .A(layer1_out[177]), .B(
    layer1_out[176]));
  NOR2XL instanceL2_g10068(.Y(instanceL2_n_11986), .A(layer1_out[178]), .B(
    layer1_out[177]));
  NAND2XL instanceL2_g10069(.Y(instanceL2_n_11987), .A(layer1_out[172]), .B(
    layer1_out[173]));
  NAND2X1 instanceL2_g10070(.Y(instanceL2_n_11092), .A(instanceL2_n_11099), .B(
    layer1_out[178]));
  INVX1 instanceL2_g10071(.Y(instanceL2_n_11095), .A(layer1_out[172]));
  INVX1 instanceL2_g10072(.Y(instanceL2_n_11097), .A(layer1_out[173]));
  INVX1 instanceL2_g10073(.Y(instanceL2_n_11099), .A(layer1_out[175]));
  INVX1 instanceL2_g10074(.Y(instanceL2_n_11101), .A(layer1_out[174]));
  INVX1 instanceL2_g10075(.Y(instanceL2_n_11103), .A(layer1_out[178]));
  INVX1 instanceL2_g10076(.Y(instanceL2_n_11988), .A(layer1_out[176]));
  INVX1 instanceL2_g10077(.Y(instanceL2_n_11107), .A(layer1_out[177]));
  MX2XL instanceL2_g10937(.Y(\instanceL2_prod_terms[6][15] [11]), .A(
    layer1_out[142]), .B(instanceL2_n_11411), .S0(instanceL2_n_11989));
  OA21X1 instanceL2_g10938(.Y(\instanceL2_prod_terms[6][15] [10]), .A0(
    instanceL2_n_11404), .A1(instanceL2_n_11991), .B0(instanceL2_n_11989));
  XNOR2X1 instanceL2_g10939(.Y(\instanceL2_prod_terms[6][15] [9]), .A(
    instanceL2_n_12022), .B(instanceL2_n_11990));
  NAND2X1 instanceL2_g10940(.Y(instanceL2_n_11989), .A(instanceL2_n_11404), .B(
    instanceL2_n_11991));
  NAND2BX1 instanceL2_g10941(.Y(\instanceL2_prod_terms[6][15] [13]), .AN(
    instanceL2_n_11992), .B(instanceL2_n_12054));
  OAI2BB1X1 instanceL2_g10942(.Y(instanceL2_n_11990), .A0N(instanceL2_n_12015),
     .A1N(instanceL2_n_11993), .B0(instanceL2_n_12016));
  XNOR2X1 instanceL2_g10943(.Y(\instanceL2_prod_terms[6][15] [8]), .A(
    instanceL2_n_12014), .B(instanceL2_n_11993));
  OAI211X1 instanceL2_g10944(.Y(instanceL2_n_11991), .A0(instanceL2_n_12034),
     .A1(instanceL2_n_12016), .B0(instanceL2_n_12033), .C0(instanceL2_n_11992));
  NAND3BXL instanceL2_g10945(.Y(instanceL2_n_11992), .AN(instanceL2_n_12034), .B(
    instanceL2_n_12015), .C(instanceL2_n_11993));
  ADDFX1 instanceL2_g10946(.CO(instanceL2_n_11993), .S(
    \instanceL2_prod_terms[6][15] [7]), .A(instanceL2_n_12025), .B(
    instanceL2_n_12019), .CI(instanceL2_n_11994));
  OAI211X1 instanceL2_g10947(.Y(\instanceL2_prod_terms[1][15] [9]), .A0(
    instanceL2_n_11404), .A1(instanceL2_n_11996), .B0(instanceL2_n_11395), .C0(
    instanceL2_n_11995));
  AND2X1 instanceL2_g10948(.Y(\instanceL2_prod_terms[1][15] [10]), .A(
    instanceL2_n_11995), .B(layer1_out[142]));
  MXI2XL instanceL2_g10949(.Y(\instanceL2_prod_terms[1][15] [8]), .A(
    instanceL2_n_11406), .B(layer1_out[140]), .S0(instanceL2_n_11996));
  ADDFX1 instanceL2_g10950(.CO(instanceL2_n_11994), .S(
    \instanceL2_prod_terms[6][15] [6]), .A(instanceL2_n_12021), .B(
    instanceL2_n_12018), .CI(instanceL2_n_11243));
  NAND2X1 instanceL2_g10951(.Y(instanceL2_n_11995), .A(instanceL2_n_12055), .B(
    instanceL2_n_11996));
  MX2XL instanceL2_g10952(.Y(\instanceL2_prod_terms[9][15] [9]), .A(
    instanceL2_n_11404), .B(layer1_out[141]), .S0(instanceL2_n_12001));
  XNOR2X1 instanceL2_g10953(.Y(\instanceL2_prod_terms[1][15] [7]), .A(
    instanceL2_n_12030), .B(instanceL2_n_11998));
  MX2XL instanceL2_g10954(.Y(\instanceL2_prod_terms[8][15] [9]), .A(
    layer1_out[142]), .B(instanceL2_n_11411), .S0(instanceL2_n_11997));
  OA22X1 instanceL2_g10955(.Y(instanceL2_n_11996), .A0(instanceL2_n_11391), .A1(
    instanceL2_n_11998), .B0(layer1_out[142]), .B1(instanceL2_n_11413));
  ADDFX1 instanceL2_g10956(.CO(instanceL2_n_11243), .S(
    \instanceL2_prod_terms[6][15] [5]), .A(instanceL2_n_12049), .B(
    instanceL2_n_12020), .CI(instanceL2_n_12004));
  AOI21X1 instanceL2_g10957(.Y(\instanceL2_prod_terms[9][15] [10]), .A0(
    instanceL2_n_11411), .A1(instanceL2_n_12000), .B0(
    \instanceL2_prod_terms[9][15] [11]));
  OAI2BB1X1 instanceL2_g10958(.Y(instanceL2_n_11997), .A0N(layer1_out[141]),
     .A1N(instanceL2_n_12005), .B0(instanceL2_n_11999));
  XNOR2X1 instanceL2_g10959(.Y(\instanceL2_prod_terms[1][15] [6]), .A(
    instanceL2_n_12029), .B(instanceL2_n_12002));
  AOI22X1 instanceL2_g10960(.Y(instanceL2_n_11998), .A0(instanceL2_n_11397), .A1(
    instanceL2_n_12002), .B0(instanceL2_n_11404), .B1(layer1_out[138]));
  OA21X1 instanceL2_g10961(.Y(\instanceL2_prod_terms[9][15] [8]), .A0(
    layer1_out[140]), .A1(instanceL2_n_12003), .B0(instanceL2_n_12001));
  NOR2X1 instanceL2_g10962(.Y(\instanceL2_prod_terms[9][15] [11]), .A(
    instanceL2_n_11411), .B(instanceL2_n_12000));
  INVX1 instanceL2_g10963(.Y(\instanceL2_prod_terms[8][15] [10]), .A(
    instanceL2_n_11999));
  XNOR2X1 instanceL2_g10964(.Y(\instanceL2_prod_terms[8][15] [8]), .A(
    instanceL2_n_11344), .B(instanceL2_n_12005));
  OAI21X1 instanceL2_g10965(.Y(instanceL2_n_11999), .A0(layer1_out[141]), .A1(
    instanceL2_n_12005), .B0(layer1_out[142]));
  NAND2BX1 instanceL2_g10966(.Y(instanceL2_n_12000), .AN(instanceL2_n_11395), .B(
    instanceL2_n_12003));
  NAND2X1 instanceL2_g10967(.Y(instanceL2_n_12001), .A(layer1_out[140]), .B(
    instanceL2_n_12003));
  XNOR2X1 instanceL2_g10968(.Y(\instanceL2_prod_terms[1][15] [5]), .A(
    instanceL2_n_12026), .B(instanceL2_n_12006));
  XNOR2X1 instanceL2_g10969(.Y(\instanceL2_prod_terms[8][15] [7]), .A(
    instanceL2_n_12036), .B(instanceL2_n_12007));
  OAI22X1 instanceL2_g10970(.Y(instanceL2_n_12002), .A0(instanceL2_n_11396), .A1(
    instanceL2_n_12006), .B0(layer1_out[140]), .B1(instanceL2_n_11409));
  ADDFX1 instanceL2_g10971(.CO(instanceL2_n_12004), .S(
    \instanceL2_prod_terms[6][15] [4]), .A(layer1_out[139]), .B(
    \instanceL2_prod_terms[9][15] [3]), .CI(instanceL2_n_12011));
  OAI2BB1X1 instanceL2_g10972(.Y(instanceL2_n_12003), .A0N(instanceL2_n_11389),
     .A1N(instanceL2_n_12009), .B0(instanceL2_n_12051));
  XNOR2X1 instanceL2_g10973(.Y(\instanceL2_prod_terms[9][15] [7]), .A(
    instanceL2_n_12030), .B(instanceL2_n_12009));
  OAI211X1 instanceL2_g10974(.Y(instanceL2_n_12005), .A0(instanceL2_n_12055),
     .A1(instanceL2_n_12008), .B0(instanceL2_n_11393), .C0(instanceL2_n_11395));
  NAND2X1 instanceL2_g10975(.Y(instanceL2_n_12007), .A(instanceL2_n_11393), .B(
    instanceL2_n_12008));
  AOI22X1 instanceL2_g10976(.Y(instanceL2_n_12006), .A0(instanceL2_n_12056), .A1(
    instanceL2_n_12010), .B0(instanceL2_n_11413), .B1(layer1_out[136]));
  XNOR2X1 instanceL2_g10977(.Y(\instanceL2_prod_terms[8][15] [5]), .A(
    instanceL2_n_12038), .B(instanceL2_n_12011));
  XNOR2X1 instanceL2_g10978(.Y(\instanceL2_prod_terms[8][15] [6]), .A(
    instanceL2_n_12031), .B(instanceL2_n_12012));
  XNOR2X1 instanceL2_g10979(.Y(\instanceL2_prod_terms[1][15] [4]), .A(
    instanceL2_n_12027), .B(instanceL2_n_12010));
  NAND2X1 instanceL2_g10980(.Y(instanceL2_n_12008), .A(instanceL2_n_12053), .B(
    instanceL2_n_12012));
  XNOR2X1 instanceL2_g10981(.Y(\instanceL2_prod_terms[9][15] [6]), .A(
    instanceL2_n_12029), .B(instanceL2_n_12013));
  OAI21X1 instanceL2_g10982(.Y(instanceL2_n_12009), .A0(instanceL2_n_12040), .A1(
    instanceL2_n_12013), .B0(instanceL2_n_12044));
  OAI21X1 instanceL2_g10983(.Y(instanceL2_n_12010), .A0(layer1_out[138]), .A1(
    instanceL2_n_12028), .B0(instanceL2_n_12049));
  OAI2BB1X1 instanceL2_g10984(.Y(instanceL2_n_12011), .A0N(instanceL2_n_12043),
     .A1N(instanceL2_n_11312), .B0(instanceL2_n_12048));
  XNOR2X1 instanceL2_g10985(.Y(\instanceL2_prod_terms[8][15] [4]), .A(
    instanceL2_n_11312), .B(instanceL2_n_12032));
  CLKXOR2X1 instanceL2_g10986(.Y(\instanceL2_prod_terms[1][15] [3]), .A(
    instanceL2_n_12028), .B(\instanceL2_prod_terms[9][15] [3]));
  OAI211X1 instanceL2_g10987(.Y(instanceL2_n_12012), .A0(instanceL2_n_12035),
     .A1(instanceL2_n_12017), .B0(instanceL2_n_12048), .C0(instanceL2_n_12045));
  NAND2XL instanceL2_g10988(.Y(instanceL2_n_12014), .A(instanceL2_n_12016), .B(
    instanceL2_n_12015));
  OAI21X1 instanceL2_g10989(.Y(instanceL2_n_12013), .A0(instanceL2_n_11372), .A1(
    instanceL2_n_12024), .B0(instanceL2_n_11387));
  XNOR2X1 instanceL2_g10990(.Y(\instanceL2_prod_terms[9][15] [5]), .A(
    instanceL2_n_12026), .B(instanceL2_n_12024));
  CLKXOR2X1 instanceL2_g10991(.Y(\instanceL2_prod_terms[8][15] [3]), .A(
    instanceL2_n_12050), .B(instanceL2_n_12039));
  INVX1 instanceL2_g10992(.Y(instanceL2_n_12017), .A(instanceL2_n_11312));
  OR2XL instanceL2_g10993(.Y(instanceL2_n_12015), .A(instanceL2_n_12030), .B(
    instanceL2_n_12023));
  NAND2X1 instanceL2_g10994(.Y(instanceL2_n_12016), .A(instanceL2_n_12030), .B(
    instanceL2_n_12023));
  NAND2XL instanceL2_g10995(.Y(instanceL2_n_11312), .A(instanceL2_n_12042), .B(
    instanceL2_n_12050));
  XNOR2X1 instanceL2_g10996(.Y(\instanceL2_prod_terms[9][15] [4]), .A(
    instanceL2_n_12047), .B(instanceL2_n_12027));
  MXI2XL instanceL2_g10997(.Y(instanceL2_n_12018), .A(instanceL2_n_11406), .B(
    layer1_out[140]), .S0(instanceL2_n_11370));
  MXI2XL instanceL2_g10998(.Y(instanceL2_n_12019), .A(layer1_out[142]), .B(
    instanceL2_n_11411), .S0(instanceL2_n_12029));
  MXI2XL instanceL2_g10999(.Y(instanceL2_n_12020), .A(instanceL2_n_11413), .B(
    layer1_out[139]), .S0(instanceL2_n_12037));
  OA21X1 instanceL2_g11000(.Y(\instanceL2_prod_terms[1][15] [2]), .A0(
    instanceL2_n_11409), .A1(instanceL2_n_12046), .B0(instanceL2_n_12028));
  OAI2BB1X1 instanceL2_g11001(.Y(instanceL2_n_12021), .A0N(instanceL2_n_12057),
     .A1N(instanceL2_n_12053), .B0(instanceL2_n_11393));
  NAND2BX1 instanceL2_g11002(.Y(instanceL2_n_12022), .AN(instanceL2_n_12034), .B(
    instanceL2_n_12033));
  OAI21X1 instanceL2_g11003(.Y(instanceL2_n_12025), .A0(layer1_out[137]), .A1(
    instanceL2_n_12055), .B0(instanceL2_n_11395));
  OAI21X1 instanceL2_g11004(.Y(instanceL2_n_12023), .A0(layer1_out[138]), .A1(
    instanceL2_n_12054), .B0(instanceL2_n_12052));
  OAI21X1 instanceL2_g11005(.Y(instanceL2_n_12024), .A0(instanceL2_n_12041), .A1(
    instanceL2_n_12047), .B0(instanceL2_n_11371));
  NOR2BX1 instanceL2_g11006(.Y(\instanceL2_prod_terms[1][15] [1]), .AN(
    instanceL2_n_12050), .B(instanceL2_n_12046));
  NAND2XL instanceL2_g11007(.Y(instanceL2_n_12031), .A(instanceL2_n_11393), .B(
    instanceL2_n_12053));
  NAND2BX1 instanceL2_g11008(.Y(instanceL2_n_11344), .AN(instanceL2_n_12054), .B(
    instanceL2_n_12052));
  NAND2XL instanceL2_g11009(.Y(instanceL2_n_12032), .A(instanceL2_n_12048), .B(
    instanceL2_n_12043));
  NAND2BX1 instanceL2_g11010(.Y(instanceL2_n_12026), .AN(instanceL2_n_11372), .B(
    instanceL2_n_11387));
  NOR2BX1 instanceL2_g11011(.Y(instanceL2_n_12027), .AN(instanceL2_n_11371), .B(
    instanceL2_n_12041));
  NAND2X1 instanceL2_g11012(.Y(instanceL2_n_12028), .A(instanceL2_n_11409), .B(
    instanceL2_n_12046));
  NOR2BX1 instanceL2_g11013(.Y(instanceL2_n_12029), .AN(instanceL2_n_12044), .B(
    instanceL2_n_12040));
  NAND2X1 instanceL2_g11014(.Y(instanceL2_n_12030), .A(instanceL2_n_12051), .B(
    instanceL2_n_11389));
  AOI21XL instanceL2_g11015(.Y(instanceL2_n_12035), .A0(layer1_out[139]), .A1(
    layer1_out[137]), .B0(layer1_out[138]));
  NAND2X1 instanceL2_g11016(.Y(instanceL2_n_12033), .A(instanceL2_n_11406), .B(
    instanceL2_n_11391));
  NAND2BX1 instanceL2_g11017(.Y(instanceL2_n_12036), .AN(instanceL2_n_12055), .B(
    instanceL2_n_11395));
  OAI22X1 instanceL2_g11018(.Y(instanceL2_n_12037), .A0(layer1_out[140]), .A1(
    layer1_out[136]), .B0(instanceL2_n_11406), .B1(instanceL2_n_12057));
  OAI21XL instanceL2_g11019(.Y(instanceL2_n_12038), .A0(layer1_out[138]), .A1(
    layer1_out[139]), .B0(instanceL2_n_12045));
  OAI2BB1X1 instanceL2_g11020(.Y(instanceL2_n_12039), .A0N(instanceL2_n_11409),
     .A1N(instanceL2_n_12057), .B0(instanceL2_n_12042));
  OAI22X1 instanceL2_g11021(.Y(instanceL2_n_11370), .A0(layer1_out[141]), .A1(
    layer1_out[137]), .B0(instanceL2_n_11404), .B1(instanceL2_n_11409));
  NOR2XL instanceL2_g11022(.Y(instanceL2_n_12034), .A(instanceL2_n_11406), .B(
    instanceL2_n_11391));
  OAI21X1 instanceL2_g11023(.Y(\instanceL2_prod_terms[9][15] [3]), .A0(
    instanceL2_n_12058), .A1(layer1_out[135]), .B0(instanceL2_n_12049));
  NAND2X1 instanceL2_g11024(.Y(instanceL2_n_11371), .A(layer1_out[136]), .B(
    layer1_out[139]));
  NOR2X1 instanceL2_g11025(.Y(instanceL2_n_11372), .A(instanceL2_n_11406), .B(
    instanceL2_n_11409));
  NOR2X1 instanceL2_g11026(.Y(instanceL2_n_12040), .A(layer1_out[141]), .B(
    layer1_out[138]));
  NOR2X1 instanceL2_g11027(.Y(instanceL2_n_12041), .A(layer1_out[136]), .B(
    layer1_out[139]));
  NAND2X1 instanceL2_g11028(.Y(instanceL2_n_12042), .A(layer1_out[137]), .B(
    layer1_out[136]));
  NAND2XL instanceL2_g11029(.Y(instanceL2_n_12043), .A(instanceL2_n_12058), .B(
    instanceL2_n_11409));
  NAND2XL instanceL2_g11030(.Y(instanceL2_n_12044), .A(layer1_out[141]), .B(
    layer1_out[138]));
  NAND2XL instanceL2_g11031(.Y(instanceL2_n_12045), .A(layer1_out[138]), .B(
    layer1_out[139]));
  NOR2X1 instanceL2_g11032(.Y(instanceL2_n_12046), .A(layer1_out[135]), .B(
    layer1_out[136]));
  NAND2X1 instanceL2_g11033(.Y(instanceL2_n_12047), .A(layer1_out[135]), .B(
    layer1_out[138]));
  NAND2X1 instanceL2_g11034(.Y(instanceL2_n_12048), .A(layer1_out[137]), .B(
    layer1_out[138]));
  NAND2X1 instanceL2_g11035(.Y(instanceL2_n_12049), .A(instanceL2_n_12058), .B(
    layer1_out[135]));
  NAND2X1 instanceL2_g11036(.Y(instanceL2_n_12050), .A(layer1_out[135]), .B(
    layer1_out[136]));
  NOR2XL instanceL2_g11037(.Y(instanceL2_n_11396), .A(layer1_out[137]), .B(
    instanceL2_n_11406));
  NAND2X1 instanceL2_g11038(.Y(instanceL2_n_11397), .A(instanceL2_n_12058), .B(
    layer1_out[141]));
  NAND2X1 instanceL2_g11039(.Y(instanceL2_n_12056), .A(layer1_out[139]), .B(
    instanceL2_n_12057));
  NAND2X1 instanceL2_g11040(.Y(instanceL2_n_12051), .A(layer1_out[142]), .B(
    layer1_out[139]));
  NAND2X1 instanceL2_g11041(.Y(instanceL2_n_11387), .A(instanceL2_n_11406), .B(
    instanceL2_n_11409));
  NAND2XL instanceL2_g11042(.Y(instanceL2_n_12052), .A(layer1_out[142]), .B(
    layer1_out[141]));
  NAND2X1 instanceL2_g11043(.Y(instanceL2_n_11389), .A(instanceL2_n_11411), .B(
    instanceL2_n_11413));
  NAND2X1 instanceL2_g11044(.Y(instanceL2_n_12053), .A(instanceL2_n_11406), .B(
    instanceL2_n_11413));
  NOR2X1 instanceL2_g11045(.Y(instanceL2_n_11391), .A(instanceL2_n_11411), .B(
    layer1_out[139]));
  NOR2X1 instanceL2_g11046(.Y(instanceL2_n_12054), .A(layer1_out[142]), .B(
    layer1_out[141]));
  NAND2X1 instanceL2_g11047(.Y(instanceL2_n_11393), .A(layer1_out[139]), .B(
    layer1_out[140]));
  NOR2X1 instanceL2_g11048(.Y(instanceL2_n_12055), .A(layer1_out[141]), .B(
    layer1_out[140]));
  NAND2X1 instanceL2_g11049(.Y(instanceL2_n_11395), .A(layer1_out[140]), .B(
    layer1_out[141]));
  INVX1 instanceL2_g11050(.Y(instanceL2_n_12057), .A(layer1_out[136]));
  INVX1 instanceL2_g11051(.Y(instanceL2_n_12058), .A(layer1_out[138]));
  INVX1 instanceL2_g11052(.Y(instanceL2_n_11404), .A(layer1_out[141]));
  INVX1 instanceL2_g11053(.Y(instanceL2_n_11406), .A(layer1_out[140]));
  INVX1 instanceL2_g11054(.Y(instanceL2_n_11409), .A(layer1_out[137]));
  INVX1 instanceL2_g11055(.Y(instanceL2_n_11411), .A(layer1_out[142]));
  INVX1 instanceL2_g11056(.Y(instanceL2_n_11413), .A(layer1_out[139]));
  XNOR2X1 instanceL2_g9594(.Y(\instanceL2_prod_terms[8][0] [10]), .A(
    instanceL2_n_10810), .B(instanceL2_n_10766));
  ADDFX1 instanceL2_g9595(.CO(instanceL2_n_10766), .S(
    \instanceL2_prod_terms[8][0] [9]), .A(instanceL2_n_10833), .B(
    instanceL2_n_12059), .CI(instanceL2_n_10768));
  ADDFX1 instanceL2_g9596(.CO(instanceL2_n_10768), .S(
    \instanceL2_prod_terms[8][0] [8]), .A(instanceL2_n_10827), .B(
    instanceL2_n_10805), .CI(instanceL2_n_10771));
  AOI21X1 instanceL2_g9597(.Y(\instanceL2_prod_terms[0][0][8] ), .A0(
    layer1_out[7]), .A1(instanceL2_n_10780), .B0(instanceL2_n_10773));
  ADDFX1 instanceL2_g9598(.CO(instanceL2_n_10771), .S(
    \instanceL2_prod_terms[8][0] [7]), .A(instanceL2_n_10802), .B(
    instanceL2_n_10804), .CI(instanceL2_n_10779));
  INVX1 instanceL2_g9599(.Y(\instanceL2_prod_terms[0][0][13] ), .A(
    instanceL2_n_10773));
  NOR2X1 instanceL2_g9600(.Y(instanceL2_n_10773), .A(layer1_out[7]), .B(
    instanceL2_n_10780));
  OA21X1 instanceL2_g9601(.Y(\instanceL2_prod_terms[0][0][7] ), .A0(
    instanceL2_n_12068), .A1(instanceL2_n_10787), .B0(instanceL2_n_10780));
  ADDFX1 instanceL2_g9602(.CO(instanceL2_n_10779), .S(
    \instanceL2_prod_terms[8][0] [6]), .A(instanceL2_n_10808), .B(
    instanceL2_n_10801), .CI(instanceL2_n_10786));
  NAND2X1 instanceL2_g9603(.Y(instanceL2_n_10780), .A(instanceL2_n_12068), .B(
    instanceL2_n_10787));
  AOI21X1 instanceL2_g9604(.Y(\instanceL2_prod_terms[0][0][6] ), .A0(
    layer1_out[5]), .A1(instanceL2_n_10795), .B0(instanceL2_n_10787));
  ADDFX1 instanceL2_g9605(.CO(instanceL2_n_10786), .S(
    \instanceL2_prod_terms[8][0] [5]), .A(instanceL2_n_12063), .B(
    instanceL2_n_10807), .CI(instanceL2_n_10793));
  NOR2X1 instanceL2_g9606(.Y(instanceL2_n_10787), .A(layer1_out[5]), .B(
    instanceL2_n_10795));
  OA21X1 instanceL2_g9607(.Y(\instanceL2_prod_terms[0][0][5] ), .A0(
    instanceL2_n_12066), .A1(instanceL2_n_10800), .B0(instanceL2_n_10795));
  ADDFX1 instanceL2_g9608(.CO(instanceL2_n_10793), .S(
    \instanceL2_prod_terms[8][0] [4]), .A(layer1_out[4]), .B(instanceL2_n_12061),
     .CI(\instanceL2_prod_terms[0][0][2] ));
  NAND2X1 instanceL2_g9609(.Y(instanceL2_n_10795), .A(instanceL2_n_12066), .B(
    instanceL2_n_10800));
  AOI21X1 instanceL2_g9610(.Y(\instanceL2_prod_terms[0][0][4] ), .A0(
    layer1_out[3]), .A1(instanceL2_n_10815), .B0(instanceL2_n_10800));
  ADDFX1 instanceL2_g9611(.CO(instanceL2_n_10802), .S(instanceL2_n_10801), .A(
    layer1_out[6]), .B(instanceL2_n_12067), .CI(layer1_out[3]));
  ADDFX1 instanceL2_g9612(.CO(instanceL2_n_10805), .S(instanceL2_n_10804), .A(
    layer1_out[7]), .B(instanceL2_n_12065), .CI(layer1_out[4]));
  ADDFX1 instanceL2_g9613(.CO(instanceL2_n_10808), .S(instanceL2_n_10807), .A(
    layer1_out[2]), .B(instanceL2_n_12064), .CI(layer1_out[5]));
  NOR2X1 instanceL2_g9614(.Y(instanceL2_n_10800), .A(layer1_out[3]), .B(
    instanceL2_n_10815));
  XNOR2X1 instanceL2_g9615(.Y(instanceL2_n_10810), .A(instanceL2_n_12062), .B(
    instanceL2_n_12070));
  OA21X1 instanceL2_g9616(.Y(\instanceL2_prod_terms[0][0][3] ), .A0(
    instanceL2_n_12067), .A1(instanceL2_n_12060), .B0(instanceL2_n_10815));
  AOI2BB1X1 instanceL2_g9617(.Y(\instanceL2_prod_terms[8][0] [3]), .A0N(
    layer1_out[0]), .A1N(layer1_out[3]), .B0(instanceL2_n_12061));
  NAND2X1 instanceL2_g9618(.Y(instanceL2_n_10815), .A(instanceL2_n_12067), .B(
    instanceL2_n_12060));
  OAI21X1 instanceL2_g9619(.Y(\instanceL2_prod_terms[0][0][2] ), .A0(
    instanceL2_n_12064), .A1(layer1_out[0]), .B0(instanceL2_n_12063));
  AOI21X1 instanceL2_g9620(.Y(instanceL2_n_12059), .A0(instanceL2_n_12068), .A1(
    layer1_out[5]), .B0(instanceL2_n_12062));
  OAI22X1 instanceL2_g9622(.Y(instanceL2_n_10827), .A0(layer1_out[5]), .A1(
    layer1_out[4]), .B0(instanceL2_n_12069), .B1(instanceL2_n_12066));
  NOR2XL instanceL2_g9623(.Y(instanceL2_n_12060), .A(layer1_out[1]), .B(
    layer1_out[0]));
  NOR2BX1 instanceL2_g9624(.Y(instanceL2_n_12061), .AN(layer1_out[0]), .B(
    instanceL2_n_12065));
  NOR2XL instanceL2_g9625(.Y(instanceL2_n_10833), .A(layer1_out[4]), .B(
    instanceL2_n_12069));
  NOR2X1 instanceL2_g9626(.Y(instanceL2_n_12062), .A(instanceL2_n_12068), .B(
    layer1_out[5]));
  NAND2X1 instanceL2_g9627(.Y(instanceL2_n_12063), .A(instanceL2_n_12064), .B(
    layer1_out[0]));
  INVX1 instanceL2_g9628(.Y(instanceL2_n_12064), .A(layer1_out[1]));
  INVX1 instanceL2_g9630(.Y(instanceL2_n_12065), .A(layer1_out[3]));
  INVX1 instanceL2_g9631(.Y(instanceL2_n_12066), .A(layer1_out[4]));
  INVX1 instanceL2_g9632(.Y(instanceL2_n_12067), .A(layer1_out[2]));
  INVX1 instanceL2_g9633(.Y(instanceL2_n_12068), .A(layer1_out[6]));
  INVX1 instanceL2_g9634(.Y(instanceL2_n_12069), .A(layer1_out[5]));
  MXI2XL instanceL2_g11057(.Y(instanceL2_n_12070), .A(layer1_out[6]), .B(
    instanceL2_n_12068), .S0(layer1_out[7]));
  XNOR2X1 instanceL2_g11058(.Y(\instanceL2_prod_terms[0][2][10] ), .A(
    layer1_out[26]), .B(instanceL2_n_12073));
  OAI211X1 instanceL2_g11059(.Y(\instanceL2_prod_terms[1][2][11] ), .A0(
    instanceL2_n_12135), .A1(instanceL2_n_12075), .B0(instanceL2_n_12136), .C0(
    instanceL2_n_12072));
  OAI21X1 instanceL2_g11060(.Y(\instanceL2_prod_terms[7][2] [8]), .A0(
    layer1_out[26]), .A1(instanceL2_n_11161), .B0(instanceL2_n_12071));
  NOR2X1 instanceL2_g11061(.Y(\instanceL2_prod_terms[1][2][12] ), .A(
    instanceL2_n_12145), .B(instanceL2_n_12074));
  OA21X1 instanceL2_g11062(.Y(instanceL2_n_12071), .A0(instanceL2_n_12136), .A1(
    instanceL2_n_12081), .B0(instanceL2_n_12135));
  MXI2XL instanceL2_g11063(.Y(\instanceL2_prod_terms[1][2][10] ), .A(
    layer1_out[25]), .B(instanceL2_n_12145), .S0(instanceL2_n_12075));
  OAI22X1 instanceL2_g11064(.Y(\instanceL2_prod_terms[7][2] [7]), .A0(
    instanceL2_n_12145), .A1(instanceL2_n_12081), .B0(layer1_out[25]), .B1(
    instanceL2_n_11161));
  XNOR2X1 instanceL2_g11065(.Y(\instanceL2_prod_terms[0][2][9] ), .A(
    instanceL2_n_12107), .B(instanceL2_n_11162));
  NAND2X1 instanceL2_g11066(.Y(instanceL2_n_12072), .A(layer1_out[26]), .B(
    instanceL2_n_12075));
  OAI21X1 instanceL2_g11067(.Y(instanceL2_n_12073), .A0(layer1_out[25]), .A1(
    instanceL2_n_12076), .B0(instanceL2_n_12114));
  OR3X1 instanceL2_g11068(.Y(\instanceL2_prod_terms[7][2] [13]), .A(
    layer1_out[26]), .B(layer1_out[25]), .C(instanceL2_n_12081));
  AOI21X1 instanceL2_g11069(.Y(instanceL2_n_12074), .A0(layer1_out[26]), .A1(
    instanceL2_n_12078), .B0(instanceL2_n_12115));
  MX2XL instanceL2_g11070(.Y(\instanceL2_prod_terms[1][2][9] ), .A(
    layer1_out[24]), .B(instanceL2_n_12148), .S0(instanceL2_n_12077));
  INVX1 instanceL2_g11071(.Y(instanceL2_n_11161), .A(instanceL2_n_12081));
  NAND2X1 instanceL2_g11072(.Y(instanceL2_n_11162), .A(instanceL2_n_12104), .B(
    instanceL2_n_12076));
  XNOR2X1 instanceL2_g11073(.Y(\instanceL2_prod_terms[0][2][8] ), .A(
    instanceL2_n_12100), .B(instanceL2_n_12079));
  NOR2X1 instanceL2_g11074(.Y(instanceL2_n_12075), .A(instanceL2_n_12115), .B(
    instanceL2_n_12078));
  NAND2X1 instanceL2_g11075(.Y(instanceL2_n_12077), .A(instanceL2_n_12130), .B(
    instanceL2_n_12080));
  NAND2X1 instanceL2_g11076(.Y(instanceL2_n_12076), .A(instanceL2_n_12103), .B(
    instanceL2_n_12079));
  OA21X1 instanceL2_g11077(.Y(\instanceL2_prod_terms[8][2] [8]), .A0(
    instanceL2_n_12148), .A1(instanceL2_n_12083), .B0(instanceL2_n_12081));
  XNOR2X1 instanceL2_g11078(.Y(\instanceL2_prod_terms[1][2][8] ), .A(
    instanceL2_n_12118), .B(instanceL2_n_12082));
  NOR2X1 instanceL2_g11079(.Y(instanceL2_n_12078), .A(instanceL2_n_12148), .B(
    instanceL2_n_12080));
  ADDFX1 instanceL2_g11080(.CO(instanceL2_n_12079), .S(
    \instanceL2_prod_terms[0][2][7] ), .A(instanceL2_n_12139), .B(
    instanceL2_n_12117), .CI(instanceL2_n_12084));
  NAND2X1 instanceL2_g11081(.Y(instanceL2_n_12080), .A(instanceL2_n_12129), .B(
    instanceL2_n_12082));
  NAND2X1 instanceL2_g11082(.Y(instanceL2_n_12081), .A(instanceL2_n_12148), .B(
    instanceL2_n_12083));
  ADDFX1 instanceL2_g11083(.CO(instanceL2_n_12082), .S(
    \instanceL2_prod_terms[1][2][7] ), .A(layer1_out[25]), .B(layer1_out[22]),
     .CI(instanceL2_n_12085));
  AOI21X1 instanceL2_g11084(.Y(\instanceL2_prod_terms[8][2] [7]), .A0(
    layer1_out[23]), .A1(instanceL2_n_12087), .B0(instanceL2_n_12083));
  ADDFX1 instanceL2_g11085(.CO(instanceL2_n_12084), .S(
    \instanceL2_prod_terms[0][2][6] ), .A(instanceL2_n_12142), .B(
    instanceL2_n_12110), .CI(instanceL2_n_12088));
  NOR2X1 instanceL2_g11086(.Y(instanceL2_n_12083), .A(layer1_out[23]), .B(
    instanceL2_n_12087));
  OAI211X1 instanceL2_g11087(.Y(\instanceL2_prod_terms[4][2] [11]), .A0(
    instanceL2_n_12135), .A1(instanceL2_n_12090), .B0(instanceL2_n_12136), .C0(
    instanceL2_n_11198));
  MX2XL instanceL2_g11088(.Y(\instanceL2_prod_terms[4][2] [10]), .A(
    instanceL2_n_12145), .B(layer1_out[25]), .S0(instanceL2_n_11200));
  ADDFX1 instanceL2_g11089(.CO(instanceL2_n_12085), .S(
    \instanceL2_prod_terms[1][2][6] ), .A(layer1_out[24]), .B(layer1_out[21]),
     .CI(instanceL2_n_12091));
  XNOR2X1 instanceL2_g11090(.Y(\instanceL2_prod_terms[4][2] [9]), .A(
    instanceL2_n_12116), .B(instanceL2_n_12089));
  NAND2X1 instanceL2_g11091(.Y(instanceL2_n_11198), .A(layer1_out[26]), .B(
    instanceL2_n_12090));
  AOI21X1 instanceL2_g11092(.Y(instanceL2_n_11200), .A0(instanceL2_n_12137), .A1(
    instanceL2_n_12092), .B0(instanceL2_n_12106));
  INVX1 instanceL2_g11093(.Y(\instanceL2_prod_terms[4][2] [12]), .A(
    instanceL2_n_12086));
  OA21X1 instanceL2_g11094(.Y(\instanceL2_prod_terms[8][2] [6]), .A0(
    instanceL2_n_12144), .A1(instanceL2_n_12095), .B0(instanceL2_n_12087));
  OAI211X1 instanceL2_g11095(.Y(instanceL2_n_12086), .A0(instanceL2_n_12106),
     .A1(instanceL2_n_12093), .B0(layer1_out[26]), .C0(layer1_out[25]));
  ADDFX1 instanceL2_g11096(.CO(instanceL2_n_12088), .S(
    \instanceL2_prod_terms[0][2][5] ), .A(instanceL2_n_12140), .B(
    instanceL2_n_12111), .CI(instanceL2_n_12094));
  NAND2BX1 instanceL2_g11097(.Y(instanceL2_n_12089), .AN(instanceL2_n_12092), .B(
    instanceL2_n_12133));
  NAND2X1 instanceL2_g11098(.Y(instanceL2_n_12087), .A(instanceL2_n_12144), .B(
    instanceL2_n_12095));
  XNOR2X1 instanceL2_g11099(.Y(\instanceL2_prod_terms[4][2] [8]), .A(
    instanceL2_n_12117), .B(instanceL2_n_12093));
  AOI21X1 instanceL2_g11100(.Y(instanceL2_n_12090), .A0(instanceL2_n_12137), .A1(
    instanceL2_n_12093), .B0(instanceL2_n_12106));
  ADDFX1 instanceL2_g11101(.CO(instanceL2_n_12091), .S(
    \instanceL2_prod_terms[1][2][5] ), .A(layer1_out[23]), .B(layer1_out[20]),
     .CI(instanceL2_n_12098));
  NOR2BX1 instanceL2_g11102(.Y(instanceL2_n_12092), .AN(instanceL2_n_12093), .B(
    instanceL2_n_12132));
  AOI21X1 instanceL2_g11103(.Y(\instanceL2_prod_terms[8][2] [5]), .A0(
    layer1_out[21]), .A1(instanceL2_n_12099), .B0(instanceL2_n_12095));
  XNOR2X1 instanceL2_g11104(.Y(\instanceL2_prod_terms[4][2] [7]), .A(
    instanceL2_n_12110), .B(instanceL2_n_12097));
  OAI21X1 instanceL2_g11105(.Y(instanceL2_n_12093), .A0(instanceL2_n_12121), .A1(
    instanceL2_n_12096), .B0(instanceL2_n_12120));
  ADDFX1 instanceL2_g11106(.CO(instanceL2_n_12094), .S(
    \instanceL2_prod_terms[0][2][4] ), .A(instanceL2_n_12141), .B(
    instanceL2_n_12112), .CI(instanceL2_n_12108));
  NOR2X1 instanceL2_g11107(.Y(instanceL2_n_12095), .A(layer1_out[21]), .B(
    instanceL2_n_12099));
  INVX1 instanceL2_g11108(.Y(instanceL2_n_12096), .A(instanceL2_n_12097));
  ADDFX1 instanceL2_g11109(.CO(instanceL2_n_12098), .S(
    \instanceL2_prod_terms[1][2][4] ), .A(layer1_out[22]), .B(layer1_out[19]),
     .CI(instanceL2_n_12128));
  OAI2BB1X1 instanceL2_g11110(.Y(instanceL2_n_12097), .A0N(instanceL2_n_12124),
     .A1N(instanceL2_n_12101), .B0(instanceL2_n_12119));
  XNOR2X1 instanceL2_g11111(.Y(\instanceL2_prod_terms[4][2] [6]), .A(
    instanceL2_n_12111), .B(instanceL2_n_12101));
  XNOR2X1 instanceL2_g11112(.Y(\instanceL2_prod_terms[0][2][3] ), .A(
    instanceL2_n_11306), .B(instanceL2_n_12102));
  OA21X1 instanceL2_g11113(.Y(\instanceL2_prod_terms[8][2] [4]), .A0(
    instanceL2_n_12146), .A1(instanceL2_n_12127), .B0(instanceL2_n_12099));
  XNOR2X1 instanceL2_g11114(.Y(\instanceL2_prod_terms[4][2] [5]), .A(
    instanceL2_n_12112), .B(instanceL2_n_12105));
  NAND2XL instanceL2_g11115(.Y(instanceL2_n_12100), .A(instanceL2_n_12104), .B(
    instanceL2_n_12103));
  NAND2X1 instanceL2_g11116(.Y(instanceL2_n_12099), .A(instanceL2_n_12146), .B(
    instanceL2_n_12127));
  XNOR2X1 instanceL2_g11117(.Y(\instanceL2_prod_terms[4][2] [4]), .A(
    instanceL2_n_11305), .B(instanceL2_n_12113));
  MXI2XL instanceL2_g11118(.Y(instanceL2_n_12102), .A(instanceL2_n_12146), .B(
    layer1_out[20]), .S0(instanceL2_n_12113));
  OAI211X1 instanceL2_g11119(.Y(instanceL2_n_12101), .A0(instanceL2_n_12126),
     .A1(instanceL2_n_12125), .B0(instanceL2_n_12123), .C0(instanceL2_n_12109));
  NAND2X1 instanceL2_g11120(.Y(instanceL2_n_12105), .A(instanceL2_n_12126), .B(
    instanceL2_n_12109));
  OR2XL instanceL2_g11121(.Y(instanceL2_n_12103), .A(instanceL2_n_12131), .B(
    instanceL2_n_12116));
  NAND2X1 instanceL2_g11122(.Y(instanceL2_n_12104), .A(instanceL2_n_12131), .B(
    instanceL2_n_12116));
  OAI211X1 instanceL2_g11123(.Y(instanceL2_n_12107), .A0(instanceL2_n_12145),
     .A1(instanceL2_n_12148), .B0(instanceL2_n_12135), .C0(instanceL2_n_12114));
  AOI2BB1X1 instanceL2_g11124(.Y(instanceL2_n_12108), .A0N(layer1_out[20]), .A1N(
    instanceL2_n_11306), .B0(instanceL2_n_12113));
  OAI21X1 instanceL2_g11125(.Y(instanceL2_n_12106), .A0(instanceL2_n_12133), .A1(
    instanceL2_n_12138), .B0(instanceL2_n_12134));
  NOR2BX1 instanceL2_g11126(.Y(\instanceL2_prod_terms[4][2] [3]), .AN(
    instanceL2_n_11305), .B(instanceL2_n_11306));
  OR2X1 instanceL2_g11127(.Y(instanceL2_n_12109), .A(instanceL2_n_12122), .B(
    instanceL2_n_11305));
  NAND2BX1 instanceL2_g11128(.Y(instanceL2_n_12110), .AN(instanceL2_n_12121), .B(
    instanceL2_n_12120));
  NAND2X1 instanceL2_g11129(.Y(instanceL2_n_12111), .A(instanceL2_n_12119), .B(
    instanceL2_n_12124));
  NAND2BX1 instanceL2_g11130(.Y(instanceL2_n_12112), .AN(instanceL2_n_12125), .B(
    instanceL2_n_12123));
  NOR2BX1 instanceL2_g11131(.Y(instanceL2_n_12113), .AN(instanceL2_n_12126), .B(
    instanceL2_n_12122));
  AOI2BB1X1 instanceL2_g11132(.Y(\instanceL2_prod_terms[1][2][3] ), .A0N(
    layer1_out[18]), .A1N(layer1_out[21]), .B0(instanceL2_n_12128));
  AOI21X1 instanceL2_g11133(.Y(\instanceL2_prod_terms[7][2] [1]), .A0(
    layer1_out[19]), .A1(layer1_out[18]), .B0(instanceL2_n_12127));
  OR2X1 instanceL2_g11134(.Y(instanceL2_n_12114), .A(layer1_out[24]), .B(
    instanceL2_n_12136));
  NAND2XL instanceL2_g11135(.Y(instanceL2_n_12118), .A(instanceL2_n_12130), .B(
    instanceL2_n_12129));
  NOR2X1 instanceL2_g11136(.Y(instanceL2_n_12115), .A(instanceL2_n_12147), .B(
    instanceL2_n_12134));
  NAND2X1 instanceL2_g11137(.Y(instanceL2_n_12116), .A(instanceL2_n_12134), .B(
    instanceL2_n_12137));
  NAND2BX1 instanceL2_g11138(.Y(instanceL2_n_12117), .AN(instanceL2_n_12132), .B(
    instanceL2_n_12133));
  NAND2X1 instanceL2_g11139(.Y(instanceL2_n_12119), .A(layer1_out[21]), .B(
    layer1_out[23]));
  NAND2X1 instanceL2_g11140(.Y(instanceL2_n_12120), .A(layer1_out[24]), .B(
    layer1_out[22]));
  NOR2X1 instanceL2_g11141(.Y(instanceL2_n_12121), .A(layer1_out[24]), .B(
    layer1_out[22]));
  NOR2XL instanceL2_g11142(.Y(instanceL2_n_12122), .A(layer1_out[21]), .B(
    layer1_out[19]));
  NAND2X1 instanceL2_g11143(.Y(instanceL2_n_12123), .A(layer1_out[20]), .B(
    layer1_out[22]));
  NAND2X1 instanceL2_g11144(.Y(instanceL2_n_12124), .A(instanceL2_n_12147), .B(
    instanceL2_n_12143));
  NOR2XL instanceL2_g11145(.Y(instanceL2_n_12125), .A(layer1_out[22]), .B(
    layer1_out[20]));
  NAND2X1 instanceL2_g11146(.Y(instanceL2_n_12126), .A(layer1_out[19]), .B(
    layer1_out[21]));
  NOR2X1 instanceL2_g11147(.Y(instanceL2_n_12127), .A(layer1_out[18]), .B(
    layer1_out[19]));
  NAND2XL instanceL2_g11148(.Y(instanceL2_n_11305), .A(layer1_out[18]), .B(
    layer1_out[20]));
  NOR2XL instanceL2_g11149(.Y(instanceL2_n_11306), .A(layer1_out[20]), .B(
    layer1_out[18]));
  AND2XL instanceL2_g11150(.Y(instanceL2_n_12128), .A(layer1_out[21]), .B(
    layer1_out[18]));
  INVX1 instanceL2_g11151(.Y(instanceL2_n_12137), .A(instanceL2_n_12138));
  NAND2X1 instanceL2_g11152(.Y(instanceL2_n_12129), .A(instanceL2_n_12149), .B(
    instanceL2_n_12147));
  NAND2X1 instanceL2_g11153(.Y(instanceL2_n_12130), .A(layer1_out[26]), .B(
    layer1_out[23]));
  NOR2XL instanceL2_g11154(.Y(instanceL2_n_12131), .A(layer1_out[23]), .B(
    instanceL2_n_12145));
  NOR2X1 instanceL2_g11155(.Y(instanceL2_n_12139), .A(layer1_out[22]), .B(
    instanceL2_n_12148));
  NOR2XL instanceL2_g11156(.Y(instanceL2_n_12132), .A(layer1_out[25]), .B(
    layer1_out[23]));
  NOR2X1 instanceL2_g11157(.Y(instanceL2_n_12140), .A(layer1_out[20]), .B(
    instanceL2_n_12144));
  NOR2X1 instanceL2_g11158(.Y(instanceL2_n_12141), .A(layer1_out[19]), .B(
    instanceL2_n_12143));
  NOR2X1 instanceL2_g11159(.Y(instanceL2_n_12142), .A(layer1_out[21]), .B(
    instanceL2_n_12147));
  NAND2X1 instanceL2_g11160(.Y(instanceL2_n_12133), .A(layer1_out[25]), .B(
    layer1_out[23]));
  NAND2X1 instanceL2_g11161(.Y(instanceL2_n_12134), .A(layer1_out[26]), .B(
    layer1_out[24]));
  NAND2X1 instanceL2_g11162(.Y(instanceL2_n_12135), .A(instanceL2_n_12149), .B(
    layer1_out[25]));
  NAND2XL instanceL2_g11163(.Y(instanceL2_n_12136), .A(layer1_out[26]), .B(
    instanceL2_n_12145));
  NOR2X1 instanceL2_g11164(.Y(instanceL2_n_12138), .A(layer1_out[26]), .B(
    layer1_out[24]));
  INVX1 instanceL2_g11165(.Y(instanceL2_n_12143), .A(layer1_out[21]));
  INVX1 instanceL2_g11166(.Y(instanceL2_n_12144), .A(layer1_out[22]));
  INVX1 instanceL2_g11167(.Y(instanceL2_n_12145), .A(layer1_out[25]));
  INVX1 instanceL2_g11168(.Y(instanceL2_n_12146), .A(layer1_out[20]));
  INVX1 instanceL2_g11169(.Y(instanceL2_n_12147), .A(layer1_out[23]));
  INVX1 instanceL2_g11170(.Y(instanceL2_n_12148), .A(layer1_out[24]));
  INVX1 instanceL2_g11171(.Y(instanceL2_n_12149), .A(layer1_out[26]));
  OAI21X1 instanceL2_g9580(.Y(\instanceL2_prod_terms[2][13] [9]), .A0(
    instanceL2_n_12177), .A1(instanceL2_n_10770), .B0(instanceL2_n_12150));
  AND2XL instanceL2_g9581(.Y(\instanceL2_prod_terms[2][13] [10]), .A(
    layer1_out[124]), .B(instanceL2_n_12150));
  AO21X1 instanceL2_g9582(.Y(\instanceL2_prod_terms[2][13] [8]), .A0(
    layer1_out[122]), .A1(instanceL2_n_10772), .B0(instanceL2_n_10770));
  NAND2BX1 instanceL2_g9583(.Y(instanceL2_n_12150), .AN(instanceL2_n_10772), .B(
    instanceL2_n_12167));
  NOR2X1 instanceL2_g9584(.Y(instanceL2_n_10770), .A(layer1_out[122]), .B(
    instanceL2_n_10772));
  ADDFX1 instanceL2_g9585(.CO(instanceL2_n_10772), .S(
    \instanceL2_prod_terms[2][13] [7]), .A(layer1_out[121]), .B(
    instanceL2_n_12176), .CI(instanceL2_n_10775));
  ADDFX1 instanceL2_g9586(.CO(instanceL2_n_10775), .S(
    \instanceL2_prod_terms[2][13] [6]), .A(instanceL2_n_12177), .B(
    layer1_out[120]), .CI(instanceL2_n_10785));
  AOI2BB1XL instanceL2_g9587(.Y(\instanceL2_prod_terms[6][13] [8]), .A0N(
    layer1_out[124]), .A1N(instanceL2_n_10783), .B0(
    \instanceL2_prod_terms[6][13] [9]));
  AND2XL instanceL2_g9588(.Y(\instanceL2_prod_terms[6][13] [9]), .A(
    layer1_out[124]), .B(instanceL2_n_10783));
  XNOR2X1 instanceL2_g9589(.Y(\instanceL2_prod_terms[6][13] [7]), .A(
    instanceL2_n_10845), .B(instanceL2_n_12151));
  OAI211X1 instanceL2_g9590(.Y(instanceL2_n_10783), .A0(instanceL2_n_12165), .A1(
    instanceL2_n_10794), .B0(instanceL2_n_10858), .C0(instanceL2_n_12171));
  ADDFX1 instanceL2_g9591(.CO(instanceL2_n_10785), .S(
    \instanceL2_prod_terms[2][13] [5]), .A(layer1_out[119]), .B(
    instanceL2_n_12180), .CI(instanceL2_n_12153));
  NAND2X1 instanceL2_g9592(.Y(instanceL2_n_12151), .A(instanceL2_n_10858), .B(
    instanceL2_n_10794));
  XNOR2X1 instanceL2_g9593(.Y(\instanceL2_prod_terms[5][13] [8]), .A(
    layer1_out[123]), .B(instanceL2_n_10811));
  XNOR2X1 instanceL2_g11172(.Y(\instanceL2_prod_terms[6][13] [6]), .A(
    instanceL2_n_12160), .B(instanceL2_n_12152));
  NAND2X1 instanceL2_g11173(.Y(\instanceL2_prod_terms[9][13] [13]), .A(
    instanceL2_n_12165), .B(instanceL2_n_10811));
  XNOR2X1 instanceL2_g11174(.Y(\instanceL2_prod_terms[6][13] [5]), .A(
    instanceL2_n_12158), .B(instanceL2_n_10806));
  NAND2BX1 instanceL2_g11175(.Y(instanceL2_n_10794), .AN(instanceL2_n_12167), .B(
    instanceL2_n_12152));
  OAI21X1 instanceL2_g11176(.Y(\instanceL2_prod_terms[5][13] [5]), .A0(
    layer1_out[120]), .A1(instanceL2_n_12162), .B0(instanceL2_n_10820));
  XNOR2X1 instanceL2_g11177(.Y(\instanceL2_prod_terms[9][13] [8]), .A(
    instanceL2_n_12176), .B(instanceL2_n_10812));
  OAI211X1 instanceL2_g11178(.Y(instanceL2_n_12152), .A0(instanceL2_n_10856),
     .A1(instanceL2_n_10814), .B0(instanceL2_n_12164), .C0(instanceL2_n_12172));
  ADDFX1 instanceL2_g11179(.CO(instanceL2_n_12153), .S(
    \instanceL2_prod_terms[2][13] [4]), .A(layer1_out[118]), .B(
    instanceL2_n_12178), .CI(instanceL2_n_12155));
  NAND2X1 instanceL2_g11180(.Y(instanceL2_n_10806), .A(instanceL2_n_12164), .B(
    instanceL2_n_10814));
  AOI21X1 instanceL2_g11181(.Y(\instanceL2_prod_terms[5][13] [7]), .A0(
    layer1_out[122]), .A1(instanceL2_n_10821), .B0(instanceL2_n_10811));
  XNOR2X1 instanceL2_g11182(.Y(\instanceL2_prod_terms[6][13] [4]), .A(
    instanceL2_n_12163), .B(instanceL2_n_12154));
  NAND2BX1 instanceL2_g11183(.Y(instanceL2_n_10812), .AN(instanceL2_n_10821), .B(
    instanceL2_n_12167));
  NOR2X1 instanceL2_g11184(.Y(instanceL2_n_10811), .A(layer1_out[122]), .B(
    instanceL2_n_10821));
  OAI21X1 instanceL2_g11185(.Y(\instanceL2_prod_terms[2][13] [3]), .A0(
    instanceL2_n_12161), .A1(instanceL2_n_12162), .B0(instanceL2_n_10820));
  XNOR2X1 instanceL2_g11186(.Y(\instanceL2_prod_terms[6][13] [3]), .A(
    instanceL2_n_12156), .B(instanceL2_n_12159));
  NAND2BX1 instanceL2_g11187(.Y(instanceL2_n_10814), .AN(instanceL2_n_12166), .B(
    instanceL2_n_12154));
  NAND2X1 instanceL2_g11188(.Y(instanceL2_n_10820), .A(instanceL2_n_12161), .B(
    instanceL2_n_12162));
  NAND2X1 instanceL2_g11189(.Y(instanceL2_n_10821), .A(instanceL2_n_12166), .B(
    instanceL2_n_12162));
  XOR2XL instanceL2_g11190(.Y(\instanceL2_prod_terms[6][13] [2]), .A(
    instanceL2_n_12168), .B(instanceL2_n_10853));
  OAI211X1 instanceL2_g11191(.Y(instanceL2_n_12154), .A0(instanceL2_n_12168),
     .A1(instanceL2_n_12174), .B0(instanceL2_n_12173), .C0(instanceL2_n_12170));
  NAND2X1 instanceL2_g11192(.Y(instanceL2_n_12155), .A(instanceL2_n_12169), .B(
    instanceL2_n_12157));
  XNOR2X1 instanceL2_g11193(.Y(\instanceL2_prod_terms[5][13] [6]), .A(
    instanceL2_n_12178), .B(instanceL2_n_12157));
  NAND2XL instanceL2_g11194(.Y(instanceL2_n_12156), .A(instanceL2_n_12173), .B(
    instanceL2_n_12168));
  AOI21X1 instanceL2_g11195(.Y(\instanceL2_prod_terms[2][13] [2]), .A0(
    layer1_out[119]), .A1(instanceL2_n_12175), .B0(instanceL2_n_12162));
  NAND2BXL instanceL2_g11196(.Y(instanceL2_n_12158), .AN(instanceL2_n_10856), .B(
    instanceL2_n_12172));
  NAND2BX1 instanceL2_g11197(.Y(instanceL2_n_12159), .AN(instanceL2_n_12174), .B(
    instanceL2_n_12170));
  NAND2BX1 instanceL2_g11198(.Y(instanceL2_n_10845), .AN(instanceL2_n_12165), .B(
    instanceL2_n_12171));
  NAND2BX1 instanceL2_g9621(.Y(instanceL2_n_12160), .AN(instanceL2_n_12167), .B(
    instanceL2_n_10858));
  NAND2BX1 instanceL2_g11199(.Y(instanceL2_n_12157), .AN(instanceL2_n_12175), .B(
    instanceL2_n_12174));
  AND2X1 instanceL2_g11200(.Y(\instanceL2_prod_terms[2][13] [1]), .A(
    instanceL2_n_12175), .B(instanceL2_n_12168));
  OAI21X1 instanceL2_g11201(.Y(instanceL2_n_12161), .A0(instanceL2_n_12179), .A1(
    layer1_out[117]), .B0(instanceL2_n_12169));
  OAI21X1 instanceL2_g11202(.Y(instanceL2_n_10853), .A0(layer1_out[119]), .A1(
    layer1_out[118]), .B0(instanceL2_n_12173));
  NAND2BXL instanceL2_g11203(.Y(instanceL2_n_12163), .AN(instanceL2_n_12166), .B(
    instanceL2_n_12164));
  NOR2X1 instanceL2_g11204(.Y(instanceL2_n_12162), .A(layer1_out[119]), .B(
    instanceL2_n_12175));
  NOR2XL instanceL2_g11205(.Y(instanceL2_n_10856), .A(layer1_out[122]), .B(
    layer1_out[121]));
  NAND2X1 instanceL2_g9629(.Y(instanceL2_n_12164), .A(layer1_out[120]), .B(
    layer1_out[121]));
  NAND2X1 instanceL2_g11206(.Y(instanceL2_n_10858), .A(layer1_out[122]), .B(
    layer1_out[123]));
  NOR2X1 instanceL2_g11207(.Y(instanceL2_n_12165), .A(layer1_out[123]), .B(
    layer1_out[124]));
  NOR2X1 instanceL2_g11208(.Y(instanceL2_n_12166), .A(layer1_out[120]), .B(
    layer1_out[121]));
  NOR2X1 instanceL2_g11209(.Y(instanceL2_n_12167), .A(layer1_out[122]), .B(
    layer1_out[123]));
  NAND2XL instanceL2_g11210(.Y(instanceL2_n_12168), .A(layer1_out[118]), .B(
    layer1_out[117]));
  NAND2X1 instanceL2_g9635(.Y(instanceL2_n_12169), .A(instanceL2_n_12179), .B(
    layer1_out[117]));
  NAND2XL instanceL2_g9636(.Y(instanceL2_n_12170), .A(layer1_out[119]), .B(
    layer1_out[120]));
  NAND2XL instanceL2_g9637(.Y(instanceL2_n_12171), .A(layer1_out[124]), .B(
    layer1_out[123]));
  NAND2XL instanceL2_g9638(.Y(instanceL2_n_12172), .A(layer1_out[121]), .B(
    layer1_out[122]));
  NAND2XL instanceL2_g9639(.Y(instanceL2_n_12173), .A(layer1_out[118]), .B(
    layer1_out[119]));
  NOR2X1 instanceL2_g9640(.Y(instanceL2_n_12174), .A(layer1_out[119]), .B(
    layer1_out[120]));
  OR2X1 instanceL2_g9641(.Y(instanceL2_n_12175), .A(layer1_out[118]), .B(
    layer1_out[117]));
  INVX1 instanceL2_g9642(.Y(instanceL2_n_12176), .A(layer1_out[124]));
  INVX1 instanceL2_g9643(.Y(instanceL2_n_12177), .A(layer1_out[123]));
  INVX1 instanceL2_g9644(.Y(instanceL2_n_12178), .A(layer1_out[121]));
  INVX1 instanceL2_g9645(.Y(instanceL2_n_12179), .A(layer1_out[120]));
  INVX1 instanceL2_g9646(.Y(instanceL2_n_12180), .A(layer1_out[122]));
  AOI2BB1X1 instanceL2_g9847(.Y(\instanceL2_prod_terms[9][3] [10]), .A0N(
    layer1_out[34]), .A1N(instanceL2_n_12183), .B0(
    \instanceL2_prod_terms[9][3] [11]));
  AND2XL instanceL2_g9848(.Y(\instanceL2_prod_terms[9][3] [11]), .A(
    layer1_out[34]), .B(instanceL2_n_12183));
  MX2X1 instanceL2_g9849(.Y(\instanceL2_prod_terms[0][3][9] ), .A(
    instanceL2_n_12186), .B(instanceL2_n_12182), .S0(layer1_out[34]));
  AOI21X1 instanceL2_g9850(.Y(\instanceL2_prod_terms[2][3] [7]), .A0(
    layer1_out[34]), .A1(instanceL2_n_12186), .B0(instanceL2_n_12181));
  AOI21X1 instanceL2_g9851(.Y(\instanceL2_prod_terms[9][3] [9]), .A0(
    instanceL2_n_12227), .A1(instanceL2_n_12184), .B0(instanceL2_n_12183));
  INVX1 instanceL2_g9852(.Y(instanceL2_n_12181), .A(
    \instanceL2_prod_terms[2][3] [13]));
  ADDFX1 instanceL2_g9853(.CO(instanceL2_n_12182), .S(
    \instanceL2_prod_terms[0][3][8] ), .A(instanceL2_n_12227), .B(
    instanceL2_n_12226), .CI(instanceL2_n_12185));
  OR2X1 instanceL2_g9854(.Y(\instanceL2_prod_terms[2][3] [13]), .A(
    layer1_out[34]), .B(instanceL2_n_12186));
  NOR2X1 instanceL2_g9855(.Y(instanceL2_n_12183), .A(instanceL2_n_12227), .B(
    instanceL2_n_12184));
  OA21X1 instanceL2_g9856(.Y(\instanceL2_prod_terms[9][3] [8]), .A0(
    layer1_out[32]), .A1(instanceL2_n_12187), .B0(instanceL2_n_12184));
  OA21X1 instanceL2_g9857(.Y(\instanceL2_prod_terms[2][3] [6]), .A0(
    instanceL2_n_12227), .A1(instanceL2_n_12188), .B0(instanceL2_n_12186));
  ADDFX1 instanceL2_g9858(.CO(instanceL2_n_12185), .S(
    \instanceL2_prod_terms[0][3][7] ), .A(instanceL2_n_10988), .B(
    instanceL2_n_12207), .CI(instanceL2_n_12189));
  NAND2X1 instanceL2_g9859(.Y(instanceL2_n_12184), .A(layer1_out[32]), .B(
    instanceL2_n_12187));
  AOI21X1 instanceL2_g9860(.Y(\instanceL2_prod_terms[1][3] [9]), .A0(
    instanceL2_n_10996), .A1(instanceL2_n_12191), .B0(
    \instanceL2_prod_terms[1][3] [10]));
  NAND2X1 instanceL2_g9861(.Y(instanceL2_n_12186), .A(instanceL2_n_12227), .B(
    instanceL2_n_12188));
  ADDFX1 instanceL2_g9862(.CO(instanceL2_n_12187), .S(
    \instanceL2_prod_terms[9][3] [7]), .A(layer1_out[34]), .B(layer1_out[31]),
     .CI(instanceL2_n_12190));
  NOR2X1 instanceL2_g9863(.Y(\instanceL2_prod_terms[1][3] [10]), .A(
    instanceL2_n_10996), .B(instanceL2_n_12191));
  AOI21X1 instanceL2_g9864(.Y(\instanceL2_prod_terms[2][3] [5]), .A0(
    layer1_out[32]), .A1(instanceL2_n_12194), .B0(instanceL2_n_12188));
  ADDFX1 instanceL2_g9865(.CO(instanceL2_n_12189), .S(
    \instanceL2_prod_terms[0][3][6] ), .A(instanceL2_n_11004), .B(
    instanceL2_n_12208), .CI(instanceL2_n_12193));
  NOR2X1 instanceL2_g9866(.Y(instanceL2_n_12188), .A(layer1_out[32]), .B(
    instanceL2_n_12194));
  OA21X1 instanceL2_g9867(.Y(\instanceL2_prod_terms[1][3] [8]), .A0(
    layer1_out[33]), .A1(instanceL2_n_12192), .B0(instanceL2_n_12191));
  ADDFX1 instanceL2_g9868(.CO(instanceL2_n_12190), .S(
    \instanceL2_prod_terms[9][3] [6]), .A(layer1_out[33]), .B(layer1_out[30]),
     .CI(instanceL2_n_12196));
  NAND2X1 instanceL2_g9869(.Y(instanceL2_n_12191), .A(layer1_out[33]), .B(
    instanceL2_n_12192));
  OAI21X1 instanceL2_g9870(.Y(instanceL2_n_12192), .A0(instanceL2_n_12222), .A1(
    instanceL2_n_12195), .B0(instanceL2_n_12224));
  OA21X1 instanceL2_g9871(.Y(\instanceL2_prod_terms[2][3] [4]), .A0(
    instanceL2_n_11001), .A1(instanceL2_n_12197), .B0(instanceL2_n_12194));
  CLKXOR2X1 instanceL2_g9872(.Y(\instanceL2_prod_terms[1][3] [7]), .A(
    instanceL2_n_12207), .B(instanceL2_n_12195));
  ADDFX1 instanceL2_g9873(.CO(instanceL2_n_12193), .S(
    \instanceL2_prod_terms[0][3][5] ), .A(instanceL2_n_10987), .B(
    instanceL2_n_12211), .CI(instanceL2_n_12198));
  NAND2X1 instanceL2_g9874(.Y(instanceL2_n_12194), .A(instanceL2_n_11001), .B(
    instanceL2_n_12197));
  ADDFX1 instanceL2_g9875(.CO(instanceL2_n_12196), .S(
    \instanceL2_prod_terms[9][3] [5]), .A(layer1_out[32]), .B(layer1_out[29]),
     .CI(instanceL2_n_12200));
  OA21X1 instanceL2_g9876(.Y(instanceL2_n_12195), .A0(instanceL2_n_12221), .A1(
    instanceL2_n_12199), .B0(instanceL2_n_12225));
  XOR2XL instanceL2_g9877(.Y(\instanceL2_prod_terms[1][3] [6]), .A(
    instanceL2_n_12208), .B(instanceL2_n_12199));
  AOI21X1 instanceL2_g9878(.Y(\instanceL2_prod_terms[2][3] [3]), .A0(
    layer1_out[30]), .A1(instanceL2_n_12203), .B0(instanceL2_n_12197));
  ADDFX1 instanceL2_g9879(.CO(instanceL2_n_12198), .S(
    \instanceL2_prod_terms[0][3][4] ), .A(instanceL2_n_11005), .B(
    instanceL2_n_12209), .CI(instanceL2_n_12205));
  NOR2X1 instanceL2_g9880(.Y(instanceL2_n_12197), .A(layer1_out[30]), .B(
    instanceL2_n_12203));
  XNOR2X1 instanceL2_g9881(.Y(\instanceL2_prod_terms[1][3] [5]), .A(
    instanceL2_n_12211), .B(instanceL2_n_12202));
  OA21X1 instanceL2_g9882(.Y(instanceL2_n_12199), .A0(instanceL2_n_12214), .A1(
    instanceL2_n_12201), .B0(instanceL2_n_12212));
  ADDFX1 instanceL2_g9883(.CO(instanceL2_n_12200), .S(
    \instanceL2_prod_terms[9][3] [4]), .A(layer1_out[31]), .B(layer1_out[28]),
     .CI(instanceL2_n_12220));
  XNOR2X1 instanceL2_g9884(.Y(\instanceL2_prod_terms[0][3][3] ), .A(
    instanceL2_n_12218), .B(instanceL2_n_12204));
  INVXL instanceL2_g9885(.Y(instanceL2_n_12201), .A(instanceL2_n_12202));
  OAI2BB1X1 instanceL2_g9886(.Y(instanceL2_n_12202), .A0N(instanceL2_n_12213),
     .A1N(instanceL2_n_12206), .B0(instanceL2_n_12216));
  OA21X1 instanceL2_g9887(.Y(\instanceL2_prod_terms[2][3] [2]), .A0(
    instanceL2_n_10992), .A1(instanceL2_n_12217), .B0(instanceL2_n_12203));
  XNOR2X1 instanceL2_g9888(.Y(\instanceL2_prod_terms[1][3] [4]), .A(
    instanceL2_n_12209), .B(instanceL2_n_12206));
  NAND2X1 instanceL2_g9889(.Y(instanceL2_n_12203), .A(instanceL2_n_10992), .B(
    instanceL2_n_12217));
  XNOR2X1 instanceL2_g9890(.Y(\instanceL2_prod_terms[1][3] [3]), .A(
    instanceL2_n_12219), .B(instanceL2_n_12210));
  MXI2XL instanceL2_g9891(.Y(instanceL2_n_12204), .A(instanceL2_n_10992), .B(
    layer1_out[29]), .S0(instanceL2_n_12210));
  AOI2BB1X1 instanceL2_g9892(.Y(instanceL2_n_12205), .A0N(layer1_out[29]), .A1N(
    instanceL2_n_12218), .B0(instanceL2_n_12210));
  AOI21X1 instanceL2_g9893(.Y(instanceL2_n_12206), .A0(instanceL2_n_12219), .A1(
    instanceL2_n_12223), .B0(instanceL2_n_12215));
  NAND2BX1 instanceL2_g9894(.Y(instanceL2_n_12207), .AN(instanceL2_n_12222), .B(
    instanceL2_n_12224));
  NAND2BX1 instanceL2_g9895(.Y(instanceL2_n_12208), .AN(instanceL2_n_12221), .B(
    instanceL2_n_12225));
  NAND2X1 instanceL2_g9896(.Y(instanceL2_n_12209), .A(instanceL2_n_12216), .B(
    instanceL2_n_12213));
  NOR2BX1 instanceL2_g9897(.Y(instanceL2_n_12210), .AN(instanceL2_n_12223), .B(
    instanceL2_n_12215));
  AOI2BB1X1 instanceL2_g9898(.Y(\instanceL2_prod_terms[9][3] [3]), .A0N(
    layer1_out[27]), .A1N(layer1_out[30]), .B0(instanceL2_n_12220));
  AOI21X1 instanceL2_g9899(.Y(\instanceL2_prod_terms[2][3] [1]), .A0(
    layer1_out[27]), .A1(layer1_out[28]), .B0(instanceL2_n_12217));
  NOR2BX1 instanceL2_g9900(.Y(\instanceL2_prod_terms[0][3][2] ), .AN(
    instanceL2_n_12219), .B(instanceL2_n_12218));
  NAND2BX1 instanceL2_g9901(.Y(instanceL2_n_12211), .AN(instanceL2_n_12214), .B(
    instanceL2_n_12212));
  NAND2XL instanceL2_g9902(.Y(instanceL2_n_12212), .A(layer1_out[32]), .B(
    layer1_out[30]));
  NAND2X1 instanceL2_g9903(.Y(instanceL2_n_12213), .A(instanceL2_n_10992), .B(
    instanceL2_n_11001));
  NOR2XL instanceL2_g9904(.Y(instanceL2_n_12214), .A(layer1_out[32]), .B(
    layer1_out[30]));
  NOR2X1 instanceL2_g9905(.Y(instanceL2_n_12215), .A(layer1_out[28]), .B(
    layer1_out[30]));
  NAND2X1 instanceL2_g9906(.Y(instanceL2_n_12216), .A(layer1_out[29]), .B(
    layer1_out[31]));
  NOR2X1 instanceL2_g9907(.Y(instanceL2_n_12217), .A(layer1_out[27]), .B(
    layer1_out[28]));
  NOR2XL instanceL2_g9908(.Y(instanceL2_n_12218), .A(layer1_out[29]), .B(
    layer1_out[27]));
  NAND2X1 instanceL2_g9909(.Y(instanceL2_n_12219), .A(layer1_out[27]), .B(
    layer1_out[29]));
  AND2XL instanceL2_g9910(.Y(instanceL2_n_12220), .A(layer1_out[30]), .B(
    layer1_out[27]));
  NOR2XL instanceL2_g9911(.Y(instanceL2_n_12221), .A(layer1_out[33]), .B(
    layer1_out[31]));
  NOR2XL instanceL2_g9912(.Y(instanceL2_n_12222), .A(layer1_out[34]), .B(
    layer1_out[32]));
  NAND2XL instanceL2_g9913(.Y(instanceL2_n_12223), .A(layer1_out[30]), .B(
    layer1_out[28]));
  NAND2XL instanceL2_g9914(.Y(instanceL2_n_12224), .A(layer1_out[34]), .B(
    layer1_out[32]));
  NAND2XL instanceL2_g9915(.Y(instanceL2_n_12225), .A(layer1_out[33]), .B(
    layer1_out[31]));
  NOR2X1 instanceL2_g9917(.Y(instanceL2_n_12226), .A(instanceL2_n_10996), .B(
    layer1_out[32]));
  NOR2X1 instanceL2_g9918(.Y(instanceL2_n_10987), .A(layer1_out[29]), .B(
    instanceL2_n_11001));
  NOR2X1 instanceL2_g9919(.Y(instanceL2_n_10988), .A(instanceL2_n_12227), .B(
    layer1_out[31]));
  INVX1 instanceL2_g9921(.Y(instanceL2_n_10992), .A(layer1_out[29]));
  INVX1 instanceL2_g9923(.Y(instanceL2_n_10996), .A(layer1_out[34]));
  INVX1 instanceL2_g9925(.Y(instanceL2_n_11001), .A(layer1_out[31]));
  INVX1 instanceL2_g9926(.Y(instanceL2_n_12227), .A(layer1_out[33]));
  NOR2BX1 instanceL2_g11211(.Y(instanceL2_n_11004), .AN(layer1_out[32]), .B(
    layer1_out[30]));
  NOR2BX1 instanceL2_g9927(.Y(instanceL2_n_11005), .AN(layer1_out[30]), .B(
    layer1_out[28]));
  AOI2BB1X1 instanceL2_g11212(.Y(\instanceL2_prod_terms[6][1] [10]), .A0N(
    layer1_out[16]), .A1N(instanceL2_n_12228), .B0(
    \instanceL2_prod_terms[6][1] [11]));
  AND2X1 instanceL2_g9916(.Y(\instanceL2_prod_terms[6][1] [11]), .A(
    instanceL2_n_12228), .B(layer1_out[16]));
  AOI21X1 instanceL2_g11213(.Y(\instanceL2_prod_terms[6][1] [9]), .A0(
    instanceL2_n_12276), .A1(instanceL2_n_11019), .B0(instanceL2_n_12228));
  NOR2X1 instanceL2_g11214(.Y(instanceL2_n_12228), .A(instanceL2_n_12276), .B(
    instanceL2_n_11019));
  XNOR2X1 instanceL2_g11215(.Y(\instanceL2_prod_terms[1][1][8] ), .A(
    instanceL2_n_12236), .B(instanceL2_n_12229));
  OA21X1 instanceL2_g9920(.Y(\instanceL2_prod_terms[6][1] [8]), .A0(
    layer1_out[14]), .A1(instanceL2_n_11025), .B0(instanceL2_n_11019));
  NAND2X1 instanceL2_g11216(.Y(instanceL2_n_11019), .A(layer1_out[14]), .B(
    instanceL2_n_11025));
  XNOR2X1 instanceL2_g9922(.Y(\instanceL2_prod_terms[1][1][7] ), .A(
    instanceL2_n_11079), .B(instanceL2_n_11027));
  OAI21X1 instanceL2_g11217(.Y(instanceL2_n_12229), .A0(instanceL2_n_12266), .A1(
    instanceL2_n_11027), .B0(instanceL2_n_11121));
  ADDFX1 instanceL2_g9924(.CO(instanceL2_n_11025), .S(
    \instanceL2_prod_terms[6][1] [7]), .A(layer1_out[16]), .B(layer1_out[13]),
     .CI(instanceL2_n_12230));
  ADDFX1 instanceL2_g11218(.CO(instanceL2_n_11027), .S(
    \instanceL2_prod_terms[1][1][6] ), .A(instanceL2_n_12268), .B(
    instanceL2_n_11135), .CI(instanceL2_n_11033));
  OR2XL instanceL2_g11219(.Y(\instanceL2_prod_terms[1][1][9] ), .A(
    instanceL2_n_12233), .B(instanceL2_n_11036));
  ADDFX1 instanceL2_g11220(.CO(instanceL2_n_12230), .S(
    \instanceL2_prod_terms[6][1] [6]), .A(layer1_out[15]), .B(layer1_out[12]),
     .CI(instanceL2_n_11044));
  ADDFX1 instanceL2_g9928(.CO(instanceL2_n_11033), .S(
    \instanceL2_prod_terms[1][1][5] ), .A(instanceL2_n_12265), .B(
    instanceL2_n_12252), .CI(instanceL2_n_11049));
  AO21X1 instanceL2_g9929(.Y(\instanceL2_prod_terms[0][1][8] ), .A0(
    instanceL2_n_12275), .A1(instanceL2_n_12231), .B0(instanceL2_n_11036));
  NOR2X1 instanceL2_g9930(.Y(instanceL2_n_11036), .A(instanceL2_n_12275), .B(
    instanceL2_n_12231));
  OAI2BB1X1 instanceL2_g9931(.Y(\instanceL2_prod_terms[9][1] [10]), .A0N(
    layer1_out[16]), .A1N(instanceL2_n_12232), .B0(instanceL2_n_12255));
  XNOR2X1 instanceL2_g9932(.Y(\instanceL2_prod_terms[9][1] [8]), .A(
    instanceL2_n_12247), .B(instanceL2_n_12232));
  ADDFX1 instanceL2_g9933(.CO(instanceL2_n_11044), .S(
    \instanceL2_prod_terms[6][1] [5]), .A(layer1_out[14]), .B(layer1_out[11]),
     .CI(instanceL2_n_11066));
  OAI211X1 instanceL2_g9934(.Y(instanceL2_n_12231), .A0(instanceL2_n_11112), .A1(
    instanceL2_n_11056), .B0(instanceL2_n_12262), .C0(instanceL2_n_12255));
  XNOR2X1 instanceL2_g9935(.Y(\instanceL2_prod_terms[9][1] [7]), .A(
    instanceL2_n_12250), .B(instanceL2_n_11056));
  ADDFX1 instanceL2_g9936(.CO(instanceL2_n_11049), .S(
    \instanceL2_prod_terms[1][1][4] ), .A(instanceL2_n_12269), .B(
    instanceL2_n_12251), .CI(instanceL2_n_12240));
  AO21X1 instanceL2_g9937(.Y(\instanceL2_prod_terms[2][1] [7]), .A0(
    layer1_out[16]), .A1(instanceL2_n_12239), .B0(instanceL2_n_12233));
  XNOR2X1 instanceL2_g9938(.Y(\instanceL2_prod_terms[9][1] [6]), .A(
    instanceL2_n_12248), .B(instanceL2_n_12235));
  OAI211X1 instanceL2_g9939(.Y(instanceL2_n_12232), .A0(instanceL2_n_12278), .A1(
    instanceL2_n_12234), .B0(instanceL2_n_12256), .C0(instanceL2_n_12262));
  NOR2XL instanceL2_g9940(.Y(instanceL2_n_12233), .A(layer1_out[16]), .B(
    instanceL2_n_12239));
  AOI31X1 instanceL2_g9941(.Y(instanceL2_n_11056), .A0(instanceL2_n_11141), .A1(
    instanceL2_n_12259), .A2(instanceL2_n_12237), .B0(instanceL2_n_12245));
  XNOR2X1 instanceL2_g9942(.Y(\instanceL2_prod_terms[2][1] [5]), .A(
    layer1_out[14]), .B(instanceL2_n_12241));
  XNOR2X1 instanceL2_g9943(.Y(\instanceL2_prod_terms[1][1][3] ), .A(
    instanceL2_n_12260), .B(instanceL2_n_11074));
  XNOR2X1 instanceL2_g9944(.Y(\instanceL2_prod_terms[0][1][4] ), .A(
    instanceL2_n_12246), .B(instanceL2_n_12237));
  INVX1 instanceL2_g9945(.Y(instanceL2_n_12234), .A(instanceL2_n_12235));
  ADDFX1 instanceL2_g9946(.CO(instanceL2_n_11066), .S(
    \instanceL2_prod_terms[6][1] [4]), .A(layer1_out[13]), .B(layer1_out[10]),
     .CI(instanceL2_n_12258));
  OAI211X1 instanceL2_g9947(.Y(instanceL2_n_12235), .A0(instanceL2_n_12244), .A1(
    instanceL2_n_12238), .B0(instanceL2_n_12264), .C0(instanceL2_n_11150));
  XNOR2X1 instanceL2_g9948(.Y(\instanceL2_prod_terms[9][1] [4]), .A(
    instanceL2_n_11128), .B(instanceL2_n_12238));
  MXI2XL instanceL2_g9949(.Y(\instanceL2_prod_terms[2][1] [3]), .A(
    instanceL2_n_12273), .B(layer1_out[12]), .S0(instanceL2_n_12243));
  XNOR2X1 instanceL2_g9950(.Y(\instanceL2_prod_terms[2][1] [6]), .A(
    layer1_out[15]), .B(instanceL2_n_11098));
  XNOR2X1 instanceL2_g9951(.Y(instanceL2_n_11074), .A(layer1_out[11]), .B(
    instanceL2_n_12279));
  MXI2XL instanceL2_g9952(.Y(instanceL2_n_12236), .A(instanceL2_n_12276), .B(
    layer1_out[15]), .S0(instanceL2_n_12270));
  CLKXOR2X1 instanceL2_g9953(.Y(\instanceL2_prod_terms[9][1] [3]), .A(
    instanceL2_n_12257), .B(instanceL2_n_12249));
  XNOR2X1 instanceL2_g9954(.Y(instanceL2_n_11079), .A(instanceL2_n_12266), .B(
    instanceL2_n_11121));
  OAI211X1 instanceL2_g9955(.Y(instanceL2_n_12237), .A0(instanceL2_n_12257), .A1(
    instanceL2_n_12267), .B0(instanceL2_n_12253), .C0(instanceL2_n_12264));
  NAND2X1 instanceL2_g9956(.Y(\instanceL2_prod_terms[2][1] [13]), .A(
    instanceL2_n_12254), .B(instanceL2_n_11098));
  NAND2BX1 instanceL2_g9957(.Y(instanceL2_n_12238), .AN(instanceL2_n_12260), .B(
    layer1_out[10]));
  AOI21X1 instanceL2_g9958(.Y(\instanceL2_prod_terms[2][1] [4]), .A0(
    layer1_out[13]), .A1(instanceL2_n_12242), .B0(instanceL2_n_12241));
  AND2XL instanceL2_g9959(.Y(instanceL2_n_12239), .A(instanceL2_n_12276), .B(
    instanceL2_n_11098));
  OA21X1 instanceL2_g9960(.Y(instanceL2_n_12240), .A0(instanceL2_n_12274), .A1(
    layer1_out[11]), .B0(instanceL2_n_12279));
  NOR2X1 instanceL2_g9961(.Y(instanceL2_n_11098), .A(instanceL2_n_12259), .B(
    instanceL2_n_12242));
  OA21X1 instanceL2_g9962(.Y(\instanceL2_prod_terms[2][1] [2]), .A0(
    instanceL2_n_12272), .A1(instanceL2_n_12261), .B0(instanceL2_n_12243));
  NOR2X1 instanceL2_g9963(.Y(instanceL2_n_12241), .A(layer1_out[13]), .B(
    instanceL2_n_12242));
  NOR2BX1 instanceL2_g9964(.Y(\instanceL2_prod_terms[2][1] [1]), .AN(
    instanceL2_n_12257), .B(instanceL2_n_12261));
  NAND2BX1 instanceL2_g9966(.Y(instanceL2_n_12244), .AN(instanceL2_n_12267), .B(
    instanceL2_n_11141));
  OR2XL instanceL2_g9967(.Y(instanceL2_n_11112), .A(instanceL2_n_12263), .B(
    instanceL2_n_12254));
  NAND2XL instanceL2_g9968(.Y(instanceL2_n_12245), .A(instanceL2_n_11150), .B(
    instanceL2_n_12256));
  NAND2XL instanceL2_g9969(.Y(instanceL2_n_12246), .A(instanceL2_n_11150), .B(
    instanceL2_n_11141));
  NAND2BXL instanceL2_g9970(.Y(instanceL2_n_12247), .AN(instanceL2_n_12254), .B(
    instanceL2_n_12255));
  NAND2XL instanceL2_g9971(.Y(instanceL2_n_12248), .A(instanceL2_n_12256), .B(
    instanceL2_n_12259));
  NAND2X1 instanceL2_g9972(.Y(instanceL2_n_12242), .A(instanceL2_n_12267), .B(
    instanceL2_n_12261));
  NAND2X1 instanceL2_g9973(.Y(instanceL2_n_12243), .A(instanceL2_n_12272), .B(
    instanceL2_n_12261));
  AOI21X1 instanceL2_g9974(.Y(\instanceL2_prod_terms[6][1] [3]), .A0(
    instanceL2_n_12274), .A1(instanceL2_n_12273), .B0(instanceL2_n_12258));
  AOI21X1 instanceL2_g9975(.Y(\instanceL2_prod_terms[1][1][2] ), .A0(
    layer1_out[9]), .A1(layer1_out[11]), .B0(instanceL2_n_12260));
  NOR2BX1 instanceL2_g9976(.Y(instanceL2_n_11128), .AN(instanceL2_n_12264), .B(
    instanceL2_n_12267));
  OAI21XL instanceL2_g9977(.Y(instanceL2_n_12249), .A0(layer1_out[10]), .A1(
    layer1_out[11]), .B0(instanceL2_n_12253));
  NOR2BX1 instanceL2_g9978(.Y(instanceL2_n_12250), .AN(instanceL2_n_12262), .B(
    instanceL2_n_12263));
  AOI21X1 instanceL2_g9979(.Y(instanceL2_n_12251), .A0(instanceL2_n_12271), .A1(
    layer1_out[11]), .B0(instanceL2_n_12265));
  AOI21X1 instanceL2_g9980(.Y(instanceL2_n_11135), .A0(instanceL2_n_12276), .A1(
    layer1_out[13]), .B0(instanceL2_n_12266));
  OAI22X1 instanceL2_g9981(.Y(instanceL2_n_12252), .A0(layer1_out[14]), .A1(
    layer1_out[12]), .B0(instanceL2_n_12277), .B1(instanceL2_n_12273));
  OAI22X1 instanceL2_g9982(.Y(instanceL2_n_11121), .A0(layer1_out[16]), .A1(
    layer1_out[14]), .B0(instanceL2_n_12275), .B1(instanceL2_n_12277));
  NAND2XL instanceL2_g9984(.Y(instanceL2_n_12253), .A(layer1_out[11]), .B(
    layer1_out[10]));
  NOR2XL instanceL2_g9985(.Y(instanceL2_n_12254), .A(layer1_out[16]), .B(
    layer1_out[15]));
  NAND2X1 instanceL2_g9986(.Y(instanceL2_n_12255), .A(layer1_out[15]), .B(
    layer1_out[16]));
  NAND2X1 instanceL2_g9987(.Y(instanceL2_n_11141), .A(instanceL2_n_12271), .B(
    instanceL2_n_12273));
  NAND2X1 instanceL2_g9988(.Y(instanceL2_n_12256), .A(layer1_out[13]), .B(
    layer1_out[14]));
  NAND2XL instanceL2_g9989(.Y(instanceL2_n_12257), .A(layer1_out[9]), .B(
    layer1_out[10]));
  NOR2X1 instanceL2_g9990(.Y(instanceL2_n_12258), .A(instanceL2_n_12274), .B(
    instanceL2_n_12273));
  NAND2X1 instanceL2_g9991(.Y(instanceL2_n_12259), .A(instanceL2_n_12271), .B(
    instanceL2_n_12277));
  NOR2X1 instanceL2_g9992(.Y(instanceL2_n_12260), .A(layer1_out[9]), .B(
    layer1_out[11]));
  NOR2X1 instanceL2_g9993(.Y(instanceL2_n_12261), .A(layer1_out[9]), .B(
    layer1_out[10]));
  NOR2X1 instanceL2_g9995(.Y(instanceL2_n_12268), .A(instanceL2_n_12277), .B(
    layer1_out[12]));
  NOR2X1 instanceL2_g9996(.Y(instanceL2_n_12269), .A(layer1_out[10]), .B(
    instanceL2_n_12273));
  NAND2X1 instanceL2_g9997(.Y(instanceL2_n_12270), .A(layer1_out[16]), .B(
    instanceL2_n_12277));
  NAND2X1 instanceL2_g9998(.Y(instanceL2_n_11150), .A(layer1_out[12]), .B(
    layer1_out[13]));
  NAND2XL instanceL2_g9999(.Y(instanceL2_n_12262), .A(layer1_out[15]), .B(
    layer1_out[14]));
  NOR2XL instanceL2_g10000(.Y(instanceL2_n_12263), .A(layer1_out[15]), .B(
    layer1_out[14]));
  NAND2X1 instanceL2_g10001(.Y(instanceL2_n_12264), .A(layer1_out[11]), .B(
    layer1_out[12]));
  NOR2X1 instanceL2_g10002(.Y(instanceL2_n_12265), .A(layer1_out[11]), .B(
    instanceL2_n_12271));
  NOR2X1 instanceL2_g10003(.Y(instanceL2_n_12266), .A(instanceL2_n_12276), .B(
    layer1_out[13]));
  NOR2X1 instanceL2_g10004(.Y(instanceL2_n_12267), .A(layer1_out[11]), .B(
    layer1_out[12]));
  INVX1 instanceL2_g10006(.Y(instanceL2_n_12271), .A(layer1_out[13]));
  INVX1 instanceL2_g10007(.Y(instanceL2_n_12272), .A(layer1_out[11]));
  INVX1 instanceL2_g10008(.Y(instanceL2_n_12273), .A(layer1_out[12]));
  INVX1 instanceL2_g10009(.Y(instanceL2_n_12274), .A(layer1_out[9]));
  INVX1 instanceL2_g10010(.Y(instanceL2_n_12275), .A(layer1_out[16]));
  INVX1 instanceL2_g10011(.Y(instanceL2_n_12276), .A(layer1_out[15]));
  INVX1 instanceL2_g10012(.Y(instanceL2_n_12277), .A(layer1_out[14]));
  NAND2BX1 instanceL2_g11221(.Y(instanceL2_n_12278), .AN(instanceL2_n_12263), .B(
    instanceL2_n_12259));
  MXI2XL instanceL2_g11222(.Y(instanceL2_n_12279), .A(layer1_out[12]), .B(
    instanceL2_n_12273), .S0(layer1_out[10]));
  AOI21X1 instanceL2_g9434(.Y(\instanceL2_prod_terms[1][10][9] ), .A0(
    instanceL2_n_10763), .A1(instanceL2_n_10704), .B0(
    \instanceL2_prod_terms[1][10][10] ));
  NOR2X1 instanceL2_g9435(.Y(\instanceL2_prod_terms[1][10][10] ), .A(
    instanceL2_n_10763), .B(instanceL2_n_10704));
  AOI21X1 instanceL2_g9436(.Y(\instanceL2_prod_terms[0][10][8] ), .A0(
    layer1_out[97]), .A1(instanceL2_n_10711), .B0(instanceL2_n_10701));
  OA21X1 instanceL2_g9437(.Y(\instanceL2_prod_terms[1][10][8] ), .A0(
    layer1_out[96]), .A1(instanceL2_n_10708), .B0(instanceL2_n_10704));
  INVX1 instanceL2_g9438(.Y(\instanceL2_prod_terms[0][10][13] ), .A(
    instanceL2_n_10701));
  NOR2X1 instanceL2_g9439(.Y(instanceL2_n_10701), .A(layer1_out[97]), .B(
    instanceL2_n_10711));
  NAND2X1 instanceL2_g9440(.Y(instanceL2_n_10704), .A(layer1_out[96]), .B(
    instanceL2_n_10708));
  ADDFX1 instanceL2_g9441(.CO(instanceL2_n_10708), .S(
    \instanceL2_prod_terms[1][10][7] ), .A(layer1_out[97]), .B(layer1_out[95]),
     .CI(instanceL2_n_10716));
  OA21X1 instanceL2_g9442(.Y(\instanceL2_prod_terms[0][10][7] ), .A0(
    instanceL2_n_10755), .A1(instanceL2_n_10719), .B0(instanceL2_n_10711));
  NAND2X1 instanceL2_g9443(.Y(instanceL2_n_10711), .A(instanceL2_n_10755), .B(
    instanceL2_n_10719));
  ADDFX1 instanceL2_g9444(.CO(instanceL2_n_10716), .S(
    \instanceL2_prod_terms[1][10][6] ), .A(layer1_out[96]), .B(layer1_out[94]),
     .CI(instanceL2_n_10723));
  AOI21X1 instanceL2_g9445(.Y(\instanceL2_prod_terms[0][10][6] ), .A0(
    layer1_out[95]), .A1(instanceL2_n_10725), .B0(instanceL2_n_10719));
  NOR2X1 instanceL2_g9446(.Y(instanceL2_n_10719), .A(layer1_out[95]), .B(
    instanceL2_n_10725));
  ADDFX1 instanceL2_g9447(.CO(instanceL2_n_10723), .S(
    \instanceL2_prod_terms[1][10][5] ), .A(layer1_out[93]), .B(layer1_out[95]),
     .CI(instanceL2_n_10730));
  OA21X1 instanceL2_g9448(.Y(\instanceL2_prod_terms[0][10][5] ), .A0(
    instanceL2_n_10757), .A1(instanceL2_n_10734), .B0(instanceL2_n_10725));
  NAND2X1 instanceL2_g9449(.Y(instanceL2_n_10725), .A(instanceL2_n_10757), .B(
    instanceL2_n_10734));
  ADDFX1 instanceL2_g9450(.CO(instanceL2_n_10730), .S(
    \instanceL2_prod_terms[1][10][4] ), .A(layer1_out[92]), .B(layer1_out[94]),
     .CI(instanceL2_n_10738));
  AOI21X1 instanceL2_g9451(.Y(\instanceL2_prod_terms[0][10][4] ), .A0(
    layer1_out[93]), .A1(instanceL2_n_10740), .B0(instanceL2_n_10734));
  NOR2X1 instanceL2_g9452(.Y(instanceL2_n_10734), .A(layer1_out[93]), .B(
    instanceL2_n_10740));
  ADDFX1 instanceL2_g9453(.CO(instanceL2_n_10738), .S(
    \instanceL2_prod_terms[1][10][3] ), .A(layer1_out[93]), .B(layer1_out[91]),
     .CI(instanceL2_n_10751));
  OA21X1 instanceL2_g9454(.Y(\instanceL2_prod_terms[0][10][3] ), .A0(
    instanceL2_n_10753), .A1(instanceL2_n_10750), .B0(instanceL2_n_10740));
  NAND2X1 instanceL2_g9455(.Y(instanceL2_n_10740), .A(instanceL2_n_10753), .B(
    instanceL2_n_10750));
  AOI21X1 instanceL2_g9456(.Y(\instanceL2_prod_terms[0][10][2] ), .A0(
    layer1_out[91]), .A1(layer1_out[90]), .B0(instanceL2_n_10750));
  AOI2BB1X1 instanceL2_g9457(.Y(\instanceL2_prod_terms[1][10][2] ), .A0N(
    layer1_out[92]), .A1N(layer1_out[90]), .B0(instanceL2_n_10751));
  NOR2X1 instanceL2_g9458(.Y(instanceL2_n_10750), .A(layer1_out[90]), .B(
    layer1_out[91]));
  AND2XL instanceL2_g9459(.Y(instanceL2_n_10751), .A(layer1_out[92]), .B(
    layer1_out[90]));
  INVX1 instanceL2_g9460(.Y(instanceL2_n_10753), .A(layer1_out[92]));
  INVX1 instanceL2_g9461(.Y(instanceL2_n_10755), .A(layer1_out[96]));
  INVX1 instanceL2_g9462(.Y(instanceL2_n_10757), .A(layer1_out[94]));
  INVX1 instanceL2_g9463(.Y(instanceL2_n_10763), .A(layer1_out[97]));
  XNOR2X1 instanceL2_g9745(.Y(\instanceL2_prod_terms[2][8][10] ), .A(
    layer1_out[80]), .B(instanceL2_n_12280));
  OA21X1 instanceL2_g9746(.Y(\instanceL2_prod_terms[1][8][9] ), .A0(
    instanceL2_n_12336), .A1(instanceL2_n_12284), .B0(
    \instanceL2_prod_terms[1][8][13] ));
  MX2X1 instanceL2_g9747(.Y(\instanceL2_prod_terms[2][8][9] ), .A(layer1_out[79]),
     .B(instanceL2_n_10991), .S0(instanceL2_n_12281));
  NAND2X1 instanceL2_g9748(.Y(\instanceL2_prod_terms[1][8][13] ), .A(
    instanceL2_n_12336), .B(instanceL2_n_12284));
  OA22X1 instanceL2_g9749(.Y(instanceL2_n_12280), .A0(instanceL2_n_10991), .A1(
    instanceL2_n_12282), .B0(instanceL2_n_12333), .B1(instanceL2_n_12303));
  OAI2BB1X1 instanceL2_g9750(.Y(instanceL2_n_12281), .A0N(layer1_out[80]), .A1N(
    layer1_out[78]), .B0(instanceL2_n_12282));
  AOI2BB1X1 instanceL2_g9751(.Y(\instanceL2_prod_terms[2][8][11] ), .A0N(
    layer1_out[78]), .A1N(instanceL2_n_12283), .B0(instanceL2_n_12303));
  XNOR2X1 instanceL2_g9752(.Y(\instanceL2_prod_terms[2][8][8] ), .A(
    instanceL2_n_12313), .B(instanceL2_n_12283));
  AOI21X1 instanceL2_g9753(.Y(\instanceL2_prod_terms[1][8][8] ), .A0(
    layer1_out[79]), .A1(instanceL2_n_12286), .B0(instanceL2_n_12284));
  OAI2BB1X1 instanceL2_g9754(.Y(instanceL2_n_12282), .A0N(instanceL2_n_12336),
     .A1N(instanceL2_n_12333), .B0(instanceL2_n_12283));
  ADDFX1 instanceL2_g9755(.CO(instanceL2_n_12283), .S(
    \instanceL2_prod_terms[2][8][7] ), .A(layer1_out[79]), .B(layer1_out[77]),
     .CI(instanceL2_n_12285));
  NOR2X1 instanceL2_g9756(.Y(instanceL2_n_12284), .A(layer1_out[79]), .B(
    instanceL2_n_12286));
  OA21X1 instanceL2_g9757(.Y(\instanceL2_prod_terms[1][8][7] ), .A0(
    instanceL2_n_12333), .A1(instanceL2_n_12287), .B0(instanceL2_n_12286));
  ADDFX1 instanceL2_g9758(.CO(instanceL2_n_12285), .S(
    \instanceL2_prod_terms[2][8][6] ), .A(layer1_out[78]), .B(layer1_out[76]),
     .CI(instanceL2_n_12288));
  NAND2X1 instanceL2_g9759(.Y(instanceL2_n_12286), .A(instanceL2_n_12333), .B(
    instanceL2_n_12287));
  XNOR2X1 instanceL2_g9760(.Y(\instanceL2_prod_terms[1][8][6] ), .A(
    layer1_out[77]), .B(instanceL2_n_12293));
  OAI2BB1X1 instanceL2_g9761(.Y(\instanceL2_prod_terms[6][8] [10]), .A0N(
    layer1_out[80]), .A1N(instanceL2_n_12290), .B0(instanceL2_n_12303));
  NOR2BX1 instanceL2_g9762(.Y(instanceL2_n_12287), .AN(instanceL2_n_12293), .B(
    layer1_out[77]));
  OAI2BB1X1 instanceL2_g9763(.Y(instanceL2_n_12288), .A0N(instanceL2_n_12328),
     .A1N(instanceL2_n_12289), .B0(instanceL2_n_12317));
  XNOR2X1 instanceL2_g9764(.Y(\instanceL2_prod_terms[6][8] [8]), .A(
    instanceL2_n_12311), .B(instanceL2_n_12290));
  OAI33X1 instanceL2_g9765(.Y(\instanceL2_prod_terms[6][8] [9]), .A0(
    instanceL2_n_12336), .A1(instanceL2_n_12321), .A2(instanceL2_n_12290), .B0(
    instanceL2_n_10991), .B1(layer1_out[80]), .B2(instanceL2_n_12291));
  XNOR2X1 instanceL2_g9766(.Y(\instanceL2_prod_terms[2][8][5] ), .A(
    instanceL2_n_12306), .B(instanceL2_n_12289));
  XNOR2X1 instanceL2_g9767(.Y(\instanceL2_prod_terms[6][8] [7]), .A(
    instanceL2_n_12307), .B(instanceL2_n_12292));
  ADDFX1 instanceL2_g9768(.CO(instanceL2_n_12289), .S(
    \instanceL2_prod_terms[2][8][4] ), .A(layer1_out[76]), .B(layer1_out[74]),
     .CI(instanceL2_n_12295));
  AOI21X1 instanceL2_g9769(.Y(\instanceL2_prod_terms[1][8][5] ), .A0(
    layer1_out[76]), .A1(instanceL2_n_12299), .B0(instanceL2_n_12293));
  INVX1 instanceL2_g9770(.Y(instanceL2_n_12291), .A(instanceL2_n_12290));
  OAI211X1 instanceL2_g9771(.Y(instanceL2_n_12290), .A0(instanceL2_n_12325), .A1(
    instanceL2_n_12294), .B0(instanceL2_n_12318), .C0(instanceL2_n_12315));
  NAND2X1 instanceL2_g9772(.Y(instanceL2_n_12292), .A(instanceL2_n_12318), .B(
    instanceL2_n_12294));
  XNOR2X1 instanceL2_g9773(.Y(\instanceL2_prod_terms[6][8] [6]), .A(
    instanceL2_n_12309), .B(instanceL2_n_12298));
  NOR2X1 instanceL2_g9774(.Y(instanceL2_n_12293), .A(layer1_out[76]), .B(
    instanceL2_n_12299));
  NAND2BX1 instanceL2_g9775(.Y(instanceL2_n_12294), .AN(instanceL2_n_12316), .B(
    instanceL2_n_12298));
  CLKXOR2X1 instanceL2_g9776(.Y(\instanceL2_prod_terms[6][8] [5]), .A(
    instanceL2_n_12312), .B(instanceL2_n_12301));
  INVX1 instanceL2_g9777(.Y(\instanceL2_prod_terms[2][8][3] ), .A(
    instanceL2_n_12296));
  INVX1 instanceL2_g9778(.Y(instanceL2_n_12295), .A(instanceL2_n_12297));
  ADDFX1 instanceL2_g9779(.CO(instanceL2_n_12297), .S(instanceL2_n_12296), .A(
    instanceL2_n_12331), .B(instanceL2_n_12334), .CI(instanceL2_n_12320));
  AOI21X1 instanceL2_g9780(.Y(\instanceL2_prod_terms[1][8][4] ), .A0(
    layer1_out[75]), .A1(instanceL2_n_12310), .B0(instanceL2_n_12300));
  OAI22X1 instanceL2_g9781(.Y(instanceL2_n_12298), .A0(instanceL2_n_12322), .A1(
    instanceL2_n_12302), .B0(instanceL2_n_12332), .B1(instanceL2_n_12329));
  INVX1 instanceL2_g9782(.Y(instanceL2_n_12299), .A(instanceL2_n_12300));
  NOR2X1 instanceL2_g9783(.Y(instanceL2_n_12300), .A(layer1_out[75]), .B(
    instanceL2_n_12310));
  XNOR2X1 instanceL2_g9784(.Y(\instanceL2_prod_terms[6][8] [4]), .A(
    instanceL2_n_12314), .B(instanceL2_n_12304));
  OAI2BB1X1 instanceL2_g9785(.Y(instanceL2_n_12301), .A0N(layer1_out[76]), .A1N(
    layer1_out[75]), .B0(instanceL2_n_12302));
  OAI2BB1X1 instanceL2_g9786(.Y(instanceL2_n_12302), .A0N(instanceL2_n_12332),
     .A1N(instanceL2_n_12331), .B0(instanceL2_n_12304));
  OAI22X1 instanceL2_g9787(.Y(\instanceL2_prod_terms[6][8] [2]), .A0(
    instanceL2_n_12330), .A1(instanceL2_n_12305), .B0(instanceL2_n_12319), .B1(
    instanceL2_n_12327));
  XNOR2X1 instanceL2_g9788(.Y(\instanceL2_prod_terms[6][8] [3]), .A(
    instanceL2_n_12305), .B(instanceL2_n_12308));
  INVX1 instanceL2_g9789(.Y(instanceL2_n_12303), .A(instanceL2_n_12321));
  OA21X1 instanceL2_g9790(.Y(\instanceL2_prod_terms[1][8][3] ), .A0(
    instanceL2_n_12335), .A1(instanceL2_n_12326), .B0(instanceL2_n_12310));
  OAI211X1 instanceL2_g9791(.Y(instanceL2_n_12304), .A0(instanceL2_n_12319), .A1(
    instanceL2_n_12323), .B0(instanceL2_n_12327), .C0(instanceL2_n_12324));
  NOR2BX1 instanceL2_g9792(.Y(\instanceL2_prod_terms[1][8][2] ), .AN(
    instanceL2_n_12319), .B(instanceL2_n_12326));
  NAND2XL instanceL2_g9793(.Y(instanceL2_n_12306), .A(instanceL2_n_12317), .B(
    instanceL2_n_12328));
  NAND2BXL instanceL2_g9794(.Y(instanceL2_n_12307), .AN(instanceL2_n_12325), .B(
    instanceL2_n_12315));
  NAND2BX1 instanceL2_g9795(.Y(instanceL2_n_12308), .AN(instanceL2_n_12323), .B(
    instanceL2_n_12324));
  NAND2BX1 instanceL2_g9796(.Y(instanceL2_n_12309), .AN(instanceL2_n_12316), .B(
    instanceL2_n_12318));
  NAND2X1 instanceL2_g9797(.Y(instanceL2_n_12305), .A(instanceL2_n_12319), .B(
    instanceL2_n_12327));
  OA21X1 instanceL2_g9798(.Y(\instanceL2_prod_terms[2][8][2] ), .A0(
    layer1_out[74]), .A1(layer1_out[72]), .B0(instanceL2_n_12320));
  OAI2BB1X1 instanceL2_g9799(.Y(instanceL2_n_12311), .A0N(instanceL2_n_12336),
     .A1N(instanceL2_n_10991), .B0(instanceL2_n_12303));
  AOI21XL instanceL2_g9800(.Y(instanceL2_n_12312), .A0(layer1_out[77]), .A1(
    layer1_out[76]), .B0(instanceL2_n_12322));
  OAI22X1 instanceL2_g9801(.Y(instanceL2_n_12313), .A0(layer1_out[80]), .A1(
    layer1_out[78]), .B0(instanceL2_n_12336), .B1(instanceL2_n_12333));
  OAI22X1 instanceL2_g9802(.Y(instanceL2_n_12314), .A0(layer1_out[76]), .A1(
    layer1_out[75]), .B0(instanceL2_n_12332), .B1(instanceL2_n_12331));
  NAND2X1 instanceL2_g9803(.Y(instanceL2_n_12310), .A(instanceL2_n_12335), .B(
    instanceL2_n_12326));
  NAND2X1 instanceL2_g9805(.Y(instanceL2_n_12315), .A(layer1_out[79]), .B(
    layer1_out[78]));
  NOR2XL instanceL2_g9806(.Y(instanceL2_n_12316), .A(layer1_out[78]), .B(
    layer1_out[77]));
  NAND2XL instanceL2_g9807(.Y(instanceL2_n_12317), .A(layer1_out[77]), .B(
    layer1_out[75]));
  NAND2X1 instanceL2_g9808(.Y(instanceL2_n_12318), .A(layer1_out[78]), .B(
    layer1_out[77]));
  NAND2X1 instanceL2_g9809(.Y(instanceL2_n_12319), .A(layer1_out[72]), .B(
    layer1_out[73]));
  NAND2X1 instanceL2_g9810(.Y(instanceL2_n_12320), .A(layer1_out[72]), .B(
    layer1_out[74]));
  NOR2X1 instanceL2_g9811(.Y(instanceL2_n_12321), .A(instanceL2_n_12336), .B(
    instanceL2_n_10991));
  INVX1 instanceL2_g9812(.Y(instanceL2_n_12328), .A(instanceL2_n_12329));
  NOR2XL instanceL2_g9813(.Y(instanceL2_n_12330), .A(layer1_out[74]), .B(
    layer1_out[73]));
  NOR2X1 instanceL2_g9814(.Y(instanceL2_n_12322), .A(layer1_out[77]), .B(
    layer1_out[76]));
  NOR2X1 instanceL2_g9815(.Y(instanceL2_n_12323), .A(layer1_out[74]), .B(
    layer1_out[75]));
  NAND2XL instanceL2_g9816(.Y(instanceL2_n_12324), .A(layer1_out[74]), .B(
    layer1_out[75]));
  NOR2X1 instanceL2_g9817(.Y(instanceL2_n_12325), .A(layer1_out[79]), .B(
    layer1_out[78]));
  NOR2X1 instanceL2_g9818(.Y(instanceL2_n_12326), .A(layer1_out[72]), .B(
    layer1_out[73]));
  NAND2XL instanceL2_g9819(.Y(instanceL2_n_12327), .A(layer1_out[73]), .B(
    layer1_out[74]));
  NOR2X1 instanceL2_g9820(.Y(instanceL2_n_12329), .A(layer1_out[77]), .B(
    layer1_out[75]));
  INVX1 instanceL2_g9821(.Y(instanceL2_n_12331), .A(layer1_out[75]));
  INVX1 instanceL2_g9822(.Y(instanceL2_n_12332), .A(layer1_out[76]));
  INVX1 instanceL2_g9823(.Y(instanceL2_n_12333), .A(layer1_out[78]));
  INVX1 instanceL2_g9824(.Y(instanceL2_n_12334), .A(layer1_out[73]));
  INVX1 instanceL2_g9825(.Y(instanceL2_n_12335), .A(layer1_out[74]));
  INVX1 instanceL2_g9826(.Y(instanceL2_n_10991), .A(layer1_out[79]));
  INVX1 instanceL2_g9827(.Y(instanceL2_n_12336), .A(layer1_out[80]));
  XNOR2X1 instanceL2_g11223(.Y(\instanceL2_prod_terms[8][18] [10]), .A(
    instanceL2_n_12359), .B(instanceL2_n_12337));
  ADDFX1 instanceL2_g11224(.CO(instanceL2_n_12337), .S(
    \instanceL2_prod_terms[8][18] [9]), .A(instanceL2_n_12368), .B(
    instanceL2_n_12365), .CI(instanceL2_n_11065));
  ADDFX1 instanceL2_g11225(.CO(instanceL2_n_11065), .S(
    \instanceL2_prod_terms[8][18] [8]), .A(instanceL2_n_12364), .B(
    instanceL2_n_12357), .CI(instanceL2_n_12338));
  ADDFX1 instanceL2_g11226(.CO(instanceL2_n_12338), .S(
    \instanceL2_prod_terms[8][18] [7]), .A(instanceL2_n_12366), .B(
    instanceL2_n_12360), .CI(instanceL2_n_12339));
  OAI2BB1X1 instanceL2_g11227(.Y(\instanceL2_prod_terms[3][18] [9]), .A0N(
    layer1_out[168]), .A1N(instanceL2_n_12341), .B0(instanceL2_n_12340));
  ADDFX1 instanceL2_g11228(.CO(instanceL2_n_12339), .S(
    \instanceL2_prod_terms[8][18] [6]), .A(instanceL2_n_12363), .B(
    instanceL2_n_12356), .CI(instanceL2_n_11088));
  AND2XL instanceL2_g11229(.Y(\instanceL2_prod_terms[3][18] [10]), .A(
    layer1_out[169]), .B(instanceL2_n_12340));
  AOI2BB1XL instanceL2_g11230(.Y(\instanceL2_prod_terms[7][18] [8]), .A0N(
    layer1_out[169]), .A1N(instanceL2_n_12343), .B0(
    \instanceL2_prod_terms[7][18] [9]));
  OAI2BB1X1 instanceL2_g11231(.Y(\instanceL2_prod_terms[3][18] [8]), .A0N(
    layer1_out[167]), .A1N(instanceL2_n_12342), .B0(instanceL2_n_12341));
  XNOR2X1 instanceL2_g11232(.Y(\instanceL2_prod_terms[4][18] [9]), .A(
    layer1_out[169]), .B(instanceL2_n_12346));
  AND2X1 instanceL2_g11233(.Y(\instanceL2_prod_terms[7][18] [9]), .A(
    instanceL2_n_12343), .B(layer1_out[169]));
  NAND2BX1 instanceL2_g11234(.Y(instanceL2_n_12340), .AN(instanceL2_n_12342), .B(
    instanceL2_n_12382));
  XNOR2X1 instanceL2_g11235(.Y(\instanceL2_prod_terms[7][18] [7]), .A(
    instanceL2_n_12370), .B(instanceL2_n_12344));
  OR2XL instanceL2_g11236(.Y(instanceL2_n_12341), .A(layer1_out[167]), .B(
    instanceL2_n_12342));
  ADDFX1 instanceL2_g11237(.CO(instanceL2_n_11088), .S(
    \instanceL2_prod_terms[8][18] [5]), .A(instanceL2_n_12400), .B(
    instanceL2_n_12348), .CI(instanceL2_n_12358));
  OAI21X1 instanceL2_g11238(.Y(instanceL2_n_12342), .A0(instanceL2_n_12397), .A1(
    instanceL2_n_12347), .B0(instanceL2_n_12398));
  XNOR2X1 instanceL2_g11239(.Y(\instanceL2_prod_terms[3][18] [7]), .A(
    instanceL2_n_12374), .B(instanceL2_n_12347));
  OAI211X1 instanceL2_g11240(.Y(instanceL2_n_12343), .A0(instanceL2_n_12386),
     .A1(instanceL2_n_12345), .B0(instanceL2_n_12384), .C0(instanceL2_n_12380));
  NAND2X1 instanceL2_g11241(.Y(instanceL2_n_12344), .A(instanceL2_n_12384), .B(
    instanceL2_n_12345));
  AOI21X1 instanceL2_g11242(.Y(\instanceL2_prod_terms[4][18] [8]), .A0(
    layer1_out[168]), .A1(instanceL2_n_12352), .B0(instanceL2_n_12346));
  XNOR2X1 instanceL2_g11243(.Y(\instanceL2_prod_terms[7][18] [6]), .A(
    instanceL2_n_12368), .B(instanceL2_n_12349));
  NAND2BX1 instanceL2_g11244(.Y(\instanceL2_prod_terms[4][18] [13]), .AN(
    instanceL2_n_12352), .B(instanceL2_n_12386));
  NAND2BX1 instanceL2_g11245(.Y(instanceL2_n_12345), .AN(instanceL2_n_12382), .B(
    instanceL2_n_12349));
  NOR2X1 instanceL2_g11246(.Y(instanceL2_n_12346), .A(layer1_out[168]), .B(
    instanceL2_n_12352));
  XNOR2X1 instanceL2_g11247(.Y(\instanceL2_prod_terms[3][18] [6]), .A(
    instanceL2_n_12376), .B(instanceL2_n_11116));
  XNOR2X1 instanceL2_g11248(.Y(\instanceL2_prod_terms[7][18] [5]), .A(
    instanceL2_n_12373), .B(instanceL2_n_12350));
  AOI21X1 instanceL2_g11249(.Y(instanceL2_n_12347), .A0(instanceL2_n_12399), .A1(
    instanceL2_n_11116), .B0(instanceL2_n_12394));
  ADDFX1 instanceL2_g11250(.CO(instanceL2_n_12348), .S(
    \instanceL2_prod_terms[8][18] [4]), .A(layer1_out[165]), .B(
    instanceL2_n_12387), .CI(\instanceL2_prod_terms[4][18] [3]));
  OAI211X1 instanceL2_g11251(.Y(instanceL2_n_12349), .A0(instanceL2_n_12379),
     .A1(instanceL2_n_12351), .B0(instanceL2_n_12402), .C0(instanceL2_n_12381));
  OA21X1 instanceL2_g11252(.Y(\instanceL2_prod_terms[4][18] [7]), .A0(
    instanceL2_n_12410), .A1(instanceL2_n_12362), .B0(instanceL2_n_12352));
  NAND2X1 instanceL2_g11253(.Y(instanceL2_n_12350), .A(instanceL2_n_12402), .B(
    instanceL2_n_12351));
  OAI2BB1X1 instanceL2_g11254(.Y(instanceL2_n_11116), .A0N(instanceL2_n_12392),
     .A1N(instanceL2_n_11134), .B0(instanceL2_n_12393));
  XNOR2X1 instanceL2_g11255(.Y(\instanceL2_prod_terms[3][18] [5]), .A(
    instanceL2_n_12375), .B(instanceL2_n_11134));
  XNOR2X1 instanceL2_g11256(.Y(\instanceL2_prod_terms[7][18] [4]), .A(
    instanceL2_n_12371), .B(instanceL2_n_12354));
  XNOR2X1 instanceL2_g11257(.Y(\instanceL2_prod_terms[3][18] [3]), .A(
    layer1_out[165]), .B(instanceL2_n_12353));
  NAND2X1 instanceL2_g11258(.Y(instanceL2_n_12351), .A(instanceL2_n_12391), .B(
    instanceL2_n_12354));
  NAND2X1 instanceL2_g11259(.Y(instanceL2_n_12352), .A(instanceL2_n_12410), .B(
    instanceL2_n_12362));
  XNOR2X1 instanceL2_g11260(.Y(\instanceL2_prod_terms[7][18] [3]), .A(
    instanceL2_n_12355), .B(instanceL2_n_12372));
  MX2X1 instanceL2_g11261(.Y(\instanceL2_prod_terms[4][18] [5]), .A(
    layer1_out[165]), .B(instanceL2_n_12411), .S0(instanceL2_n_12369));
  NAND2XL instanceL2_g11262(.Y(instanceL2_n_12353), .A(instanceL2_n_11237), .B(
    instanceL2_n_12369));
  OAI2BB1X1 instanceL2_g11263(.Y(instanceL2_n_11134), .A0N(instanceL2_n_12395),
     .A1N(instanceL2_n_12361), .B0(instanceL2_n_12396));
  XNOR2X1 instanceL2_g11264(.Y(\instanceL2_prod_terms[3][18] [4]), .A(
    instanceL2_n_12377), .B(instanceL2_n_12361));
  XOR2XL instanceL2_g11265(.Y(\instanceL2_prod_terms[7][18] [2]), .A(
    instanceL2_n_11213), .B(instanceL2_n_12378));
  OAI211X1 instanceL2_g11266(.Y(instanceL2_n_12354), .A0(instanceL2_n_11213),
     .A1(instanceL2_n_12401), .B0(instanceL2_n_12383), .C0(instanceL2_n_11204));
  AOI21X1 instanceL2_g11267(.Y(\instanceL2_prod_terms[4][18] [6]), .A0(
    layer1_out[166]), .A1(instanceL2_n_12367), .B0(instanceL2_n_12362));
  NAND2X1 instanceL2_g11268(.Y(instanceL2_n_12355), .A(instanceL2_n_11213), .B(
    instanceL2_n_12383));
  MXI2XL instanceL2_g11269(.Y(instanceL2_n_12356), .A(layer1_out[165]), .B(
    instanceL2_n_12411), .S0(instanceL2_n_12375));
  MXI2XL instanceL2_g11270(.Y(instanceL2_n_12357), .A(instanceL2_n_12410), .B(
    layer1_out[167]), .S0(instanceL2_n_12374));
  XNOR2X1 instanceL2_g11271(.Y(instanceL2_n_12358), .A(layer1_out[164]), .B(
    instanceL2_n_12377));
  XNOR2X1 instanceL2_g11272(.Y(instanceL2_n_12359), .A(instanceL2_n_12404), .B(
    instanceL2_n_12370));
  XNOR2X1 instanceL2_g11273(.Y(instanceL2_n_12360), .A(layer1_out[166]), .B(
    instanceL2_n_12376));
  OA21X1 instanceL2_g11274(.Y(\instanceL2_prod_terms[4][18] [4]), .A0(
    instanceL2_n_12406), .A1(instanceL2_n_12385), .B0(instanceL2_n_12369));
  OAI2BB1X1 instanceL2_g11275(.Y(instanceL2_n_12361), .A0N(layer1_out[162]),
     .A1N(instanceL2_n_12411), .B0(instanceL2_n_12367));
  NOR2X1 instanceL2_g11276(.Y(instanceL2_n_12362), .A(layer1_out[166]), .B(
    instanceL2_n_12367));
  OAI22X1 instanceL2_g11277(.Y(instanceL2_n_12363), .A0(layer1_out[163]), .A1(
    instanceL2_n_12388), .B0(instanceL2_n_12407), .B1(instanceL2_n_12406));
  OAI22X1 instanceL2_g11278(.Y(instanceL2_n_12364), .A0(layer1_out[165]), .A1(
    instanceL2_n_12389), .B0(instanceL2_n_12405), .B1(instanceL2_n_12407));
  OAI22X1 instanceL2_g11279(.Y(instanceL2_n_12365), .A0(layer1_out[166]), .A1(
    instanceL2_n_12390), .B0(instanceL2_n_12409), .B1(instanceL2_n_12410));
  OAI22X1 instanceL2_g11280(.Y(instanceL2_n_12366), .A0(layer1_out[164]), .A1(
    instanceL2_n_12403), .B0(instanceL2_n_12410), .B1(instanceL2_n_12411));
  NAND2XL instanceL2_g11281(.Y(instanceL2_n_12371), .A(instanceL2_n_12402), .B(
    instanceL2_n_12391));
  NAND2BX1 instanceL2_g11282(.Y(instanceL2_n_12372), .AN(instanceL2_n_12401), .B(
    instanceL2_n_11204));
  NAND2BX1 instanceL2_g11283(.Y(instanceL2_n_12373), .AN(instanceL2_n_12379), .B(
    instanceL2_n_12381));
  NAND2X1 instanceL2_g11284(.Y(instanceL2_n_12367), .A(instanceL2_n_12385), .B(
    instanceL2_n_12401));
  NAND2BX1 instanceL2_g11285(.Y(instanceL2_n_12368), .AN(instanceL2_n_12382), .B(
    instanceL2_n_12384));
  NAND2X1 instanceL2_g11286(.Y(instanceL2_n_12369), .A(instanceL2_n_12406), .B(
    instanceL2_n_12385));
  NAND2BX1 instanceL2_g11287(.Y(instanceL2_n_12370), .AN(instanceL2_n_12386), .B(
    instanceL2_n_12380));
  AOI21X1 instanceL2_g11288(.Y(\instanceL2_prod_terms[8][18] [3]), .A0(
    instanceL2_n_11237), .A1(instanceL2_n_12406), .B0(instanceL2_n_12387));
  OAI21X1 instanceL2_g11289(.Y(instanceL2_n_12378), .A0(layer1_out[164]), .A1(
    layer1_out[163]), .B0(instanceL2_n_12383));
  NOR2BX1 instanceL2_g11290(.Y(instanceL2_n_12374), .AN(instanceL2_n_12398), .B(
    instanceL2_n_12397));
  NAND2X1 instanceL2_g11291(.Y(instanceL2_n_12375), .A(instanceL2_n_12392), .B(
    instanceL2_n_12393));
  OAI2BB1X1 instanceL2_g11292(.Y(\instanceL2_prod_terms[4][18] [3]), .A0N(
    layer1_out[163]), .A1N(instanceL2_n_11237), .B0(instanceL2_n_12400));
  NAND2BX1 instanceL2_g11293(.Y(instanceL2_n_12376), .AN(instanceL2_n_12394), .B(
    instanceL2_n_12399));
  NAND2X1 instanceL2_g10277(.Y(instanceL2_n_12377), .A(instanceL2_n_12395), .B(
    instanceL2_n_12396));
  NOR2XL instanceL2_g10278(.Y(instanceL2_n_12388), .A(layer1_out[166]), .B(
    layer1_out[164]));
  NOR2XL instanceL2_g10279(.Y(instanceL2_n_12389), .A(layer1_out[168]), .B(
    layer1_out[166]));
  NOR2XL instanceL2_g10280(.Y(instanceL2_n_12390), .A(layer1_out[169]), .B(
    layer1_out[167]));
  NAND2XL instanceL2_g10281(.Y(instanceL2_n_11204), .A(layer1_out[164]), .B(
    layer1_out[165]));
  NOR2X1 instanceL2_g10282(.Y(instanceL2_n_12379), .A(layer1_out[167]), .B(
    layer1_out[166]));
  NAND2X1 instanceL2_g10283(.Y(instanceL2_n_12380), .A(layer1_out[169]), .B(
    layer1_out[168]));
  NAND2XL instanceL2_g10284(.Y(instanceL2_n_12381), .A(layer1_out[167]), .B(
    layer1_out[166]));
  NOR2XL instanceL2_g10285(.Y(instanceL2_n_12382), .A(layer1_out[168]), .B(
    layer1_out[167]));
  NAND2XL instanceL2_g10286(.Y(instanceL2_n_12383), .A(layer1_out[163]), .B(
    layer1_out[164]));
  NAND2X1 instanceL2_g10287(.Y(instanceL2_n_12384), .A(layer1_out[167]), .B(
    layer1_out[168]));
  NOR2X1 instanceL2_g10288(.Y(instanceL2_n_12385), .A(layer1_out[162]), .B(
    layer1_out[163]));
  NOR2X1 instanceL2_g10289(.Y(instanceL2_n_12386), .A(layer1_out[169]), .B(
    layer1_out[168]));
  NAND2XL instanceL2_g10290(.Y(instanceL2_n_11213), .A(layer1_out[162]), .B(
    layer1_out[163]));
  NOR2X1 instanceL2_g10291(.Y(instanceL2_n_12387), .A(instanceL2_n_11237), .B(
    instanceL2_n_12406));
  NOR2XL instanceL2_g10292(.Y(instanceL2_n_12403), .A(layer1_out[167]), .B(
    layer1_out[165]));
  NAND2X1 instanceL2_g10293(.Y(instanceL2_n_12391), .A(instanceL2_n_12407), .B(
    instanceL2_n_12411));
  NAND2X1 instanceL2_g10294(.Y(instanceL2_n_12392), .A(layer1_out[167]), .B(
    instanceL2_n_12406));
  NAND2X1 instanceL2_g10295(.Y(instanceL2_n_12393), .A(instanceL2_n_12410), .B(
    layer1_out[164]));
  NOR2XL instanceL2_g10296(.Y(instanceL2_n_12394), .A(layer1_out[168]), .B(
    instanceL2_n_12411));
  NAND2XL instanceL2_g10297(.Y(instanceL2_n_12395), .A(instanceL2_n_12408), .B(
    layer1_out[166]));
  NAND2X1 instanceL2_g10298(.Y(instanceL2_n_12396), .A(layer1_out[163]), .B(
    instanceL2_n_12407));
  NOR2X1 instanceL2_g10299(.Y(instanceL2_n_12397), .A(instanceL2_n_12409), .B(
    layer1_out[166]));
  NAND2X1 instanceL2_g10300(.Y(instanceL2_n_12398), .A(instanceL2_n_12409), .B(
    layer1_out[166]));
  NOR2XL instanceL2_g10301(.Y(instanceL2_n_12404), .A(instanceL2_n_12405), .B(
    layer1_out[167]));
  NAND2X1 instanceL2_g10302(.Y(instanceL2_n_12399), .A(layer1_out[168]), .B(
    instanceL2_n_12411));
  NAND2X1 instanceL2_g10303(.Y(instanceL2_n_12400), .A(layer1_out[162]), .B(
    instanceL2_n_12408));
  NOR2X1 instanceL2_g10304(.Y(instanceL2_n_12401), .A(layer1_out[164]), .B(
    layer1_out[165]));
  NAND2XL instanceL2_g10305(.Y(instanceL2_n_12402), .A(layer1_out[166]), .B(
    layer1_out[165]));
  INVX1 instanceL2_g10306(.Y(instanceL2_n_11237), .A(layer1_out[162]));
  INVX1 instanceL2_g10307(.Y(instanceL2_n_12405), .A(layer1_out[168]));
  INVX1 instanceL2_g10308(.Y(instanceL2_n_12406), .A(layer1_out[164]));
  INVX1 instanceL2_g11294(.Y(instanceL2_n_12407), .A(layer1_out[166]));
  INVX1 instanceL2_g11295(.Y(instanceL2_n_12408), .A(layer1_out[163]));
  INVX1 instanceL2_g11296(.Y(instanceL2_n_12409), .A(layer1_out[169]));
  INVX1 instanceL2_g11297(.Y(instanceL2_n_12410), .A(layer1_out[167]));
  INVX1 instanceL2_g11298(.Y(instanceL2_n_12411), .A(layer1_out[165]));
  XNOR2X1 instanceL2_g11299(.Y(\instanceL2_prod_terms[7][9][11] ), .A(
    layer1_out[89]), .B(instanceL2_n_12412));
  XNOR2X1 instanceL2_g11300(.Y(\instanceL2_prod_terms[7][9][10] ), .A(
    layer1_out[88]), .B(instanceL2_n_12413));
  NOR2X1 instanceL2_g11301(.Y(\instanceL2_prod_terms[7][9][12] ), .A(
    instanceL2_n_11035), .B(instanceL2_n_12413));
  MX2XL instanceL2_g11302(.Y(\instanceL2_prod_terms[7][9][9] ), .A(
    layer1_out[87]), .B(instanceL2_n_11040), .S0(instanceL2_n_12414));
  OA22X1 instanceL2_g11303(.Y(instanceL2_n_12412), .A0(instanceL2_n_12447), .A1(
    instanceL2_n_12415), .B0(instanceL2_n_11035), .B1(instanceL2_n_12434));
  AND2X1 instanceL2_g11304(.Y(instanceL2_n_12413), .A(instanceL2_n_12415), .B(
    instanceL2_n_12434));
  NAND2XL instanceL2_g11305(.Y(instanceL2_n_12414), .A(instanceL2_n_12444), .B(
    instanceL2_n_12416));
  XNOR2X1 instanceL2_g11306(.Y(\instanceL2_prod_terms[7][9][8] ), .A(
    instanceL2_n_10999), .B(instanceL2_n_12417));
  OR2XL instanceL2_g11307(.Y(instanceL2_n_12415), .A(instanceL2_n_11040), .B(
    instanceL2_n_12416));
  NAND2BX1 instanceL2_g11308(.Y(instanceL2_n_12416), .AN(instanceL2_n_11018), .B(
    instanceL2_n_12417));
  OA21X1 instanceL2_g11309(.Y(\instanceL2_prod_terms[2][9] [10]), .A0(
    instanceL2_n_11048), .A1(instanceL2_n_12419), .B0(
    \instanceL2_prod_terms[2][9] [13]));
  XNOR2X1 instanceL2_g11310(.Y(\instanceL2_prod_terms[3][9] [9]), .A(
    layer1_out[89]), .B(instanceL2_n_12418));
  ADDFX1 instanceL2_g11311(.CO(instanceL2_n_12417), .S(
    \instanceL2_prod_terms[7][9][7] ), .A(layer1_out[85]), .B(layer1_out[88]),
     .CI(instanceL2_n_12420));
  NAND2X1 instanceL2_g11312(.Y(\instanceL2_prod_terms[2][9] [13]), .A(
    instanceL2_n_11048), .B(instanceL2_n_12419));
  AOI21X1 instanceL2_g11313(.Y(instanceL2_n_12418), .A0(layer1_out[88]), .A1(
    instanceL2_n_12421), .B0(\instanceL2_prod_terms[3][9] [10]));
  OAI2BB1X1 instanceL2_g11314(.Y(\instanceL2_prod_terms[3][9] [10]), .A0N(
    layer1_out[89]), .A1N(instanceL2_n_12421), .B0(instanceL2_n_11035));
  AOI21X1 instanceL2_g11315(.Y(\instanceL2_prod_terms[2][9] [9]), .A0(
    layer1_out[88]), .A1(instanceL2_n_12423), .B0(instanceL2_n_12419));
  XNOR2X1 instanceL2_g11316(.Y(\instanceL2_prod_terms[3][9] [8]), .A(
    instanceL2_n_12438), .B(instanceL2_n_12421));
  ADDFX1 instanceL2_g11317(.CO(instanceL2_n_12420), .S(
    \instanceL2_prod_terms[7][9][6] ), .A(layer1_out[84]), .B(layer1_out[87]),
     .CI(instanceL2_n_12424));
  NOR2X1 instanceL2_g11318(.Y(instanceL2_n_12419), .A(layer1_out[88]), .B(
    instanceL2_n_12423));
  XNOR2X1 instanceL2_g11319(.Y(\instanceL2_prod_terms[3][9] [7]), .A(
    instanceL2_n_11009), .B(instanceL2_n_12422));
  OAI211X1 instanceL2_g11320(.Y(instanceL2_n_12421), .A0(instanceL2_n_11028),
     .A1(instanceL2_n_12425), .B0(instanceL2_n_11034), .C0(instanceL2_n_12440));
  NAND2X1 instanceL2_g11321(.Y(instanceL2_n_12422), .A(instanceL2_n_11034), .B(
    instanceL2_n_12425));
  OA21X1 instanceL2_g11322(.Y(\instanceL2_prod_terms[2][9] [8]), .A0(
    instanceL2_n_11040), .A1(instanceL2_n_12429), .B0(instanceL2_n_12423));
  XNOR2X1 instanceL2_g11323(.Y(\instanceL2_prod_terms[3][9] [6]), .A(
    instanceL2_n_10994), .B(instanceL2_n_12426));
  ADDFX1 instanceL2_g11324(.CO(instanceL2_n_12424), .S(
    \instanceL2_prod_terms[7][9][5] ), .A(layer1_out[86]), .B(layer1_out[83]),
     .CI(instanceL2_n_12430));
  NAND2X1 instanceL2_g11325(.Y(instanceL2_n_12423), .A(instanceL2_n_11040), .B(
    instanceL2_n_12429));
  XNOR2X1 instanceL2_g11326(.Y(\instanceL2_prod_terms[3][9] [5]), .A(
    instanceL2_n_11006), .B(instanceL2_n_12427));
  NAND2BX1 instanceL2_g11327(.Y(instanceL2_n_12425), .AN(instanceL2_n_12443), .B(
    instanceL2_n_12426));
  OAI211X1 instanceL2_g11328(.Y(instanceL2_n_12426), .A0(instanceL2_n_11029),
     .A1(instanceL2_n_12428), .B0(instanceL2_n_11032), .C0(instanceL2_n_12445));
  NAND2X1 instanceL2_g11329(.Y(instanceL2_n_12427), .A(instanceL2_n_11032), .B(
    instanceL2_n_12428));
  AOI21X1 instanceL2_g11330(.Y(\instanceL2_prod_terms[2][9] [7]), .A0(
    layer1_out[86]), .A1(instanceL2_n_12431), .B0(instanceL2_n_12429));
  XNOR2X1 instanceL2_g11331(.Y(\instanceL2_prod_terms[3][9] [4]), .A(
    instanceL2_n_12436), .B(instanceL2_n_12432));
  ADDFX1 instanceL2_g11332(.CO(instanceL2_n_12430), .S(
    \instanceL2_prod_terms[7][9][4] ), .A(layer1_out[85]), .B(layer1_out[82]),
     .CI(instanceL2_n_11024));
  NAND2BX1 instanceL2_g11333(.Y(instanceL2_n_12428), .AN(instanceL2_n_12446), .B(
    instanceL2_n_12432));
  NOR2X1 instanceL2_g11334(.Y(instanceL2_n_12429), .A(layer1_out[86]), .B(
    instanceL2_n_12431));
  XNOR2X1 instanceL2_g11335(.Y(\instanceL2_prod_terms[3][9] [3]), .A(
    instanceL2_n_12435), .B(instanceL2_n_12433));
  XNOR2X1 instanceL2_g11336(.Y(\instanceL2_prod_terms[2][9] [5]), .A(
    layer1_out[84]), .B(instanceL2_n_12437));
  NAND2X1 instanceL2_g11337(.Y(instanceL2_n_12431), .A(instanceL2_n_12446), .B(
    instanceL2_n_12437));
  XOR2XL instanceL2_g11338(.Y(\instanceL2_prod_terms[3][9] [2]), .A(
    instanceL2_n_12442), .B(instanceL2_n_11015));
  OAI211X1 instanceL2_g11339(.Y(instanceL2_n_12432), .A0(instanceL2_n_12441),
     .A1(instanceL2_n_12442), .B0(instanceL2_n_11021), .C0(instanceL2_n_12439));
  NAND2XL instanceL2_g11340(.Y(instanceL2_n_12433), .A(instanceL2_n_11021), .B(
    instanceL2_n_12442));
  AOI21X1 instanceL2_g11341(.Y(\instanceL2_prod_terms[2][9] [4]), .A0(
    layer1_out[83]), .A1(instanceL2_n_11022), .B0(instanceL2_n_12437));
  AND2X1 instanceL2_g11342(.Y(\instanceL2_prod_terms[2][9] [3]), .A(
    instanceL2_n_11022), .B(instanceL2_n_12442));
  NAND2BX1 instanceL2_g11343(.Y(instanceL2_n_10994), .AN(instanceL2_n_12443), .B(
    instanceL2_n_11034));
  NAND2BXL instanceL2_g11344(.Y(instanceL2_n_12435), .AN(instanceL2_n_12441), .B(
    instanceL2_n_12439));
  NAND2BX1 instanceL2_g11345(.Y(instanceL2_n_10999), .AN(instanceL2_n_11018), .B(
    instanceL2_n_12444));
  NAND2BX1 instanceL2_g11346(.Y(instanceL2_n_12436), .AN(instanceL2_n_12446), .B(
    instanceL2_n_11032));
  OR2XL instanceL2_g11347(.Y(instanceL2_n_12434), .A(instanceL2_n_11048), .B(
    instanceL2_n_11034));
  AOI2BB1X1 instanceL2_g11348(.Y(\instanceL2_prod_terms[7][9][3] ), .A0N(
    layer1_out[84]), .A1N(layer1_out[81]), .B0(instanceL2_n_11024));
  NAND2BX1 instanceL2_g11349(.Y(instanceL2_n_11006), .AN(instanceL2_n_11029), .B(
    instanceL2_n_12445));
  NAND2BXL instanceL2_g11350(.Y(instanceL2_n_11009), .AN(instanceL2_n_11028), .B(
    instanceL2_n_12440));
  NAND2BX1 instanceL2_g11351(.Y(instanceL2_n_11012), .AN(instanceL2_n_11022), .B(
    instanceL2_n_12441));
  OAI2BB1X1 instanceL2_g11352(.Y(instanceL2_n_12438), .A0N(instanceL2_n_12447),
     .A1N(instanceL2_n_11048), .B0(instanceL2_n_11035));
  OAI21X1 instanceL2_g11353(.Y(instanceL2_n_11015), .A0(layer1_out[83]), .A1(
    layer1_out[82]), .B0(instanceL2_n_11021));
  NOR2X1 instanceL2_g11354(.Y(instanceL2_n_12437), .A(layer1_out[83]), .B(
    instanceL2_n_11022));
  NAND2XL instanceL2_g11355(.Y(instanceL2_n_12439), .A(layer1_out[84]), .B(
    layer1_out[83]));
  NOR2XL instanceL2_g11356(.Y(instanceL2_n_11018), .A(layer1_out[86]), .B(
    layer1_out[89]));
  NAND2XL instanceL2_g11357(.Y(instanceL2_n_12440), .A(layer1_out[88]), .B(
    layer1_out[87]));
  NOR2X1 instanceL2_g11358(.Y(instanceL2_n_12441), .A(layer1_out[84]), .B(
    layer1_out[83]));
  NAND2XL instanceL2_g11359(.Y(instanceL2_n_11021), .A(layer1_out[82]), .B(
    layer1_out[83]));
  OR2X1 instanceL2_g11360(.Y(instanceL2_n_11022), .A(layer1_out[82]), .B(
    layer1_out[81]));
  AND2XL instanceL2_g11361(.Y(instanceL2_n_11024), .A(layer1_out[84]), .B(
    layer1_out[81]));
  NAND2XL instanceL2_g11362(.Y(instanceL2_n_12442), .A(layer1_out[82]), .B(
    layer1_out[81]));
  NOR2XL instanceL2_g11363(.Y(instanceL2_n_12443), .A(layer1_out[86]), .B(
    layer1_out[87]));
  NOR2XL instanceL2_g11364(.Y(instanceL2_n_11028), .A(layer1_out[88]), .B(
    layer1_out[87]));
  NOR2X1 instanceL2_g11365(.Y(instanceL2_n_11029), .A(layer1_out[85]), .B(
    layer1_out[86]));
  NAND2XL instanceL2_g11366(.Y(instanceL2_n_12444), .A(layer1_out[86]), .B(
    layer1_out[89]));
  NAND2XL instanceL2_g11367(.Y(instanceL2_n_12445), .A(layer1_out[85]), .B(
    layer1_out[86]));
  NAND2X1 instanceL2_g11368(.Y(instanceL2_n_11032), .A(layer1_out[84]), .B(
    layer1_out[85]));
  NOR2X1 instanceL2_g11369(.Y(instanceL2_n_12446), .A(layer1_out[84]), .B(
    layer1_out[85]));
  NAND2X1 instanceL2_g11370(.Y(instanceL2_n_11034), .A(layer1_out[86]), .B(
    layer1_out[87]));
  NAND2X1 instanceL2_g11371(.Y(instanceL2_n_11035), .A(layer1_out[88]), .B(
    layer1_out[89]));
  INVX1 instanceL2_g11372(.Y(instanceL2_n_11040), .A(layer1_out[87]));
  INVX1 instanceL2_g11373(.Y(instanceL2_n_12447), .A(layer1_out[88]));
  INVX1 instanceL2_g11374(.Y(instanceL2_n_11048), .A(layer1_out[89]));
  CLKXOR2X1 instanceL2_g11375(.Y(\instanceL2_prod_terms[2][9] [6]), .A(
    layer1_out[85]), .B(instanceL2_n_11012));
  XNOR2X1 instanceL2_g11376(.Y(\instanceL2_prod_terms[8][7] [10]), .A(
    layer1_out[70]), .B(instanceL2_n_10790));
  AOI2BB1X1 instanceL2_g9648(.Y(\instanceL2_prod_terms[3][7] [8]), .A0N(
    layer1_out[70]), .A1N(instanceL2_n_10791), .B0(
    \instanceL2_prod_terms[3][7] [9]));
  AOI21X1 instanceL2_g9649(.Y(\instanceL2_prod_terms[8][7] [11]), .A0(
    instanceL2_n_12487), .A1(instanceL2_n_12448), .B0(instanceL2_n_12481));
  OAI21X1 instanceL2_g9650(.Y(instanceL2_n_10784), .A0(instanceL2_n_12486), .A1(
    instanceL2_n_12448), .B0(instanceL2_n_12487));
  AND2X1 instanceL2_g9651(.Y(\instanceL2_prod_terms[3][7] [9]), .A(
    instanceL2_n_10791), .B(layer1_out[70]));
  XNOR2X1 instanceL2_g9652(.Y(\instanceL2_prod_terms[8][7] [8]), .A(
    instanceL2_n_12463), .B(instanceL2_n_12448));
  XNOR2X1 instanceL2_g9653(.Y(\instanceL2_prod_terms[3][7] [7]), .A(
    instanceL2_n_12466), .B(instanceL2_n_10797));
  AOI22X1 instanceL2_g9654(.Y(instanceL2_n_10790), .A0(instanceL2_n_12461), .A1(
    instanceL2_n_12449), .B0(layer1_out[68]), .B1(instanceL2_n_10888));
  OAI211X1 instanceL2_g9655(.Y(instanceL2_n_10791), .A0(instanceL2_n_12492), .A1(
    instanceL2_n_12450), .B0(instanceL2_n_12481), .C0(instanceL2_n_12489));
  INVX1 instanceL2_g9656(.Y(instanceL2_n_12448), .A(instanceL2_n_12449));
  ADDFX1 instanceL2_g9657(.CO(instanceL2_n_12449), .S(
    \instanceL2_prod_terms[8][7] [7]), .A(layer1_out[69]), .B(layer1_out[67]),
     .CI(instanceL2_n_10809));
  NAND2X1 instanceL2_g9658(.Y(instanceL2_n_10797), .A(instanceL2_n_12489), .B(
    instanceL2_n_12450));
  XNOR2X1 instanceL2_g9659(.Y(\instanceL2_prod_terms[3][7] [6]), .A(
    instanceL2_n_10874), .B(instanceL2_n_12451));
  NAND2BX1 instanceL2_g9660(.Y(instanceL2_n_12450), .AN(instanceL2_n_12479), .B(
    instanceL2_n_12451));
  CLKXOR2X1 instanceL2_g9661(.Y(\instanceL2_prod_terms[3][7] [5]), .A(
    instanceL2_n_12469), .B(instanceL2_n_12452));
  OAI22X1 instanceL2_g9662(.Y(instanceL2_n_12451), .A0(instanceL2_n_12476), .A1(
    instanceL2_n_10816), .B0(instanceL2_n_12494), .B1(instanceL2_n_12490));
  XNOR2X1 instanceL2_g9663(.Y(\instanceL2_prod_terms[0][7] [8]), .A(
    layer1_out[70]), .B(instanceL2_n_10817));
  XNOR2X1 instanceL2_g9664(.Y(\instanceL2_prod_terms[3][7] [4]), .A(
    instanceL2_n_12470), .B(instanceL2_n_12456));
  NAND2X1 instanceL2_g9665(.Y(instanceL2_n_12452), .A(instanceL2_n_12473), .B(
    instanceL2_n_10816));
  OAI21X1 instanceL2_g9666(.Y(instanceL2_n_10809), .A0(instanceL2_n_12490), .A1(
    instanceL2_n_12455), .B0(instanceL2_n_12484));
  XNOR2X1 instanceL2_g9667(.Y(\instanceL2_prod_terms[8][7] [6]), .A(
    instanceL2_n_12465), .B(instanceL2_n_12455));
  XNOR2X1 instanceL2_g9668(.Y(\instanceL2_prod_terms[8][7] [5]), .A(
    instanceL2_n_12462), .B(instanceL2_n_12454));
  XNOR2X1 instanceL2_g9669(.Y(\instanceL2_prod_terms[0][7] [6]), .A(
    layer1_out[68]), .B(instanceL2_n_12453));
  AND2XL instanceL2_g9670(.Y(instanceL2_n_10817), .A(instanceL2_n_12479), .B(
    instanceL2_n_12453));
  NAND2BX1 instanceL2_g9671(.Y(instanceL2_n_10816), .AN(instanceL2_n_12488), .B(
    instanceL2_n_12456));
  XNOR2X1 instanceL2_g9672(.Y(\instanceL2_prod_terms[3][7] [3]), .A(
    instanceL2_n_12458), .B(instanceL2_n_12472));
  XNOR2X1 instanceL2_g9673(.Y(\instanceL2_prod_terms[0][7] [7]), .A(
    layer1_out[69]), .B(instanceL2_n_12457));
  XNOR2X1 instanceL2_g9674(.Y(\instanceL2_prod_terms[0][7] [4]), .A(
    layer1_out[66]), .B(instanceL2_n_12468));
  NAND2X2 instanceL2_g9675(.Y(\instanceL2_prod_terms[0][7] [13]), .A(
    instanceL2_n_12492), .B(instanceL2_n_12457));
  NAND2BX1 instanceL2_g9676(.Y(instanceL2_n_12454), .AN(instanceL2_n_12459), .B(
    instanceL2_n_12478));
  AND2XL instanceL2_g9677(.Y(instanceL2_n_12453), .A(instanceL2_n_12488), .B(
    instanceL2_n_12468));
  XNOR2X1 instanceL2_g9678(.Y(\instanceL2_prod_terms[8][7] [4]), .A(
    instanceL2_n_12480), .B(instanceL2_n_12464));
  CLKXOR2X1 instanceL2_g9679(.Y(\instanceL2_prod_terms[3][7] [2]), .A(
    instanceL2_n_12482), .B(instanceL2_n_12471));
  NOR2X1 instanceL2_g9680(.Y(instanceL2_n_12455), .A(instanceL2_n_12459), .B(
    instanceL2_n_12460));
  OAI211X1 instanceL2_g9681(.Y(instanceL2_n_12456), .A0(instanceL2_n_12482), .A1(
    instanceL2_n_12491), .B0(instanceL2_n_12477), .C0(instanceL2_n_12483));
  NAND2XL instanceL2_g9682(.Y(instanceL2_n_12458), .A(instanceL2_n_12477), .B(
    instanceL2_n_12482));
  NOR2BX1 instanceL2_g9683(.Y(instanceL2_n_12457), .AN(instanceL2_n_12476), .B(
    instanceL2_n_12467));
  XNOR2X1 instanceL2_g9684(.Y(\instanceL2_prod_terms[4][7] [6]), .A(
    instanceL2_n_12494), .B(instanceL2_n_12467));
  NOR2X1 instanceL2_g9685(.Y(instanceL2_n_12459), .A(instanceL2_n_12474), .B(
    instanceL2_n_12480));
  OAI21X1 instanceL2_g9686(.Y(instanceL2_n_12460), .A0(instanceL2_n_12478), .A1(
    instanceL2_n_12475), .B0(instanceL2_n_12485));
  AOI21X1 instanceL2_g9687(.Y(\instanceL2_prod_terms[0][7] [3]), .A0(
    layer1_out[65]), .A1(instanceL2_n_12493), .B0(instanceL2_n_12468));
  AND2X1 instanceL2_g9688(.Y(\instanceL2_prod_terms[0][7] [2]), .A(
    instanceL2_n_12493), .B(instanceL2_n_12482));
  NAND2XL instanceL2_g9689(.Y(instanceL2_n_12461), .A(instanceL2_n_12481), .B(
    instanceL2_n_12489));
  NAND2BXL instanceL2_g9690(.Y(instanceL2_n_12462), .AN(instanceL2_n_12475), .B(
    instanceL2_n_12485));
  NOR2BX1 instanceL2_g9691(.Y(instanceL2_n_12463), .AN(instanceL2_n_12487), .B(
    instanceL2_n_12486));
  NOR2BX1 instanceL2_g9692(.Y(instanceL2_n_12464), .AN(instanceL2_n_12478), .B(
    instanceL2_n_12474));
  NOR2BX1 instanceL2_g9693(.Y(instanceL2_n_12465), .AN(instanceL2_n_12484), .B(
    instanceL2_n_12490));
  NAND2BXL instanceL2_g9694(.Y(instanceL2_n_12466), .AN(instanceL2_n_12492), .B(
    instanceL2_n_12481));
  OA21X1 instanceL2_g9695(.Y(\instanceL2_prod_terms[8][7] [3]), .A0(
    layer1_out[65]), .A1(layer1_out[63]), .B0(instanceL2_n_12480));
  AOI21XL instanceL2_g9696(.Y(instanceL2_n_12469), .A0(layer1_out[68]), .A1(
    layer1_out[67]), .B0(instanceL2_n_12476));
  NAND2BXL instanceL2_g9697(.Y(instanceL2_n_12470), .AN(instanceL2_n_12488), .B(
    instanceL2_n_12473));
  NAND2BXL instanceL2_g9698(.Y(instanceL2_n_10874), .AN(instanceL2_n_12479), .B(
    instanceL2_n_12489));
  OAI21X1 instanceL2_g9699(.Y(instanceL2_n_12471), .A0(layer1_out[64]), .A1(
    layer1_out[65]), .B0(instanceL2_n_12477));
  NAND2BX1 instanceL2_g9700(.Y(instanceL2_n_12472), .AN(instanceL2_n_12491), .B(
    instanceL2_n_12483));
  NAND2BX1 instanceL2_g9701(.Y(instanceL2_n_12467), .AN(instanceL2_n_12493), .B(
    instanceL2_n_12491));
  NOR2X1 instanceL2_g9702(.Y(instanceL2_n_12468), .A(layer1_out[65]), .B(
    instanceL2_n_12493));
  INVX1 instanceL2_g9703(.Y(instanceL2_n_10888), .A(instanceL2_n_12481));
  NAND2XL instanceL2_g9704(.Y(instanceL2_n_12473), .A(layer1_out[66]), .B(
    layer1_out[67]));
  NOR2X1 instanceL2_g9705(.Y(instanceL2_n_12474), .A(layer1_out[64]), .B(
    layer1_out[66]));
  NOR2X1 instanceL2_g9706(.Y(instanceL2_n_12475), .A(layer1_out[65]), .B(
    layer1_out[67]));
  NOR2X1 instanceL2_g9707(.Y(instanceL2_n_12476), .A(layer1_out[68]), .B(
    layer1_out[67]));
  NAND2X1 instanceL2_g9708(.Y(instanceL2_n_12477), .A(layer1_out[64]), .B(
    layer1_out[65]));
  NAND2X1 instanceL2_g9709(.Y(instanceL2_n_12478), .A(layer1_out[64]), .B(
    layer1_out[66]));
  NOR2X1 instanceL2_g9710(.Y(instanceL2_n_12479), .A(layer1_out[69]), .B(
    layer1_out[68]));
  NAND2X1 instanceL2_g9711(.Y(instanceL2_n_12480), .A(layer1_out[65]), .B(
    layer1_out[63]));
  NAND2X1 instanceL2_g9712(.Y(instanceL2_n_12481), .A(layer1_out[69]), .B(
    layer1_out[70]));
  NAND2X1 instanceL2_g9713(.Y(instanceL2_n_12482), .A(layer1_out[64]), .B(
    layer1_out[63]));
  NAND2XL instanceL2_g9714(.Y(instanceL2_n_12483), .A(layer1_out[66]), .B(
    layer1_out[65]));
  NAND2XL instanceL2_g9715(.Y(instanceL2_n_12484), .A(layer1_out[66]), .B(
    layer1_out[68]));
  NAND2XL instanceL2_g9716(.Y(instanceL2_n_12485), .A(layer1_out[65]), .B(
    layer1_out[67]));
  NOR2X1 instanceL2_g9717(.Y(instanceL2_n_12486), .A(layer1_out[70]), .B(
    layer1_out[68]));
  NAND2X1 instanceL2_g9718(.Y(instanceL2_n_12487), .A(layer1_out[70]), .B(
    layer1_out[68]));
  NOR2X1 instanceL2_g9719(.Y(instanceL2_n_12488), .A(layer1_out[66]), .B(
    layer1_out[67]));
  NAND2X1 instanceL2_g9720(.Y(instanceL2_n_12489), .A(layer1_out[69]), .B(
    layer1_out[68]));
  NOR2X1 instanceL2_g9721(.Y(instanceL2_n_12490), .A(layer1_out[66]), .B(
    layer1_out[68]));
  NOR2X1 instanceL2_g9722(.Y(instanceL2_n_12491), .A(layer1_out[65]), .B(
    layer1_out[66]));
  NOR2X1 instanceL2_g9723(.Y(instanceL2_n_12492), .A(layer1_out[69]), .B(
    layer1_out[70]));
  OR2X1 instanceL2_g9724(.Y(instanceL2_n_12493), .A(layer1_out[64]), .B(
    layer1_out[63]));
  INVX1 instanceL2_g9726(.Y(instanceL2_n_12494), .A(layer1_out[67]));
  XOR2XL instanceL2_g11377(.Y(\instanceL2_prod_terms[8][7] [9]), .A(
    layer1_out[69]), .B(instanceL2_n_10784));
  XNOR2X1 instanceL2_g11378(.Y(\instanceL2_prod_terms[7][5] [10]), .A(
    instanceL2_n_11110), .B(instanceL2_n_12495));
  ADDFX1 instanceL2_g11379(.CO(instanceL2_n_12495), .S(
    \instanceL2_prod_terms[7][5] [9]), .A(instanceL2_n_12553), .B(
    instanceL2_n_12533), .CI(instanceL2_n_12496));
  ADDFX1 instanceL2_g11380(.CO(instanceL2_n_12496), .S(
    \instanceL2_prod_terms[7][5] [8]), .A(instanceL2_n_12531), .B(
    instanceL2_n_12514), .CI(instanceL2_n_12498));
  NAND2X1 instanceL2_g11381(.Y(\instanceL2_prod_terms[0][5][9] ), .A(
    instanceL2_n_12499), .B(instanceL2_n_12497));
  OAI211X1 instanceL2_g11382(.Y(instanceL2_n_12497), .A0(instanceL2_n_12548),
     .A1(instanceL2_n_12500), .B0(instanceL2_n_12561), .C0(layer1_out[52]));
  XNOR2X1 instanceL2_g11383(.Y(\instanceL2_prod_terms[0][5][8] ), .A(
    instanceL2_n_12519), .B(instanceL2_n_12500));
  ADDFX1 instanceL2_g11384(.CO(instanceL2_n_12498), .S(
    \instanceL2_prod_terms[7][5] [7]), .A(instanceL2_n_12516), .B(
    instanceL2_n_12513), .CI(instanceL2_n_11046));
  OAI2BB1X1 instanceL2_g11385(.Y(instanceL2_n_12499), .A0N(instanceL2_n_12561),
     .A1N(instanceL2_n_12502), .B0(instanceL2_n_12559));
  ADDFX1 instanceL2_g11386(.CO(instanceL2_n_12500), .S(
    \instanceL2_prod_terms[0][5][7] ), .A(instanceL2_n_12552), .B(
    instanceL2_n_12529), .CI(instanceL2_n_12501));
  XNOR2X1 instanceL2_g11387(.Y(\instanceL2_prod_terms[2][5] [7]), .A(
    layer1_out[51]), .B(instanceL2_n_12502));
  ADDFX1 instanceL2_g11388(.CO(instanceL2_n_11046), .S(
    \instanceL2_prod_terms[7][5] [6]), .A(instanceL2_n_12518), .B(
    instanceL2_n_12515), .CI(instanceL2_n_11058));
  ADDFX1 instanceL2_g11389(.CO(instanceL2_n_12501), .S(
    \instanceL2_prod_terms[0][5][6] ), .A(instanceL2_n_12551), .B(
    instanceL2_n_12530), .CI(instanceL2_n_12504));
  MXI2XL instanceL2_g11390(.Y(\instanceL2_prod_terms[1][5] [10]), .A(
    layer1_out[52]), .B(instanceL2_n_12559), .S0(instanceL2_n_12503));
  AOI21X1 instanceL2_g11391(.Y(\instanceL2_prod_terms[2][5] [6]), .A0(
    layer1_out[50]), .A1(instanceL2_n_12507), .B0(instanceL2_n_12502));
  MX2XL instanceL2_g11392(.Y(\instanceL2_prod_terms[1][5] [9]), .A(
    layer1_out[51]), .B(instanceL2_n_12561), .S0(instanceL2_n_12505));
  ADDFX1 instanceL2_g11393(.CO(instanceL2_n_11058), .S(
    \instanceL2_prod_terms[7][5] [5]), .A(instanceL2_n_12540), .B(
    instanceL2_n_12517), .CI(instanceL2_n_12508));
  NOR2X1 instanceL2_g11394(.Y(\instanceL2_prod_terms[1][5] [11]), .A(
    instanceL2_n_12559), .B(instanceL2_n_12506));
  NOR2X1 instanceL2_g11395(.Y(instanceL2_n_12502), .A(layer1_out[50]), .B(
    instanceL2_n_12507));
  OR4X1 instanceL2_g11396(.Y(\instanceL2_prod_terms[9][5] [13]), .A(
    layer1_out[52]), .B(layer1_out[51]), .C(layer1_out[50]), .D(
    instanceL2_n_12507));
  AOI21X1 instanceL2_g11397(.Y(instanceL2_n_12503), .A0(layer1_out[51]), .A1(
    instanceL2_n_11075), .B0(instanceL2_n_11130));
  ADDFX1 instanceL2_g11398(.CO(instanceL2_n_12504), .S(
    \instanceL2_prod_terms[0][5][5] ), .A(instanceL2_n_12550), .B(
    instanceL2_n_12527), .CI(instanceL2_n_12510));
  NAND2BX1 instanceL2_g11399(.Y(instanceL2_n_12505), .AN(instanceL2_n_11075), .B(
    instanceL2_n_12538));
  AOI21X1 instanceL2_g11400(.Y(instanceL2_n_12506), .A0(layer1_out[51]), .A1(
    instanceL2_n_12509), .B0(instanceL2_n_11130));
  XNOR2X1 instanceL2_g11401(.Y(\instanceL2_prod_terms[1][5] [8]), .A(
    instanceL2_n_12529), .B(instanceL2_n_12509));
  OA21X1 instanceL2_g11402(.Y(instanceL2_n_11075), .A0(layer1_out[52]), .A1(
    layer1_out[50]), .B0(instanceL2_n_12509));
  OA21X1 instanceL2_g11403(.Y(\instanceL2_prod_terms[5][5] [6]), .A0(
    instanceL2_n_12557), .A1(instanceL2_n_12512), .B0(instanceL2_n_12507));
  ADDFX1 instanceL2_g11404(.CO(instanceL2_n_12508), .S(
    \instanceL2_prod_terms[7][5] [4]), .A(layer1_out[49]), .B(
    instanceL2_n_12542), .CI(\instanceL2_prod_terms[2][5] [2]));
  NAND2X1 instanceL2_g11405(.Y(instanceL2_n_12507), .A(instanceL2_n_12557), .B(
    instanceL2_n_12512));
  XNOR2X1 instanceL2_g11406(.Y(\instanceL2_prod_terms[1][5] [7]), .A(
    instanceL2_n_12530), .B(instanceL2_n_12511));
  OAI2BB1X1 instanceL2_g11407(.Y(instanceL2_n_12509), .A0N(instanceL2_n_12544),
     .A1N(instanceL2_n_12511), .B0(instanceL2_n_12545));
  ADDFX1 instanceL2_g11408(.CO(instanceL2_n_12510), .S(
    \instanceL2_prod_terms[0][5][4] ), .A(instanceL2_n_12549), .B(
    instanceL2_n_11132), .CI(instanceL2_n_12524));
  AOI21X1 instanceL2_g11409(.Y(\instanceL2_prod_terms[2][5] [4]), .A0(
    layer1_out[48]), .A1(instanceL2_n_12526), .B0(instanceL2_n_12512));
  OAI2BB1X1 instanceL2_g11410(.Y(instanceL2_n_12511), .A0N(instanceL2_n_12534),
     .A1N(instanceL2_n_12521), .B0(instanceL2_n_12537));
  XNOR2X1 instanceL2_g11411(.Y(\instanceL2_prod_terms[0][5][3] ), .A(
    instanceL2_n_12541), .B(instanceL2_n_12522));
  XNOR2X1 instanceL2_g11412(.Y(\instanceL2_prod_terms[1][5] [6]), .A(
    instanceL2_n_12527), .B(instanceL2_n_12521));
  ADDFX1 instanceL2_g11413(.CO(instanceL2_n_12514), .S(instanceL2_n_12513), .A(
    layer1_out[52]), .B(layer1_out[49]), .CI(instanceL2_n_12556));
  ADDFX1 instanceL2_g11414(.CO(instanceL2_n_12516), .S(instanceL2_n_12515), .A(
    layer1_out[48]), .B(layer1_out[51]), .CI(instanceL2_n_12555));
  ADDFX1 instanceL2_g11415(.CO(instanceL2_n_12518), .S(instanceL2_n_12517), .A(
    instanceL2_n_12558), .B(layer1_out[50]), .CI(layer1_out[47]));
  OAI21XL instanceL2_g11416(.Y(instanceL2_n_12519), .A0(instanceL2_n_12561), .A1(
    instanceL2_n_12548), .B0(instanceL2_n_12520));
  NOR2X1 instanceL2_g11417(.Y(instanceL2_n_12512), .A(layer1_out[48]), .B(
    instanceL2_n_12526));
  XNOR2X1 instanceL2_g11418(.Y(\instanceL2_prod_terms[1][5] [5]), .A(
    instanceL2_n_11132), .B(instanceL2_n_12523));
  XNOR2X1 instanceL2_g11419(.Y(instanceL2_n_11110), .A(instanceL2_n_12547), .B(
    instanceL2_n_12532));
  NAND2X1 instanceL2_g11420(.Y(instanceL2_n_12520), .A(instanceL2_n_12561), .B(
    instanceL2_n_12548));
  OAI211X1 instanceL2_g11421(.Y(instanceL2_n_12521), .A0(instanceL2_n_12539),
     .A1(instanceL2_n_12543), .B0(instanceL2_n_12546), .C0(instanceL2_n_12525));
  XNOR2X1 instanceL2_g11422(.Y(\instanceL2_prod_terms[1][5] [4]), .A(
    instanceL2_n_11165), .B(instanceL2_n_12528));
  MXI2XL instanceL2_g11423(.Y(instanceL2_n_12522), .A(instanceL2_n_12555), .B(
    layer1_out[47]), .S0(instanceL2_n_12528));
  NAND2X1 instanceL2_g11424(.Y(instanceL2_n_12523), .A(instanceL2_n_12539), .B(
    instanceL2_n_12525));
  OA21X1 instanceL2_g11425(.Y(\instanceL2_prod_terms[2][5] [3]), .A0(
    instanceL2_n_12555), .A1(instanceL2_n_12535), .B0(instanceL2_n_12526));
  AOI2BB1X1 instanceL2_g11426(.Y(instanceL2_n_12524), .A0N(layer1_out[47]), .A1N(
    instanceL2_n_12541), .B0(instanceL2_n_12528));
  NOR2BX1 instanceL2_g11427(.Y(\instanceL2_prod_terms[1][5] [3]), .AN(
    instanceL2_n_11165), .B(instanceL2_n_12541));
  OR2X1 instanceL2_g11428(.Y(instanceL2_n_12525), .A(instanceL2_n_12536), .B(
    instanceL2_n_11165));
  NOR2X1 instanceL2_g11429(.Y(instanceL2_n_11130), .A(instanceL2_n_12561), .B(
    instanceL2_n_12538));
  NAND2X1 instanceL2_g11430(.Y(instanceL2_n_12526), .A(instanceL2_n_12555), .B(
    instanceL2_n_12535));
  NAND2BX1 instanceL2_g11431(.Y(instanceL2_n_11132), .AN(instanceL2_n_12543), .B(
    instanceL2_n_12546));
  NAND2X1 instanceL2_g11432(.Y(instanceL2_n_12527), .A(instanceL2_n_12537), .B(
    instanceL2_n_12534));
  NOR2BX1 instanceL2_g11433(.Y(instanceL2_n_12528), .AN(instanceL2_n_12539), .B(
    instanceL2_n_12536));
  AOI21X1 instanceL2_g11434(.Y(\instanceL2_prod_terms[7][5] [3]), .A0(
    instanceL2_n_12554), .A1(instanceL2_n_12556), .B0(instanceL2_n_12542));
  OAI22X1 instanceL2_g11435(.Y(instanceL2_n_12531), .A0(layer1_out[50]), .A1(
    layer1_out[49]), .B0(instanceL2_n_12560), .B1(instanceL2_n_12557));
  OAI22X1 instanceL2_g11436(.Y(instanceL2_n_12532), .A0(layer1_out[52]), .A1(
    layer1_out[51]), .B0(instanceL2_n_12559), .B1(instanceL2_n_12561));
  AOI21X1 instanceL2_g11437(.Y(instanceL2_n_12533), .A0(instanceL2_n_12561), .A1(
    layer1_out[50]), .B0(instanceL2_n_12547));
  AOI21X1 instanceL2_g11438(.Y(instanceL2_n_12529), .A0(instanceL2_n_12559), .A1(
    layer1_out[50]), .B0(instanceL2_n_12548));
  NAND2X1 instanceL2_g11439(.Y(instanceL2_n_12530), .A(instanceL2_n_12545), .B(
    instanceL2_n_12544));
  OAI21X1 instanceL2_g11440(.Y(\instanceL2_prod_terms[2][5] [2]), .A0(
    instanceL2_n_12558), .A1(layer1_out[45]), .B0(instanceL2_n_12540));
  NAND2X1 instanceL2_g11441(.Y(instanceL2_n_12534), .A(instanceL2_n_12560), .B(
    instanceL2_n_12556));
  NOR2X1 instanceL2_g11442(.Y(instanceL2_n_12535), .A(layer1_out[46]), .B(
    layer1_out[45]));
  NOR2X1 instanceL2_g11443(.Y(instanceL2_n_12536), .A(layer1_out[46]), .B(
    layer1_out[48]));
  NAND2X1 instanceL2_g11444(.Y(instanceL2_n_12537), .A(layer1_out[50]), .B(
    layer1_out[48]));
  NAND2XL instanceL2_g11445(.Y(instanceL2_n_12538), .A(layer1_out[52]), .B(
    layer1_out[50]));
  NAND2X1 instanceL2_g11446(.Y(instanceL2_n_12539), .A(layer1_out[46]), .B(
    layer1_out[48]));
  NAND2X1 instanceL2_g11447(.Y(instanceL2_n_12540), .A(instanceL2_n_12558), .B(
    layer1_out[45]));
  NAND2X1 instanceL2_g11448(.Y(instanceL2_n_11165), .A(layer1_out[45]), .B(
    layer1_out[47]));
  NOR2X1 instanceL2_g11449(.Y(instanceL2_n_12541), .A(layer1_out[45]), .B(
    layer1_out[47]));
  NOR2X1 instanceL2_g11450(.Y(instanceL2_n_12542), .A(instanceL2_n_12554), .B(
    instanceL2_n_12556));
  NOR2XL instanceL2_g11451(.Y(instanceL2_n_12543), .A(layer1_out[49]), .B(
    layer1_out[47]));
  NAND2X1 instanceL2_g11452(.Y(instanceL2_n_12544), .A(instanceL2_n_12561), .B(
    instanceL2_n_12557));
  NAND2X1 instanceL2_g11453(.Y(instanceL2_n_12545), .A(layer1_out[51]), .B(
    layer1_out[49]));
  NOR2X1 instanceL2_g11454(.Y(instanceL2_n_12549), .A(layer1_out[46]), .B(
    instanceL2_n_12556));
  NAND2X1 instanceL2_g11455(.Y(instanceL2_n_12546), .A(layer1_out[47]), .B(
    layer1_out[49]));
  NOR2X1 instanceL2_g11456(.Y(instanceL2_n_12550), .A(layer1_out[47]), .B(
    instanceL2_n_12557));
  NOR2X1 instanceL2_g11457(.Y(instanceL2_n_12551), .A(layer1_out[48]), .B(
    instanceL2_n_12560));
  NOR2X1 instanceL2_g11458(.Y(instanceL2_n_12552), .A(instanceL2_n_12561), .B(
    layer1_out[49]));
  NOR2XL instanceL2_g11459(.Y(instanceL2_n_12553), .A(layer1_out[49]), .B(
    instanceL2_n_12560));
  NOR2X1 instanceL2_g11460(.Y(instanceL2_n_12547), .A(instanceL2_n_12561), .B(
    layer1_out[50]));
  NOR2X1 instanceL2_g11461(.Y(instanceL2_n_12548), .A(instanceL2_n_12559), .B(
    layer1_out[50]));
  INVX1 instanceL2_g11462(.Y(instanceL2_n_12554), .A(layer1_out[45]));
  INVX1 instanceL2_g11463(.Y(instanceL2_n_12555), .A(layer1_out[47]));
  INVX1 instanceL2_g11464(.Y(instanceL2_n_12556), .A(layer1_out[48]));
  INVX1 instanceL2_g11465(.Y(instanceL2_n_12557), .A(layer1_out[49]));
  INVX1 instanceL2_g11466(.Y(instanceL2_n_12558), .A(layer1_out[46]));
  INVX1 instanceL2_g11467(.Y(instanceL2_n_12559), .A(layer1_out[52]));
  INVX1 instanceL2_g11468(.Y(instanceL2_n_12560), .A(layer1_out[50]));
  INVX1 instanceL2_g11469(.Y(instanceL2_n_12561), .A(layer1_out[51]));
  OAI21X1 instanceL2_g11470(.Y(\instanceL2_prod_terms[2][5] [8]), .A0(
    instanceL2_n_12520), .A1(instanceL2_n_12507), .B0(instanceL2_n_12499));
  XNOR2X1 instanceL2_g11471(.Y(\instanceL2_prod_terms[0][17][9] ), .A(
    instanceL2_n_11102), .B(instanceL2_n_10995));
  ADDFX1 instanceL2_g11472(.CO(instanceL2_n_10995), .S(
    \instanceL2_prod_terms[0][17][8] ), .A(instanceL2_n_12637), .B(
    instanceL2_n_12599), .CI(instanceL2_n_10997));
  ADDFX1 instanceL2_g11473(.CO(instanceL2_n_10997), .S(
    \instanceL2_prod_terms[0][17][7] ), .A(instanceL2_n_12646), .B(
    instanceL2_n_12598), .CI(instanceL2_n_12563));
  XNOR2X1 instanceL2_g11474(.Y(\instanceL2_prod_terms[3][17] [10]), .A(
    layer1_out[161]), .B(instanceL2_n_12562));
  MXI2XL instanceL2_g11475(.Y(\instanceL2_prod_terms[3][17] [9]), .A(
    instanceL2_n_12639), .B(layer1_out[160]), .S0(instanceL2_n_12564));
  NAND2X1 instanceL2_g11476(.Y(\instanceL2_prod_terms[0][17][10] ), .A(
    instanceL2_n_12570), .B(instanceL2_n_12566));
  AOI22X1 instanceL2_g11477(.Y(instanceL2_n_12562), .A0(layer1_out[160]), .A1(
    instanceL2_n_12565), .B0(layer1_out[159]), .B1(instanceL2_n_12635));
  ADDFX1 instanceL2_g11478(.CO(instanceL2_n_12563), .S(
    \instanceL2_prod_terms[0][17][6] ), .A(instanceL2_n_12642), .B(
    instanceL2_n_12591), .CI(instanceL2_n_12569));
  NAND2BX1 instanceL2_g11479(.Y(instanceL2_n_12564), .AN(instanceL2_n_12565), .B(
    instanceL2_n_12625));
  OA21X1 instanceL2_g11480(.Y(\instanceL2_prod_terms[3][17] [11]), .A0(
    layer1_out[159]), .A1(instanceL2_n_12567), .B0(instanceL2_n_12635));
  XNOR2X1 instanceL2_g11481(.Y(\instanceL2_prod_terms[3][17] [8]), .A(
    instanceL2_n_12599), .B(instanceL2_n_12567));
  NOR2BX1 instanceL2_g11482(.Y(instanceL2_n_12565), .AN(instanceL2_n_12567), .B(
    instanceL2_n_12624));
  OAI21X1 instanceL2_g11483(.Y(\instanceL2_prod_terms[9][17] [9]), .A0(
    layer1_out[161]), .A1(instanceL2_n_12568), .B0(instanceL2_n_12566));
  XNOR2X1 instanceL2_g11484(.Y(\instanceL2_prod_terms[4][17] [7]), .A(
    layer1_out[160]), .B(instanceL2_n_12572));
  NAND2X1 instanceL2_g11485(.Y(instanceL2_n_12566), .A(layer1_out[161]), .B(
    instanceL2_n_12568));
  OAI21X1 instanceL2_g11486(.Y(instanceL2_n_12567), .A0(instanceL2_n_12605), .A1(
    instanceL2_n_11037), .B0(instanceL2_n_12608));
  XOR2XL instanceL2_g11487(.Y(\instanceL2_prod_terms[3][17] [7]), .A(
    instanceL2_n_12598), .B(instanceL2_n_11037));
  XNOR2X1 instanceL2_g11488(.Y(\instanceL2_prod_terms[4][17] [5]), .A(
    layer1_out[158]), .B(instanceL2_n_11047));
  ADDFX1 instanceL2_g11489(.CO(instanceL2_n_12569), .S(
    \instanceL2_prod_terms[0][17][5] ), .A(instanceL2_n_12643), .B(
    instanceL2_n_11108), .CI(instanceL2_n_12575));
  OAI2BB1X1 instanceL2_g11490(.Y(\instanceL2_prod_terms[4][17] [8]), .A0N(
    layer1_out[161]), .A1N(instanceL2_n_12571), .B0(instanceL2_n_12570));
  AOI21X1 instanceL2_g11491(.Y(instanceL2_n_12568), .A0(instanceL2_n_12644), .A1(
    instanceL2_n_12573), .B0(instanceL2_n_12635));
  OAI2BB1X1 instanceL2_g11492(.Y(\instanceL2_prod_terms[9][17] [10]), .A0N(
    layer1_out[161]), .A1N(instanceL2_n_12573), .B0(instanceL2_n_12634));
  XNOR2X1 instanceL2_g11493(.Y(\instanceL2_prod_terms[9][17] [8]), .A(
    instanceL2_n_12603), .B(instanceL2_n_12573));
  AOI21X1 instanceL2_g11494(.Y(\instanceL2_prod_terms[4][17] [6]), .A0(
    layer1_out[159]), .A1(instanceL2_n_12574), .B0(instanceL2_n_12572));
  OR2X1 instanceL2_g11495(.Y(instanceL2_n_12570), .A(layer1_out[161]), .B(
    instanceL2_n_12571));
  XNOR2X1 instanceL2_g11496(.Y(\instanceL2_prod_terms[3][17] [6]), .A(
    instanceL2_n_12591), .B(instanceL2_n_12578));
  XNOR2X1 instanceL2_g11497(.Y(\instanceL2_prod_terms[9][17] [7]), .A(
    instanceL2_n_12601), .B(instanceL2_n_12576));
  OA21X1 instanceL2_g11498(.Y(instanceL2_n_11037), .A0(instanceL2_n_12610), .A1(
    instanceL2_n_12577), .B0(instanceL2_n_12613));
  NOR2X1 instanceL2_g11499(.Y(instanceL2_n_12571), .A(instanceL2_n_12627), .B(
    instanceL2_n_12574));
  NOR2X1 instanceL2_g11500(.Y(instanceL2_n_12572), .A(layer1_out[159]), .B(
    instanceL2_n_12574));
  AOI21X1 instanceL2_g11501(.Y(\instanceL2_prod_terms[4][17] [4]), .A0(
    layer1_out[157]), .A1(instanceL2_n_12581), .B0(instanceL2_n_11047));
  OAI211X1 instanceL2_g11502(.Y(instanceL2_n_12573), .A0(instanceL2_n_12628),
     .A1(instanceL2_n_11062), .B0(instanceL2_n_12615), .C0(instanceL2_n_12629));
  ADDFX1 instanceL2_g11503(.CO(instanceL2_n_12575), .S(
    \instanceL2_prod_terms[0][17][4] ), .A(instanceL2_n_12645), .B(
    instanceL2_n_12590), .CI(instanceL2_n_12586));
  NAND2X1 instanceL2_g11504(.Y(instanceL2_n_12576), .A(instanceL2_n_12615), .B(
    instanceL2_n_11062));
  NOR2X1 instanceL2_g11505(.Y(instanceL2_n_11047), .A(layer1_out[157]), .B(
    instanceL2_n_12581));
  NAND2BX1 instanceL2_g11506(.Y(instanceL2_n_12574), .AN(instanceL2_n_12581), .B(
    instanceL2_n_12632));
  INVXL instanceL2_g11507(.Y(instanceL2_n_12577), .A(instanceL2_n_12578));
  XNOR2X1 instanceL2_g11508(.Y(\instanceL2_prod_terms[3][17] [5]), .A(
    instanceL2_n_11108), .B(instanceL2_n_12580));
  XNOR2X1 instanceL2_g11509(.Y(\instanceL2_prod_terms[9][17] [6]), .A(
    instanceL2_n_12594), .B(instanceL2_n_11069));
  OAI21X1 instanceL2_g11510(.Y(instanceL2_n_12578), .A0(instanceL2_n_12607), .A1(
    instanceL2_n_12579), .B0(instanceL2_n_12612));
  NAND2BX1 instanceL2_g11511(.Y(instanceL2_n_11062), .AN(instanceL2_n_12614), .B(
    instanceL2_n_11069));
  XNOR2X1 instanceL2_g11512(.Y(\instanceL2_prod_terms[0][17][3] ), .A(
    instanceL2_n_12621), .B(instanceL2_n_12584));
  XNOR2X1 instanceL2_g11513(.Y(\instanceL2_prod_terms[9][17] [5]), .A(
    instanceL2_n_12604), .B(instanceL2_n_12583));
  INVX1 instanceL2_g11514(.Y(instanceL2_n_12579), .A(instanceL2_n_12580));
  AOI21X1 instanceL2_g11515(.Y(\instanceL2_prod_terms[4][17] [3]), .A0(
    layer1_out[156]), .A1(instanceL2_n_12597), .B0(instanceL2_n_12582));
  OAI21X1 instanceL2_g11516(.Y(instanceL2_n_12580), .A0(instanceL2_n_12606), .A1(
    instanceL2_n_12587), .B0(instanceL2_n_12609));
  XOR2XL instanceL2_g11517(.Y(\instanceL2_prod_terms[3][17] [4]), .A(
    instanceL2_n_12590), .B(instanceL2_n_12587));
  OAI211X1 instanceL2_g11518(.Y(instanceL2_n_11069), .A0(instanceL2_n_12632),
     .A1(instanceL2_n_12585), .B0(instanceL2_n_12616), .C0(instanceL2_n_12611));
  INVX1 instanceL2_g11519(.Y(instanceL2_n_12581), .A(instanceL2_n_12582));
  NAND2X1 instanceL2_g11520(.Y(instanceL2_n_12583), .A(instanceL2_n_12616), .B(
    instanceL2_n_12585));
  NOR2X1 instanceL2_g11521(.Y(instanceL2_n_12582), .A(layer1_out[156]), .B(
    instanceL2_n_12597));
  XNOR2X1 instanceL2_g11522(.Y(\instanceL2_prod_terms[9][17] [4]), .A(
    instanceL2_n_12595), .B(instanceL2_n_12589));
  XNOR2X1 instanceL2_g11523(.Y(\instanceL2_prod_terms[3][17] [3]), .A(
    instanceL2_n_12620), .B(instanceL2_n_12588));
  XNOR2X1 instanceL2_g11524(.Y(instanceL2_n_12584), .A(layer1_out[155]), .B(
    instanceL2_n_12600));
  OAI22X1 instanceL2_g11525(.Y(\instanceL2_prod_terms[9][17] [2]), .A0(
    instanceL2_n_12623), .A1(instanceL2_n_12596), .B0(instanceL2_n_12633), .B1(
    instanceL2_n_12617));
  NAND2BX1 instanceL2_g11526(.Y(instanceL2_n_12585), .AN(instanceL2_n_12630), .B(
    instanceL2_n_12589));
  AOI2BB1X1 instanceL2_g11527(.Y(instanceL2_n_12586), .A0N(layer1_out[155]),
     .A1N(instanceL2_n_12621), .B0(instanceL2_n_12588));
  OR4X1 instanceL2_g11528(.Y(\instanceL2_prod_terms[4][17] [13]), .A(
    layer1_out[154]), .B(instanceL2_n_12622), .C(instanceL2_n_12644), .D(
    instanceL2_n_12592));
  XNOR2X1 instanceL2_g11529(.Y(\instanceL2_prod_terms[9][17] [3]), .A(
    instanceL2_n_12602), .B(instanceL2_n_12596));
  OAI22X1 instanceL2_g11530(.Y(instanceL2_n_12587), .A0(layer1_out[154]), .A1(
    instanceL2_n_12593), .B0(layer1_out[156]), .B1(instanceL2_n_12619));
  INVX1 instanceL2_g11531(.Y(instanceL2_n_12588), .A(instanceL2_n_12600));
  OA21X1 instanceL2_g11532(.Y(\instanceL2_prod_terms[4][17] [2]), .A0(
    instanceL2_n_12638), .A1(instanceL2_n_12618), .B0(instanceL2_n_12597));
  OAI221X1 instanceL2_g10078(.Y(instanceL2_n_11102), .A0(layer1_out[159]), .A1(
    instanceL2_n_12636), .B0(layer1_out[161]), .B1(instanceL2_n_12639), .C0(
    instanceL2_n_12629));
  OAI211X1 instanceL2_g10079(.Y(instanceL2_n_12589), .A0(instanceL2_n_12626),
     .A1(instanceL2_n_12633), .B0(instanceL2_n_12617), .C0(instanceL2_n_12631));
  NOR2BX1 instanceL2_g10080(.Y(\instanceL2_prod_terms[4][17] [1]), .AN(
    instanceL2_n_12633), .B(instanceL2_n_12618));
  NOR2X1 instanceL2_g10081(.Y(\instanceL2_prod_terms[0][17][2] ), .A(
    instanceL2_n_12619), .B(instanceL2_n_12621));
  NAND2XL instanceL2_g10082(.Y(instanceL2_n_12592), .A(instanceL2_n_12614), .B(
    instanceL2_n_12630));
  NOR2BX1 instanceL2_g10083(.Y(instanceL2_n_12593), .AN(instanceL2_n_12640), .B(
    instanceL2_n_12631));
  NAND2BXL instanceL2_g10084(.Y(instanceL2_n_12594), .AN(instanceL2_n_12614), .B(
    instanceL2_n_12615));
  NAND2BXL instanceL2_g10085(.Y(instanceL2_n_12595), .AN(instanceL2_n_12630), .B(
    instanceL2_n_12616));
  NAND2BX1 instanceL2_g10086(.Y(instanceL2_n_12590), .AN(instanceL2_n_12606), .B(
    instanceL2_n_12609));
  NAND2BX1 instanceL2_g10087(.Y(instanceL2_n_11108), .AN(instanceL2_n_12607), .B(
    instanceL2_n_12612));
  NAND2BX1 instanceL2_g10088(.Y(instanceL2_n_12591), .AN(instanceL2_n_12610), .B(
    instanceL2_n_12613));
  NAND2XL instanceL2_g10089(.Y(instanceL2_n_12601), .A(instanceL2_n_12629), .B(
    instanceL2_n_12627));
  NAND2BX1 instanceL2_g10090(.Y(instanceL2_n_12602), .AN(instanceL2_n_12626), .B(
    instanceL2_n_12631));
  NAND2XL instanceL2_g10091(.Y(instanceL2_n_12603), .A(instanceL2_n_12634), .B(
    instanceL2_n_12644));
  NAND2BX1 instanceL2_g10092(.Y(instanceL2_n_12604), .AN(instanceL2_n_12632), .B(
    instanceL2_n_12611));
  NAND2X1 instanceL2_g10093(.Y(instanceL2_n_12596), .A(instanceL2_n_12633), .B(
    instanceL2_n_12617));
  NAND2X1 instanceL2_g10094(.Y(instanceL2_n_12597), .A(instanceL2_n_12638), .B(
    instanceL2_n_12618));
  NAND2BX1 instanceL2_g10095(.Y(instanceL2_n_12598), .AN(instanceL2_n_12605), .B(
    instanceL2_n_12608));
  NAND2BX1 instanceL2_g10096(.Y(instanceL2_n_12599), .AN(instanceL2_n_12624), .B(
    instanceL2_n_12625));
  XNOR2X1 instanceL2_g10097(.Y(instanceL2_n_12600), .A(layer1_out[156]), .B(
    layer1_out[154]));
  INVX1 instanceL2_g10098(.Y(instanceL2_n_12619), .A(instanceL2_n_12620));
  INVXL instanceL2_g10099(.Y(instanceL2_n_12622), .A(instanceL2_n_12621));
  NOR2XL instanceL2_g10100(.Y(instanceL2_n_12623), .A(layer1_out[154]), .B(
    layer1_out[155]));
  NOR2XL instanceL2_g10101(.Y(instanceL2_n_12605), .A(layer1_out[160]), .B(
    layer1_out[158]));
  NOR2XL instanceL2_g10102(.Y(instanceL2_n_12606), .A(layer1_out[157]), .B(
    layer1_out[155]));
  NOR2X1 instanceL2_g10103(.Y(instanceL2_n_12607), .A(layer1_out[158]), .B(
    layer1_out[156]));
  NAND2X1 instanceL2_g10104(.Y(instanceL2_n_12608), .A(layer1_out[160]), .B(
    layer1_out[158]));
  NAND2X1 instanceL2_g10105(.Y(instanceL2_n_12609), .A(layer1_out[155]), .B(
    layer1_out[157]));
  NOR2XL instanceL2_g10106(.Y(instanceL2_n_12610), .A(layer1_out[159]), .B(
    layer1_out[157]));
  NAND2X1 instanceL2_g10107(.Y(instanceL2_n_12611), .A(layer1_out[158]), .B(
    layer1_out[157]));
  NAND2X1 instanceL2_g10108(.Y(instanceL2_n_12612), .A(layer1_out[158]), .B(
    layer1_out[156]));
  NAND2XL instanceL2_g10109(.Y(instanceL2_n_12613), .A(layer1_out[159]), .B(
    layer1_out[157]));
  NOR2XL instanceL2_g11533(.Y(instanceL2_n_12614), .A(layer1_out[159]), .B(
    layer1_out[158]));
  NAND2X1 instanceL2_g11534(.Y(instanceL2_n_12615), .A(layer1_out[158]), .B(
    layer1_out[159]));
  NAND2X1 instanceL2_g11535(.Y(instanceL2_n_12616), .A(layer1_out[157]), .B(
    layer1_out[156]));
  NAND2XL instanceL2_g11536(.Y(instanceL2_n_12617), .A(layer1_out[155]), .B(
    layer1_out[154]));
  NOR2X1 instanceL2_g11537(.Y(instanceL2_n_12618), .A(instanceL2_n_12640), .B(
    layer1_out[154]));
  NAND2XL instanceL2_g11538(.Y(instanceL2_n_12620), .A(instanceL2_n_12640), .B(
    layer1_out[155]));
  NOR2X1 instanceL2_g11539(.Y(instanceL2_n_12621), .A(instanceL2_n_12640), .B(
    layer1_out[155]));
  INVX1 instanceL2_g11540(.Y(instanceL2_n_12627), .A(instanceL2_n_12628));
  INVX1 instanceL2_g11541(.Y(instanceL2_n_12635), .A(instanceL2_n_12634));
  NAND2XL instanceL2_g11542(.Y(instanceL2_n_12636), .A(layer1_out[161]), .B(
    instanceL2_n_12639));
  NOR2X1 instanceL2_g11543(.Y(instanceL2_n_12637), .A(layer1_out[158]), .B(
    instanceL2_n_12639));
  NOR2XL instanceL2_g11544(.Y(instanceL2_n_12624), .A(layer1_out[161]), .B(
    layer1_out[159]));
  NAND2X1 instanceL2_g11545(.Y(instanceL2_n_12625), .A(layer1_out[161]), .B(
    layer1_out[159]));
  NOR2X1 instanceL2_g11546(.Y(instanceL2_n_12626), .A(layer1_out[155]), .B(
    layer1_out[156]));
  NOR2X1 instanceL2_g11547(.Y(instanceL2_n_12628), .A(layer1_out[160]), .B(
    layer1_out[159]));
  NAND2XL instanceL2_g11548(.Y(instanceL2_n_12629), .A(layer1_out[160]), .B(
    layer1_out[159]));
  NOR2XL instanceL2_g11549(.Y(instanceL2_n_12630), .A(layer1_out[157]), .B(
    layer1_out[156]));
  NAND2XL instanceL2_g11550(.Y(instanceL2_n_12631), .A(layer1_out[155]), .B(
    layer1_out[156]));
  NOR2X1 instanceL2_g11551(.Y(instanceL2_n_12632), .A(layer1_out[158]), .B(
    layer1_out[157]));
  NAND2X1 instanceL2_g11552(.Y(instanceL2_n_12633), .A(instanceL2_n_12640), .B(
    layer1_out[154]));
  NAND2XL instanceL2_g11553(.Y(instanceL2_n_12634), .A(layer1_out[161]), .B(
    layer1_out[160]));
  INVX1 instanceL2_g11554(.Y(instanceL2_n_12638), .A(layer1_out[155]));
  INVX1 instanceL2_g11555(.Y(instanceL2_n_12639), .A(layer1_out[160]));
  INVX1 instanceL2_drc_bufs(.Y(instanceL2_n_12640), .A(instanceL2_n_12641));
  INVX1 instanceL2_drc_bufs10144(.Y(instanceL2_n_12641), .A(layer1_out[153]));
  NOR2BX1 instanceL2_g11556(.Y(instanceL2_n_12642), .AN(layer1_out[158]), .B(
    layer1_out[156]));
  NOR2BX1 instanceL2_g11557(.Y(instanceL2_n_12643), .AN(layer1_out[157]), .B(
    layer1_out[155]));
  NAND2BX1 instanceL2_g11558(.Y(instanceL2_n_12644), .AN(layer1_out[161]), .B(
    instanceL2_n_12639));
  NOR2BX1 instanceL2_g11559(.Y(instanceL2_n_12645), .AN(layer1_out[156]), .B(
    layer1_out[154]));
  NOR2BX1 instanceL2_g11560(.Y(instanceL2_n_12646), .AN(layer1_out[159]), .B(
    layer1_out[157]));
endmodule

