//
// Conformal-LEC: Version 24.10-s400 (28-Apr-2025) (64 bit executable)
//
module VDW_WMUX2 (Z, A, B, S);
// conformal library_module
output [1:0] Z;
input [1:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_ADD_2_1_0_CIM(SUM, A, B);
// conformal library_module
input   [1:0] A;
input   [1:0] B;
output  [1:0] SUM;
wire   [1:0] SUM;
wire   [1:0] B;
wire   [1:0] A;
  xor U$1(SUM[1], A[1], A[0]);
  not U$2(SUM[0], A[0]);
endmodule

module VDW_LT_u2_CIM(Z, A, B);
// conformal library_module
output Z;
input   [1:0] A;
input   [1:0] B;
wire  Z;
wire   [1:0] B;
wire   [1:0] A;
  nand U$1(Z, A[0], A[1]);
endmodule

module VDW_WMUX5 (Z, A, B, S);
// conformal library_module
output [4:0] Z;
input [4:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_ADD_10_1_0(SUM, A, B);
input   [9:0] A;
input   [9:0] B;
output  [9:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42;
wire   [9:0] SUM;
wire   [9:0] B;
wire   [9:0] A;
  xor U$1(SUM[9], N$2, N$1);
  xor U$2(N$2, A[9], B[9]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[8], N$6);
  and U$5(N$4, B[8], N$6);
  and U$6(N$5, A[8], B[8]);
  xor U$7(SUM[8], N$7, N$6);
  xor U$8(N$7, A[8], B[8]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[7], N$11);
  and U$11(N$9, B[7], N$11);
  and U$12(N$10, A[7], B[7]);
  xor U$13(SUM[7], N$12, N$11);
  xor U$14(N$12, A[7], B[7]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[6], N$16);
  and U$17(N$14, B[6], N$16);
  and U$18(N$15, A[6], B[6]);
  xor U$19(SUM[6], N$17, N$16);
  xor U$20(N$17, A[6], B[6]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[5], N$21);
  and U$23(N$19, B[5], N$21);
  and U$24(N$20, A[5], B[5]);
  xor U$25(SUM[5], N$22, N$21);
  xor U$26(N$22, A[5], B[5]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[4], N$26);
  and U$29(N$24, B[4], N$26);
  and U$30(N$25, A[4], B[4]);
  xor U$31(SUM[4], N$27, N$26);
  xor U$32(N$27, A[4], B[4]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[3], N$31);
  and U$35(N$29, B[3], N$31);
  and U$36(N$30, A[3], B[3]);
  xor U$37(SUM[3], N$32, N$31);
  xor U$38(N$32, A[3], B[3]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[2], N$36);
  and U$41(N$34, B[2], N$36);
  and U$42(N$35, A[2], B[2]);
  xor U$43(SUM[2], N$37, N$36);
  xor U$44(N$37, A[2], B[2]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[1], N$41);
  and U$47(N$39, B[1], N$41);
  and U$48(N$40, A[1], B[1]);
  xor U$49(SUM[1], N$42, N$41);
  xor U$50(N$42, A[1], B[1]);
  and U$51(N$41, A[0], B[0]);
  xor U$52(SUM[0], A[0], B[0]);
endmodule

module VDW_WMUX256 (Z, A, B, S);
// conformal library_module
output [255:0] Z;
input [255:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX9 (Z, A, B, S);
// conformal library_module
output [8:0] Z;
input [8:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module ReLU_10bit(in_data, out_data);
input   [9:0] in_data;
output  [8:0] out_data;
wire  n196;
wire   [8:0] out_data;
wire   [9:0] in_data;
  VDW_WMUX9 U$1(.Z({ out_data[8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ in_data[8:0] }), .S(n196));
  not U$2(n196, in_data[9]);
endmodule

module VDW_ADD_6_1_0(SUM, A, B);
input   [5:0] A;
input   [5:0] B;
output  [5:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22;
wire   [5:0] SUM;
wire   [5:0] B;
wire   [5:0] A;
  xor U$1(SUM[5], N$2, N$1);
  xor U$2(N$2, A[5], B[5]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[4], N$6);
  and U$5(N$4, B[4], N$6);
  and U$6(N$5, A[4], B[4]);
  xor U$7(SUM[4], N$7, N$6);
  xor U$8(N$7, A[4], B[4]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[3], N$11);
  and U$11(N$9, B[3], N$11);
  and U$12(N$10, A[3], B[3]);
  xor U$13(SUM[3], N$12, N$11);
  xor U$14(N$12, A[3], B[3]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[2], N$16);
  and U$17(N$14, B[2], N$16);
  and U$18(N$15, A[2], B[2]);
  xor U$19(SUM[2], N$17, N$16);
  xor U$20(N$17, A[2], B[2]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[1], N$21);
  and U$23(N$19, B[1], N$21);
  and U$24(N$20, A[1], B[1]);
  xor U$25(SUM[1], N$22, N$21);
  xor U$26(N$22, A[1], B[1]);
  and U$27(N$21, A[0], B[0]);
  xor U$28(SUM[0], A[0], B[0]);
endmodule

module adder_5to6(a, b, sum);
input   [4:0] a;
input   [4:0] b;
output  [5:0] sum;
wire   [5:0] sum;
wire   [4:0] b;
wire   [4:0] a;
  VDW_ADD_6_1_0 add_6_20(.SUM({ sum[5:0] }), .A({a[4],  a[4:0] }), .B({b[4],  b[4:0] }));
endmodule

module VDW_ADD_7_1_0(SUM, A, B);
input   [6:0] A;
input   [6:0] B;
output  [6:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27;
wire   [6:0] SUM;
wire   [6:0] B;
wire   [6:0] A;
  xor U$1(SUM[6], N$2, N$1);
  xor U$2(N$2, A[6], B[6]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[5], N$6);
  and U$5(N$4, B[5], N$6);
  and U$6(N$5, A[5], B[5]);
  xor U$7(SUM[5], N$7, N$6);
  xor U$8(N$7, A[5], B[5]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[4], N$11);
  and U$11(N$9, B[4], N$11);
  and U$12(N$10, A[4], B[4]);
  xor U$13(SUM[4], N$12, N$11);
  xor U$14(N$12, A[4], B[4]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[3], N$16);
  and U$17(N$14, B[3], N$16);
  and U$18(N$15, A[3], B[3]);
  xor U$19(SUM[3], N$17, N$16);
  xor U$20(N$17, A[3], B[3]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[2], N$21);
  and U$23(N$19, B[2], N$21);
  and U$24(N$20, A[2], B[2]);
  xor U$25(SUM[2], N$22, N$21);
  xor U$26(N$22, A[2], B[2]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[1], N$26);
  and U$29(N$24, B[1], N$26);
  and U$30(N$25, A[1], B[1]);
  xor U$31(SUM[1], N$27, N$26);
  xor U$32(N$27, A[1], B[1]);
  and U$33(N$26, A[0], B[0]);
  xor U$34(SUM[0], A[0], B[0]);
endmodule

module adder_6to7(a, b, sum);
input   [5:0] a;
input   [5:0] b;
output  [6:0] sum;
wire   [6:0] sum;
wire   [5:0] b;
wire   [5:0] a;
  VDW_ADD_7_1_0 add_14_20(.SUM({ sum[6:0] }), .A({a[5],  a[5:0] }), .B({b[5],  b[5:0] }));
endmodule

module VDW_ADD_8_1_0(SUM, A, B);
input   [7:0] A;
input   [7:0] B;
output  [7:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32;
wire   [7:0] SUM;
wire   [7:0] B;
wire   [7:0] A;
  xor U$1(SUM[7], N$2, N$1);
  xor U$2(N$2, A[7], B[7]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[6], N$6);
  and U$5(N$4, B[6], N$6);
  and U$6(N$5, A[6], B[6]);
  xor U$7(SUM[6], N$7, N$6);
  xor U$8(N$7, A[6], B[6]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[5], N$11);
  and U$11(N$9, B[5], N$11);
  and U$12(N$10, A[5], B[5]);
  xor U$13(SUM[5], N$12, N$11);
  xor U$14(N$12, A[5], B[5]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[4], N$16);
  and U$17(N$14, B[4], N$16);
  and U$18(N$15, A[4], B[4]);
  xor U$19(SUM[4], N$17, N$16);
  xor U$20(N$17, A[4], B[4]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[3], N$21);
  and U$23(N$19, B[3], N$21);
  and U$24(N$20, A[3], B[3]);
  xor U$25(SUM[3], N$22, N$21);
  xor U$26(N$22, A[3], B[3]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[2], N$26);
  and U$29(N$24, B[2], N$26);
  and U$30(N$25, A[2], B[2]);
  xor U$31(SUM[2], N$27, N$26);
  xor U$32(N$27, A[2], B[2]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[1], N$31);
  and U$35(N$29, B[1], N$31);
  and U$36(N$30, A[1], B[1]);
  xor U$37(SUM[1], N$32, N$31);
  xor U$38(N$32, A[1], B[1]);
  and U$39(N$31, A[0], B[0]);
  xor U$40(SUM[0], A[0], B[0]);
endmodule

module adder_7to8(a, b, sum);
input   [6:0] a;
input   [6:0] b;
output  [7:0] sum;
wire   [7:0] sum;
wire   [6:0] b;
wire   [6:0] a;
  VDW_ADD_8_1_0 add_22_20(.SUM({ sum[7:0] }), .A({a[6],  a[6:0] }), .B({b[6],  b[6:0] }));
endmodule

module VDW_ADD_9_1_0(SUM, A, B);
input   [8:0] A;
input   [8:0] B;
output  [8:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37;
wire   [8:0] SUM;
wire   [8:0] B;
wire   [8:0] A;
  xor U$1(SUM[8], N$2, N$1);
  xor U$2(N$2, A[8], B[8]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[7], N$6);
  and U$5(N$4, B[7], N$6);
  and U$6(N$5, A[7], B[7]);
  xor U$7(SUM[7], N$7, N$6);
  xor U$8(N$7, A[7], B[7]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[6], N$11);
  and U$11(N$9, B[6], N$11);
  and U$12(N$10, A[6], B[6]);
  xor U$13(SUM[6], N$12, N$11);
  xor U$14(N$12, A[6], B[6]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[5], N$16);
  and U$17(N$14, B[5], N$16);
  and U$18(N$15, A[5], B[5]);
  xor U$19(SUM[5], N$17, N$16);
  xor U$20(N$17, A[5], B[5]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[4], N$21);
  and U$23(N$19, B[4], N$21);
  and U$24(N$20, A[4], B[4]);
  xor U$25(SUM[4], N$22, N$21);
  xor U$26(N$22, A[4], B[4]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[3], N$26);
  and U$29(N$24, B[3], N$26);
  and U$30(N$25, A[3], B[3]);
  xor U$31(SUM[3], N$27, N$26);
  xor U$32(N$27, A[3], B[3]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[2], N$31);
  and U$35(N$29, B[2], N$31);
  and U$36(N$30, A[2], B[2]);
  xor U$37(SUM[2], N$32, N$31);
  xor U$38(N$32, A[2], B[2]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[1], N$36);
  and U$41(N$34, B[1], N$36);
  and U$42(N$35, A[1], B[1]);
  xor U$43(SUM[1], N$37, N$36);
  xor U$44(N$37, A[1], B[1]);
  and U$45(N$36, A[0], B[0]);
  xor U$46(SUM[0], A[0], B[0]);
endmodule

module adder_8to9(a, b, sum);
input   [7:0] a;
input   [7:0] b;
output  [8:0] sum;
wire   [8:0] sum;
wire   [7:0] b;
wire   [7:0] a;
  VDW_ADD_9_1_0 add_30_20(.SUM({ sum[8:0] }), .A({a[7],  a[7:0] }), .B({b[7],  b[7:0] }));
endmodule

module adder_9to10(a, b, sum);
input   [8:0] a;
input   [8:0] b;
output  [9:0] sum;
wire   [9:0] sum;
wire   [8:0] b;
wire   [8:0] a;
  VDW_ADD_10_1_0 add_38_20(.SUM({ sum[9:0] }), .A({a[8],  a[8:0] }), .B({b[8],  b[8:0] }));
endmodule

module VDW_ADD_11_1_0(SUM, A, B);
input   [10:0] A;
input   [10:0] B;
output  [10:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47;
wire   [10:0] SUM;
wire   [10:0] B;
wire   [10:0] A;
  xor U$1(SUM[10], N$2, N$1);
  xor U$2(N$2, A[10], B[10]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[9], N$6);
  and U$5(N$4, B[9], N$6);
  and U$6(N$5, A[9], B[9]);
  xor U$7(SUM[9], N$7, N$6);
  xor U$8(N$7, A[9], B[9]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[8], N$11);
  and U$11(N$9, B[8], N$11);
  and U$12(N$10, A[8], B[8]);
  xor U$13(SUM[8], N$12, N$11);
  xor U$14(N$12, A[8], B[8]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[7], N$16);
  and U$17(N$14, B[7], N$16);
  and U$18(N$15, A[7], B[7]);
  xor U$19(SUM[7], N$17, N$16);
  xor U$20(N$17, A[7], B[7]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[6], N$21);
  and U$23(N$19, B[6], N$21);
  and U$24(N$20, A[6], B[6]);
  xor U$25(SUM[6], N$22, N$21);
  xor U$26(N$22, A[6], B[6]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[5], N$26);
  and U$29(N$24, B[5], N$26);
  and U$30(N$25, A[5], B[5]);
  xor U$31(SUM[5], N$27, N$26);
  xor U$32(N$27, A[5], B[5]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[4], N$31);
  and U$35(N$29, B[4], N$31);
  and U$36(N$30, A[4], B[4]);
  xor U$37(SUM[4], N$32, N$31);
  xor U$38(N$32, A[4], B[4]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[3], N$36);
  and U$41(N$34, B[3], N$36);
  and U$42(N$35, A[3], B[3]);
  xor U$43(SUM[3], N$37, N$36);
  xor U$44(N$37, A[3], B[3]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[2], N$41);
  and U$47(N$39, B[2], N$41);
  and U$48(N$40, A[2], B[2]);
  xor U$49(SUM[2], N$42, N$41);
  xor U$50(N$42, A[2], B[2]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[1], N$46);
  and U$53(N$44, B[1], N$46);
  and U$54(N$45, A[1], B[1]);
  xor U$55(SUM[1], N$47, N$46);
  xor U$56(N$47, A[1], B[1]);
  and U$57(N$46, A[0], B[0]);
  xor U$58(SUM[0], A[0], B[0]);
endmodule

module adder_10to10(a, b, sum);
input   [9:0] a;
input   [9:0] b;
output  [9:0] sum;
wire   [10:0] result;
wire   [9:0] sum;
wire   [9:0] b;
wire   [9:0] a;
  VDW_ADD_11_1_0 add_47_23(.SUM({dummy$0,  result[9:0] }), .A({a[9],  a[9:0] }), .B({b[9],  b[9:0] }));
  assign sum[0] = result[0];
  assign sum[1] = result[1];
  assign sum[2] = result[2];
  assign sum[3] = result[3];
  assign sum[4] = result[4];
  assign sum[5] = result[5];
  assign sum[6] = result[6];
  assign sum[7] = result[7];
  assign sum[8] = result[8];
  assign sum[9] = result[9];
endmodule

module layer1(clk, rst_n, updown, in, out);
input  clk, rst_n, updown;
input   [0:127] in;
output  [179:0] out;
wire  n5413, updown, rst_n, clk;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76, N$77, N$78, N$79, N$80, N$81, N$82, N$83, N$84, N$85, N$86, 
    N$87, N$88, N$89, N$90, N$91, N$92, N$93, N$94, N$95, N$96, N$97, N$98, 
    N$99, N$100, N$101, N$102, N$103, N$104, N$105, N$106, N$107, N$108, N$109, 
    N$110, N$111, N$112, N$113, N$114, N$115, N$116, N$117, N$118, N$119, 
    N$120, N$121, N$122, N$123, N$124, N$125, N$126, N$127, N$128, N$129, 
    N$130, N$131, N$132, N$133, N$134, N$135, N$136, N$137, N$138, N$139, 
    N$140, N$141, N$142, N$143, N$144, N$145, N$146, N$147, N$148, N$149, 
    N$150, N$151, N$152, N$153, N$154, N$155, N$156, N$157, N$158, N$159, 
    N$160, N$161, N$162, N$163, N$164, N$165, N$166, N$167, N$168, N$169, 
    N$170, N$171, N$172, N$173, N$174, N$175, N$176, N$177, N$178, N$179, 
    N$180, N$181, N$182, N$183, N$184, N$185, N$186, N$187, N$188, N$189, 
    N$190, N$191, N$192, N$193, N$194, N$195, N$196, N$197, N$198, N$199, 
    N$200, N$201, N$202, N$203, N$204, N$205, N$206, N$207, N$208, N$209, 
    N$210, N$211, N$212, N$213, N$214, N$215, N$216, N$217, N$218, N$219, 
    N$220, N$221, N$222, N$223, N$224, N$225, N$226, N$227, N$228, N$229, 
    N$230, N$231, N$232, N$233, N$234, N$235, N$236, N$237, N$238, N$239, 
    N$240, N$241, N$242, N$243, N$244, N$245, N$246, N$247, N$248, N$249, 
    N$250, N$251, N$252, N$253, N$254, N$255, N$256, N$257, N$258, N$259, 
    N$260, N$261, N$262, N$263, N$264, N$265;
wire   [255:0] n5418;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[19].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[18].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[17].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[16].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[15].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[14].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[13].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[12].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[11].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[10].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[9].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[8].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[7].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[6].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[5].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[4].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[3].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[2].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[1].product_terms[255] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[0] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[1] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[2] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[3] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[4] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[5] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[6] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[7] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[8] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[9] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[10] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[11] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[12] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[13] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[14] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[15] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[16] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[17] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[18] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[19] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[20] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[21] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[22] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[23] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[24] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[25] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[26] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[27] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[28] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[29] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[30] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[31] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[32] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[33] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[34] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[35] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[36] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[37] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[38] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[39] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[40] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[41] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[42] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[43] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[44] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[45] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[46] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[47] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[48] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[49] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[50] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[51] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[52] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[53] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[54] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[55] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[56] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[57] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[58] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[59] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[60] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[61] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[62] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[63] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[64] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[65] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[66] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[67] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[68] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[69] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[70] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[71] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[72] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[73] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[74] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[75] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[76] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[77] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[78] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[79] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[80] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[81] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[82] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[83] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[84] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[85] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[86] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[87] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[88] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[89] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[90] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[91] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[92] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[93] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[94] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[95] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[96] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[97] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[98] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[99] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[100] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[101] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[102] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[103] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[104] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[105] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[106] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[107] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[108] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[109] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[110] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[111] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[112] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[113] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[114] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[115] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[116] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[117] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[118] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[119] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[120] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[121] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[122] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[123] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[124] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[125] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[126] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[127] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[128] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[129] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[130] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[131] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[132] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[133] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[134] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[135] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[136] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[137] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[138] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[139] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[140] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[141] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[142] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[143] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[144] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[145] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[146] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[147] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[148] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[149] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[150] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[151] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[152] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[153] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[154] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[155] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[156] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[157] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[158] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[159] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[160] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[161] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[162] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[163] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[164] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[165] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[166] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[167] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[168] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[169] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[170] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[171] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[172] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[173] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[174] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[175] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[176] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[177] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[178] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[179] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[180] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[181] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[182] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[183] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[184] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[185] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[186] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[187] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[188] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[189] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[190] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[191] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[192] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[193] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[194] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[195] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[196] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[197] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[198] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[199] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[200] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[201] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[202] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[203] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[204] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[205] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[206] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[207] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[208] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[209] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[210] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[211] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[212] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[213] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[214] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[215] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[216] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[217] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[218] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[219] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[220] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[221] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[222] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[223] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[224] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[225] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[226] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[227] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[228] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[229] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[230] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[231] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[232] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[233] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[234] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[235] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[236] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[237] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[238] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[239] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[240] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[241] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[242] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[243] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[244] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[245] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[246] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[247] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[248] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[249] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[250] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[251] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[252] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[253] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[254] ;
wire   [4:0] \dot_product_and_ReLU[0].product_terms[255] ;
wire   [8:0] \out_sig[0] ;
wire   [8:0] \out_sig[1] ;
wire   [8:0] \out_sig[2] ;
wire   [8:0] \out_sig[3] ;
wire   [8:0] \out_sig[4] ;
wire   [8:0] \out_sig[5] ;
wire   [8:0] \out_sig[6] ;
wire   [8:0] \out_sig[7] ;
wire   [8:0] \out_sig[8] ;
wire   [8:0] \out_sig[9] ;
wire   [8:0] \out_sig[10] ;
wire   [8:0] \out_sig[11] ;
wire   [8:0] \out_sig[12] ;
wire   [8:0] \out_sig[13] ;
wire   [8:0] \out_sig[14] ;
wire   [8:0] \out_sig[15] ;
wire   [8:0] \out_sig[16] ;
wire   [8:0] \out_sig[17] ;
wire   [8:0] \out_sig[18] ;
wire   [8:0] \out_sig[19] ;
wire   [8:0] \out_reg[0] ;
wire   [8:0] \out_reg[1] ;
wire   [8:0] \out_reg[2] ;
wire   [8:0] \out_reg[3] ;
wire   [8:0] \out_reg[4] ;
wire   [8:0] \out_reg[5] ;
wire   [8:0] \out_reg[6] ;
wire   [8:0] \out_reg[7] ;
wire   [8:0] \out_reg[8] ;
wire   [8:0] \out_reg[9] ;
wire   [8:0] \out_reg[10] ;
wire   [8:0] \out_reg[11] ;
wire   [8:0] \out_reg[12] ;
wire   [8:0] \out_reg[13] ;
wire   [8:0] \out_reg[14] ;
wire   [8:0] \out_reg[15] ;
wire   [8:0] \out_reg[16] ;
wire   [8:0] \out_reg[17] ;
wire   [8:0] \out_reg[18] ;
wire   [8:0] \out_reg[19] ;
wire   [9:0] \final_sums[0] ;
wire   [9:0] \final_sums[1] ;
wire   [9:0] \final_sums[2] ;
wire   [9:0] \final_sums[3] ;
wire   [9:0] \final_sums[4] ;
wire   [9:0] \final_sums[5] ;
wire   [9:0] \final_sums[6] ;
wire   [9:0] \final_sums[7] ;
wire   [9:0] \final_sums[8] ;
wire   [9:0] \final_sums[9] ;
wire   [9:0] \final_sums[10] ;
wire   [9:0] \final_sums[11] ;
wire   [9:0] \final_sums[12] ;
wire   [9:0] \final_sums[13] ;
wire   [9:0] \final_sums[14] ;
wire   [9:0] \final_sums[15] ;
wire   [9:0] \final_sums[16] ;
wire   [9:0] \final_sums[17] ;
wire   [9:0] \final_sums[18] ;
wire   [9:0] \final_sums[19] ;
wire   [9:0] \level_8_sums[0] ;
wire   [9:0] \level_8_sums[1] ;
wire   [9:0] \level_8_sums[2] ;
wire   [9:0] \level_8_sums[3] ;
wire   [9:0] \level_8_sums[4] ;
wire   [9:0] \level_8_sums[5] ;
wire   [9:0] \level_8_sums[6] ;
wire   [9:0] \level_8_sums[7] ;
wire   [9:0] \level_8_sums[8] ;
wire   [9:0] \level_8_sums[9] ;
wire   [9:0] \level_8_sums[10] ;
wire   [9:0] \level_8_sums[11] ;
wire   [9:0] \level_8_sums[12] ;
wire   [9:0] \level_8_sums[13] ;
wire   [9:0] \level_8_sums[14] ;
wire   [9:0] \level_8_sums[15] ;
wire   [9:0] \level_8_sums[16] ;
wire   [9:0] \level_8_sums[17] ;
wire   [9:0] \level_8_sums[18] ;
wire   [9:0] \level_8_sums[19] ;
wire   [9:0] \level_7_sums[0][0] ;
wire   [9:0] \level_7_sums[0][1] ;
wire   [9:0] \level_7_sums[1][0] ;
wire   [9:0] \level_7_sums[1][1] ;
wire   [9:0] \level_7_sums[2][0] ;
wire   [9:0] \level_7_sums[2][1] ;
wire   [9:0] \level_7_sums[3][0] ;
wire   [9:0] \level_7_sums[3][1] ;
wire   [9:0] \level_7_sums[4][0] ;
wire   [9:0] \level_7_sums[4][1] ;
wire   [9:0] \level_7_sums[5][0] ;
wire   [9:0] \level_7_sums[5][1] ;
wire   [9:0] \level_7_sums[6][0] ;
wire   [9:0] \level_7_sums[6][1] ;
wire   [9:0] \level_7_sums[7][0] ;
wire   [9:0] \level_7_sums[7][1] ;
wire   [9:0] \level_7_sums[8][0] ;
wire   [9:0] \level_7_sums[8][1] ;
wire   [9:0] \level_7_sums[9][0] ;
wire   [9:0] \level_7_sums[9][1] ;
wire   [9:0] \level_7_sums[10][0] ;
wire   [9:0] \level_7_sums[10][1] ;
wire   [9:0] \level_7_sums[11][0] ;
wire   [9:0] \level_7_sums[11][1] ;
wire   [9:0] \level_7_sums[12][0] ;
wire   [9:0] \level_7_sums[12][1] ;
wire   [9:0] \level_7_sums[13][0] ;
wire   [9:0] \level_7_sums[13][1] ;
wire   [9:0] \level_7_sums[14][0] ;
wire   [9:0] \level_7_sums[14][1] ;
wire   [9:0] \level_7_sums[15][0] ;
wire   [9:0] \level_7_sums[15][1] ;
wire   [9:0] \level_7_sums[16][0] ;
wire   [9:0] \level_7_sums[16][1] ;
wire   [9:0] \level_7_sums[17][0] ;
wire   [9:0] \level_7_sums[17][1] ;
wire   [9:0] \level_7_sums[18][0] ;
wire   [9:0] \level_7_sums[18][1] ;
wire   [9:0] \level_7_sums[19][0] ;
wire   [9:0] \level_7_sums[19][1] ;
wire   [9:0] \level_6_sums[0][0] ;
wire   [9:0] \level_6_sums[0][1] ;
wire   [9:0] \level_6_sums[0][2] ;
wire   [9:0] \level_6_sums[0][3] ;
wire   [9:0] \level_6_sums[1][0] ;
wire   [9:0] \level_6_sums[1][1] ;
wire   [9:0] \level_6_sums[1][2] ;
wire   [9:0] \level_6_sums[1][3] ;
wire   [9:0] \level_6_sums[2][0] ;
wire   [9:0] \level_6_sums[2][1] ;
wire   [9:0] \level_6_sums[2][2] ;
wire   [9:0] \level_6_sums[2][3] ;
wire   [9:0] \level_6_sums[3][0] ;
wire   [9:0] \level_6_sums[3][1] ;
wire   [9:0] \level_6_sums[3][2] ;
wire   [9:0] \level_6_sums[3][3] ;
wire   [9:0] \level_6_sums[4][0] ;
wire   [9:0] \level_6_sums[4][1] ;
wire   [9:0] \level_6_sums[4][2] ;
wire   [9:0] \level_6_sums[4][3] ;
wire   [9:0] \level_6_sums[5][0] ;
wire   [9:0] \level_6_sums[5][1] ;
wire   [9:0] \level_6_sums[5][2] ;
wire   [9:0] \level_6_sums[5][3] ;
wire   [9:0] \level_6_sums[6][0] ;
wire   [9:0] \level_6_sums[6][1] ;
wire   [9:0] \level_6_sums[6][2] ;
wire   [9:0] \level_6_sums[6][3] ;
wire   [9:0] \level_6_sums[7][0] ;
wire   [9:0] \level_6_sums[7][1] ;
wire   [9:0] \level_6_sums[7][2] ;
wire   [9:0] \level_6_sums[7][3] ;
wire   [9:0] \level_6_sums[8][0] ;
wire   [9:0] \level_6_sums[8][1] ;
wire   [9:0] \level_6_sums[8][2] ;
wire   [9:0] \level_6_sums[8][3] ;
wire   [9:0] \level_6_sums[9][0] ;
wire   [9:0] \level_6_sums[9][1] ;
wire   [9:0] \level_6_sums[9][2] ;
wire   [9:0] \level_6_sums[9][3] ;
wire   [9:0] \level_6_sums[10][0] ;
wire   [9:0] \level_6_sums[10][1] ;
wire   [9:0] \level_6_sums[10][2] ;
wire   [9:0] \level_6_sums[10][3] ;
wire   [9:0] \level_6_sums[11][0] ;
wire   [9:0] \level_6_sums[11][1] ;
wire   [9:0] \level_6_sums[11][2] ;
wire   [9:0] \level_6_sums[11][3] ;
wire   [9:0] \level_6_sums[12][0] ;
wire   [9:0] \level_6_sums[12][1] ;
wire   [9:0] \level_6_sums[12][2] ;
wire   [9:0] \level_6_sums[12][3] ;
wire   [9:0] \level_6_sums[13][0] ;
wire   [9:0] \level_6_sums[13][1] ;
wire   [9:0] \level_6_sums[13][2] ;
wire   [9:0] \level_6_sums[13][3] ;
wire   [9:0] \level_6_sums[14][0] ;
wire   [9:0] \level_6_sums[14][1] ;
wire   [9:0] \level_6_sums[14][2] ;
wire   [9:0] \level_6_sums[14][3] ;
wire   [9:0] \level_6_sums[15][0] ;
wire   [9:0] \level_6_sums[15][1] ;
wire   [9:0] \level_6_sums[15][2] ;
wire   [9:0] \level_6_sums[15][3] ;
wire   [9:0] \level_6_sums[16][0] ;
wire   [9:0] \level_6_sums[16][1] ;
wire   [9:0] \level_6_sums[16][2] ;
wire   [9:0] \level_6_sums[16][3] ;
wire   [9:0] \level_6_sums[17][0] ;
wire   [9:0] \level_6_sums[17][1] ;
wire   [9:0] \level_6_sums[17][2] ;
wire   [9:0] \level_6_sums[17][3] ;
wire   [9:0] \level_6_sums[18][0] ;
wire   [9:0] \level_6_sums[18][1] ;
wire   [9:0] \level_6_sums[18][2] ;
wire   [9:0] \level_6_sums[18][3] ;
wire   [9:0] \level_6_sums[19][0] ;
wire   [9:0] \level_6_sums[19][1] ;
wire   [9:0] \level_6_sums[19][2] ;
wire   [9:0] \level_6_sums[19][3] ;
wire   [9:0] \level_5_sums[0][0] ;
wire   [9:0] \level_5_sums[0][1] ;
wire   [9:0] \level_5_sums[0][2] ;
wire   [9:0] \level_5_sums[0][3] ;
wire   [9:0] \level_5_sums[0][4] ;
wire   [9:0] \level_5_sums[0][5] ;
wire   [9:0] \level_5_sums[0][6] ;
wire   [9:0] \level_5_sums[0][7] ;
wire   [9:0] \level_5_sums[1][0] ;
wire   [9:0] \level_5_sums[1][1] ;
wire   [9:0] \level_5_sums[1][2] ;
wire   [9:0] \level_5_sums[1][3] ;
wire   [9:0] \level_5_sums[1][4] ;
wire   [9:0] \level_5_sums[1][5] ;
wire   [9:0] \level_5_sums[1][6] ;
wire   [9:0] \level_5_sums[1][7] ;
wire   [9:0] \level_5_sums[2][0] ;
wire   [9:0] \level_5_sums[2][1] ;
wire   [9:0] \level_5_sums[2][2] ;
wire   [9:0] \level_5_sums[2][3] ;
wire   [9:0] \level_5_sums[2][4] ;
wire   [9:0] \level_5_sums[2][5] ;
wire   [9:0] \level_5_sums[2][6] ;
wire   [9:0] \level_5_sums[2][7] ;
wire   [9:0] \level_5_sums[3][0] ;
wire   [9:0] \level_5_sums[3][1] ;
wire   [9:0] \level_5_sums[3][2] ;
wire   [9:0] \level_5_sums[3][3] ;
wire   [9:0] \level_5_sums[3][4] ;
wire   [9:0] \level_5_sums[3][5] ;
wire   [9:0] \level_5_sums[3][6] ;
wire   [9:0] \level_5_sums[3][7] ;
wire   [9:0] \level_5_sums[4][0] ;
wire   [9:0] \level_5_sums[4][1] ;
wire   [9:0] \level_5_sums[4][2] ;
wire   [9:0] \level_5_sums[4][3] ;
wire   [9:0] \level_5_sums[4][4] ;
wire   [9:0] \level_5_sums[4][5] ;
wire   [9:0] \level_5_sums[4][6] ;
wire   [9:0] \level_5_sums[4][7] ;
wire   [9:0] \level_5_sums[5][0] ;
wire   [9:0] \level_5_sums[5][1] ;
wire   [9:0] \level_5_sums[5][2] ;
wire   [9:0] \level_5_sums[5][3] ;
wire   [9:0] \level_5_sums[5][4] ;
wire   [9:0] \level_5_sums[5][5] ;
wire   [9:0] \level_5_sums[5][6] ;
wire   [9:0] \level_5_sums[5][7] ;
wire   [9:0] \level_5_sums[6][0] ;
wire   [9:0] \level_5_sums[6][1] ;
wire   [9:0] \level_5_sums[6][2] ;
wire   [9:0] \level_5_sums[6][3] ;
wire   [9:0] \level_5_sums[6][4] ;
wire   [9:0] \level_5_sums[6][5] ;
wire   [9:0] \level_5_sums[6][6] ;
wire   [9:0] \level_5_sums[6][7] ;
wire   [9:0] \level_5_sums[7][0] ;
wire   [9:0] \level_5_sums[7][1] ;
wire   [9:0] \level_5_sums[7][2] ;
wire   [9:0] \level_5_sums[7][3] ;
wire   [9:0] \level_5_sums[7][4] ;
wire   [9:0] \level_5_sums[7][5] ;
wire   [9:0] \level_5_sums[7][6] ;
wire   [9:0] \level_5_sums[7][7] ;
wire   [9:0] \level_5_sums[8][0] ;
wire   [9:0] \level_5_sums[8][1] ;
wire   [9:0] \level_5_sums[8][2] ;
wire   [9:0] \level_5_sums[8][3] ;
wire   [9:0] \level_5_sums[8][4] ;
wire   [9:0] \level_5_sums[8][5] ;
wire   [9:0] \level_5_sums[8][6] ;
wire   [9:0] \level_5_sums[8][7] ;
wire   [9:0] \level_5_sums[9][0] ;
wire   [9:0] \level_5_sums[9][1] ;
wire   [9:0] \level_5_sums[9][2] ;
wire   [9:0] \level_5_sums[9][3] ;
wire   [9:0] \level_5_sums[9][4] ;
wire   [9:0] \level_5_sums[9][5] ;
wire   [9:0] \level_5_sums[9][6] ;
wire   [9:0] \level_5_sums[9][7] ;
wire   [9:0] \level_5_sums[10][0] ;
wire   [9:0] \level_5_sums[10][1] ;
wire   [9:0] \level_5_sums[10][2] ;
wire   [9:0] \level_5_sums[10][3] ;
wire   [9:0] \level_5_sums[10][4] ;
wire   [9:0] \level_5_sums[10][5] ;
wire   [9:0] \level_5_sums[10][6] ;
wire   [9:0] \level_5_sums[10][7] ;
wire   [9:0] \level_5_sums[11][0] ;
wire   [9:0] \level_5_sums[11][1] ;
wire   [9:0] \level_5_sums[11][2] ;
wire   [9:0] \level_5_sums[11][3] ;
wire   [9:0] \level_5_sums[11][4] ;
wire   [9:0] \level_5_sums[11][5] ;
wire   [9:0] \level_5_sums[11][6] ;
wire   [9:0] \level_5_sums[11][7] ;
wire   [9:0] \level_5_sums[12][0] ;
wire   [9:0] \level_5_sums[12][1] ;
wire   [9:0] \level_5_sums[12][2] ;
wire   [9:0] \level_5_sums[12][3] ;
wire   [9:0] \level_5_sums[12][4] ;
wire   [9:0] \level_5_sums[12][5] ;
wire   [9:0] \level_5_sums[12][6] ;
wire   [9:0] \level_5_sums[12][7] ;
wire   [9:0] \level_5_sums[13][0] ;
wire   [9:0] \level_5_sums[13][1] ;
wire   [9:0] \level_5_sums[13][2] ;
wire   [9:0] \level_5_sums[13][3] ;
wire   [9:0] \level_5_sums[13][4] ;
wire   [9:0] \level_5_sums[13][5] ;
wire   [9:0] \level_5_sums[13][6] ;
wire   [9:0] \level_5_sums[13][7] ;
wire   [9:0] \level_5_sums[14][0] ;
wire   [9:0] \level_5_sums[14][1] ;
wire   [9:0] \level_5_sums[14][2] ;
wire   [9:0] \level_5_sums[14][3] ;
wire   [9:0] \level_5_sums[14][4] ;
wire   [9:0] \level_5_sums[14][5] ;
wire   [9:0] \level_5_sums[14][6] ;
wire   [9:0] \level_5_sums[14][7] ;
wire   [9:0] \level_5_sums[15][0] ;
wire   [9:0] \level_5_sums[15][1] ;
wire   [9:0] \level_5_sums[15][2] ;
wire   [9:0] \level_5_sums[15][3] ;
wire   [9:0] \level_5_sums[15][4] ;
wire   [9:0] \level_5_sums[15][5] ;
wire   [9:0] \level_5_sums[15][6] ;
wire   [9:0] \level_5_sums[15][7] ;
wire   [9:0] \level_5_sums[16][0] ;
wire   [9:0] \level_5_sums[16][1] ;
wire   [9:0] \level_5_sums[16][2] ;
wire   [9:0] \level_5_sums[16][3] ;
wire   [9:0] \level_5_sums[16][4] ;
wire   [9:0] \level_5_sums[16][5] ;
wire   [9:0] \level_5_sums[16][6] ;
wire   [9:0] \level_5_sums[16][7] ;
wire   [9:0] \level_5_sums[17][0] ;
wire   [9:0] \level_5_sums[17][1] ;
wire   [9:0] \level_5_sums[17][2] ;
wire   [9:0] \level_5_sums[17][3] ;
wire   [9:0] \level_5_sums[17][4] ;
wire   [9:0] \level_5_sums[17][5] ;
wire   [9:0] \level_5_sums[17][6] ;
wire   [9:0] \level_5_sums[17][7] ;
wire   [9:0] \level_5_sums[18][0] ;
wire   [9:0] \level_5_sums[18][1] ;
wire   [9:0] \level_5_sums[18][2] ;
wire   [9:0] \level_5_sums[18][3] ;
wire   [9:0] \level_5_sums[18][4] ;
wire   [9:0] \level_5_sums[18][5] ;
wire   [9:0] \level_5_sums[18][6] ;
wire   [9:0] \level_5_sums[18][7] ;
wire   [9:0] \level_5_sums[19][0] ;
wire   [9:0] \level_5_sums[19][1] ;
wire   [9:0] \level_5_sums[19][2] ;
wire   [9:0] \level_5_sums[19][3] ;
wire   [9:0] \level_5_sums[19][4] ;
wire   [9:0] \level_5_sums[19][5] ;
wire   [9:0] \level_5_sums[19][6] ;
wire   [9:0] \level_5_sums[19][7] ;
wire   [8:0] \level_4_sums[0][0] ;
wire   [8:0] \level_4_sums[0][1] ;
wire   [8:0] \level_4_sums[0][2] ;
wire   [8:0] \level_4_sums[0][3] ;
wire   [8:0] \level_4_sums[0][4] ;
wire   [8:0] \level_4_sums[0][5] ;
wire   [8:0] \level_4_sums[0][6] ;
wire   [8:0] \level_4_sums[0][7] ;
wire   [8:0] \level_4_sums[0][8] ;
wire   [8:0] \level_4_sums[0][9] ;
wire   [8:0] \level_4_sums[0][10] ;
wire   [8:0] \level_4_sums[0][11] ;
wire   [8:0] \level_4_sums[0][12] ;
wire   [8:0] \level_4_sums[0][13] ;
wire   [8:0] \level_4_sums[0][14] ;
wire   [8:0] \level_4_sums[0][15] ;
wire   [8:0] \level_4_sums[1][0] ;
wire   [8:0] \level_4_sums[1][1] ;
wire   [8:0] \level_4_sums[1][2] ;
wire   [8:0] \level_4_sums[1][3] ;
wire   [8:0] \level_4_sums[1][4] ;
wire   [8:0] \level_4_sums[1][5] ;
wire   [8:0] \level_4_sums[1][6] ;
wire   [8:0] \level_4_sums[1][7] ;
wire   [8:0] \level_4_sums[1][8] ;
wire   [8:0] \level_4_sums[1][9] ;
wire   [8:0] \level_4_sums[1][10] ;
wire   [8:0] \level_4_sums[1][11] ;
wire   [8:0] \level_4_sums[1][12] ;
wire   [8:0] \level_4_sums[1][13] ;
wire   [8:0] \level_4_sums[1][14] ;
wire   [8:0] \level_4_sums[1][15] ;
wire   [8:0] \level_4_sums[2][0] ;
wire   [8:0] \level_4_sums[2][1] ;
wire   [8:0] \level_4_sums[2][2] ;
wire   [8:0] \level_4_sums[2][3] ;
wire   [8:0] \level_4_sums[2][4] ;
wire   [8:0] \level_4_sums[2][5] ;
wire   [8:0] \level_4_sums[2][6] ;
wire   [8:0] \level_4_sums[2][7] ;
wire   [8:0] \level_4_sums[2][8] ;
wire   [8:0] \level_4_sums[2][9] ;
wire   [8:0] \level_4_sums[2][10] ;
wire   [8:0] \level_4_sums[2][11] ;
wire   [8:0] \level_4_sums[2][12] ;
wire   [8:0] \level_4_sums[2][13] ;
wire   [8:0] \level_4_sums[2][14] ;
wire   [8:0] \level_4_sums[2][15] ;
wire   [8:0] \level_4_sums[3][0] ;
wire   [8:0] \level_4_sums[3][1] ;
wire   [8:0] \level_4_sums[3][2] ;
wire   [8:0] \level_4_sums[3][3] ;
wire   [8:0] \level_4_sums[3][4] ;
wire   [8:0] \level_4_sums[3][5] ;
wire   [8:0] \level_4_sums[3][6] ;
wire   [8:0] \level_4_sums[3][7] ;
wire   [8:0] \level_4_sums[3][8] ;
wire   [8:0] \level_4_sums[3][9] ;
wire   [8:0] \level_4_sums[3][10] ;
wire   [8:0] \level_4_sums[3][11] ;
wire   [8:0] \level_4_sums[3][12] ;
wire   [8:0] \level_4_sums[3][13] ;
wire   [8:0] \level_4_sums[3][14] ;
wire   [8:0] \level_4_sums[3][15] ;
wire   [8:0] \level_4_sums[4][0] ;
wire   [8:0] \level_4_sums[4][1] ;
wire   [8:0] \level_4_sums[4][2] ;
wire   [8:0] \level_4_sums[4][3] ;
wire   [8:0] \level_4_sums[4][4] ;
wire   [8:0] \level_4_sums[4][5] ;
wire   [8:0] \level_4_sums[4][6] ;
wire   [8:0] \level_4_sums[4][7] ;
wire   [8:0] \level_4_sums[4][8] ;
wire   [8:0] \level_4_sums[4][9] ;
wire   [8:0] \level_4_sums[4][10] ;
wire   [8:0] \level_4_sums[4][11] ;
wire   [8:0] \level_4_sums[4][12] ;
wire   [8:0] \level_4_sums[4][13] ;
wire   [8:0] \level_4_sums[4][14] ;
wire   [8:0] \level_4_sums[4][15] ;
wire   [8:0] \level_4_sums[5][0] ;
wire   [8:0] \level_4_sums[5][1] ;
wire   [8:0] \level_4_sums[5][2] ;
wire   [8:0] \level_4_sums[5][3] ;
wire   [8:0] \level_4_sums[5][4] ;
wire   [8:0] \level_4_sums[5][5] ;
wire   [8:0] \level_4_sums[5][6] ;
wire   [8:0] \level_4_sums[5][7] ;
wire   [8:0] \level_4_sums[5][8] ;
wire   [8:0] \level_4_sums[5][9] ;
wire   [8:0] \level_4_sums[5][10] ;
wire   [8:0] \level_4_sums[5][11] ;
wire   [8:0] \level_4_sums[5][12] ;
wire   [8:0] \level_4_sums[5][13] ;
wire   [8:0] \level_4_sums[5][14] ;
wire   [8:0] \level_4_sums[5][15] ;
wire   [8:0] \level_4_sums[6][0] ;
wire   [8:0] \level_4_sums[6][1] ;
wire   [8:0] \level_4_sums[6][2] ;
wire   [8:0] \level_4_sums[6][3] ;
wire   [8:0] \level_4_sums[6][4] ;
wire   [8:0] \level_4_sums[6][5] ;
wire   [8:0] \level_4_sums[6][6] ;
wire   [8:0] \level_4_sums[6][7] ;
wire   [8:0] \level_4_sums[6][8] ;
wire   [8:0] \level_4_sums[6][9] ;
wire   [8:0] \level_4_sums[6][10] ;
wire   [8:0] \level_4_sums[6][11] ;
wire   [8:0] \level_4_sums[6][12] ;
wire   [8:0] \level_4_sums[6][13] ;
wire   [8:0] \level_4_sums[6][14] ;
wire   [8:0] \level_4_sums[6][15] ;
wire   [8:0] \level_4_sums[7][0] ;
wire   [8:0] \level_4_sums[7][1] ;
wire   [8:0] \level_4_sums[7][2] ;
wire   [8:0] \level_4_sums[7][3] ;
wire   [8:0] \level_4_sums[7][4] ;
wire   [8:0] \level_4_sums[7][5] ;
wire   [8:0] \level_4_sums[7][6] ;
wire   [8:0] \level_4_sums[7][7] ;
wire   [8:0] \level_4_sums[7][8] ;
wire   [8:0] \level_4_sums[7][9] ;
wire   [8:0] \level_4_sums[7][10] ;
wire   [8:0] \level_4_sums[7][11] ;
wire   [8:0] \level_4_sums[7][12] ;
wire   [8:0] \level_4_sums[7][13] ;
wire   [8:0] \level_4_sums[7][14] ;
wire   [8:0] \level_4_sums[7][15] ;
wire   [8:0] \level_4_sums[8][0] ;
wire   [8:0] \level_4_sums[8][1] ;
wire   [8:0] \level_4_sums[8][2] ;
wire   [8:0] \level_4_sums[8][3] ;
wire   [8:0] \level_4_sums[8][4] ;
wire   [8:0] \level_4_sums[8][5] ;
wire   [8:0] \level_4_sums[8][6] ;
wire   [8:0] \level_4_sums[8][7] ;
wire   [8:0] \level_4_sums[8][8] ;
wire   [8:0] \level_4_sums[8][9] ;
wire   [8:0] \level_4_sums[8][10] ;
wire   [8:0] \level_4_sums[8][11] ;
wire   [8:0] \level_4_sums[8][12] ;
wire   [8:0] \level_4_sums[8][13] ;
wire   [8:0] \level_4_sums[8][14] ;
wire   [8:0] \level_4_sums[8][15] ;
wire   [8:0] \level_4_sums[9][0] ;
wire   [8:0] \level_4_sums[9][1] ;
wire   [8:0] \level_4_sums[9][2] ;
wire   [8:0] \level_4_sums[9][3] ;
wire   [8:0] \level_4_sums[9][4] ;
wire   [8:0] \level_4_sums[9][5] ;
wire   [8:0] \level_4_sums[9][6] ;
wire   [8:0] \level_4_sums[9][7] ;
wire   [8:0] \level_4_sums[9][8] ;
wire   [8:0] \level_4_sums[9][9] ;
wire   [8:0] \level_4_sums[9][10] ;
wire   [8:0] \level_4_sums[9][11] ;
wire   [8:0] \level_4_sums[9][12] ;
wire   [8:0] \level_4_sums[9][13] ;
wire   [8:0] \level_4_sums[9][14] ;
wire   [8:0] \level_4_sums[9][15] ;
wire   [8:0] \level_4_sums[10][0] ;
wire   [8:0] \level_4_sums[10][1] ;
wire   [8:0] \level_4_sums[10][2] ;
wire   [8:0] \level_4_sums[10][3] ;
wire   [8:0] \level_4_sums[10][4] ;
wire   [8:0] \level_4_sums[10][5] ;
wire   [8:0] \level_4_sums[10][6] ;
wire   [8:0] \level_4_sums[10][7] ;
wire   [8:0] \level_4_sums[10][8] ;
wire   [8:0] \level_4_sums[10][9] ;
wire   [8:0] \level_4_sums[10][10] ;
wire   [8:0] \level_4_sums[10][11] ;
wire   [8:0] \level_4_sums[10][12] ;
wire   [8:0] \level_4_sums[10][13] ;
wire   [8:0] \level_4_sums[10][14] ;
wire   [8:0] \level_4_sums[10][15] ;
wire   [8:0] \level_4_sums[11][0] ;
wire   [8:0] \level_4_sums[11][1] ;
wire   [8:0] \level_4_sums[11][2] ;
wire   [8:0] \level_4_sums[11][3] ;
wire   [8:0] \level_4_sums[11][4] ;
wire   [8:0] \level_4_sums[11][5] ;
wire   [8:0] \level_4_sums[11][6] ;
wire   [8:0] \level_4_sums[11][7] ;
wire   [8:0] \level_4_sums[11][8] ;
wire   [8:0] \level_4_sums[11][9] ;
wire   [8:0] \level_4_sums[11][10] ;
wire   [8:0] \level_4_sums[11][11] ;
wire   [8:0] \level_4_sums[11][12] ;
wire   [8:0] \level_4_sums[11][13] ;
wire   [8:0] \level_4_sums[11][14] ;
wire   [8:0] \level_4_sums[11][15] ;
wire   [8:0] \level_4_sums[12][0] ;
wire   [8:0] \level_4_sums[12][1] ;
wire   [8:0] \level_4_sums[12][2] ;
wire   [8:0] \level_4_sums[12][3] ;
wire   [8:0] \level_4_sums[12][4] ;
wire   [8:0] \level_4_sums[12][5] ;
wire   [8:0] \level_4_sums[12][6] ;
wire   [8:0] \level_4_sums[12][7] ;
wire   [8:0] \level_4_sums[12][8] ;
wire   [8:0] \level_4_sums[12][9] ;
wire   [8:0] \level_4_sums[12][10] ;
wire   [8:0] \level_4_sums[12][11] ;
wire   [8:0] \level_4_sums[12][12] ;
wire   [8:0] \level_4_sums[12][13] ;
wire   [8:0] \level_4_sums[12][14] ;
wire   [8:0] \level_4_sums[12][15] ;
wire   [8:0] \level_4_sums[13][0] ;
wire   [8:0] \level_4_sums[13][1] ;
wire   [8:0] \level_4_sums[13][2] ;
wire   [8:0] \level_4_sums[13][3] ;
wire   [8:0] \level_4_sums[13][4] ;
wire   [8:0] \level_4_sums[13][5] ;
wire   [8:0] \level_4_sums[13][6] ;
wire   [8:0] \level_4_sums[13][7] ;
wire   [8:0] \level_4_sums[13][8] ;
wire   [8:0] \level_4_sums[13][9] ;
wire   [8:0] \level_4_sums[13][10] ;
wire   [8:0] \level_4_sums[13][11] ;
wire   [8:0] \level_4_sums[13][12] ;
wire   [8:0] \level_4_sums[13][13] ;
wire   [8:0] \level_4_sums[13][14] ;
wire   [8:0] \level_4_sums[13][15] ;
wire   [8:0] \level_4_sums[14][0] ;
wire   [8:0] \level_4_sums[14][1] ;
wire   [8:0] \level_4_sums[14][2] ;
wire   [8:0] \level_4_sums[14][3] ;
wire   [8:0] \level_4_sums[14][4] ;
wire   [8:0] \level_4_sums[14][5] ;
wire   [8:0] \level_4_sums[14][6] ;
wire   [8:0] \level_4_sums[14][7] ;
wire   [8:0] \level_4_sums[14][8] ;
wire   [8:0] \level_4_sums[14][9] ;
wire   [8:0] \level_4_sums[14][10] ;
wire   [8:0] \level_4_sums[14][11] ;
wire   [8:0] \level_4_sums[14][12] ;
wire   [8:0] \level_4_sums[14][13] ;
wire   [8:0] \level_4_sums[14][14] ;
wire   [8:0] \level_4_sums[14][15] ;
wire   [8:0] \level_4_sums[15][0] ;
wire   [8:0] \level_4_sums[15][1] ;
wire   [8:0] \level_4_sums[15][2] ;
wire   [8:0] \level_4_sums[15][3] ;
wire   [8:0] \level_4_sums[15][4] ;
wire   [8:0] \level_4_sums[15][5] ;
wire   [8:0] \level_4_sums[15][6] ;
wire   [8:0] \level_4_sums[15][7] ;
wire   [8:0] \level_4_sums[15][8] ;
wire   [8:0] \level_4_sums[15][9] ;
wire   [8:0] \level_4_sums[15][10] ;
wire   [8:0] \level_4_sums[15][11] ;
wire   [8:0] \level_4_sums[15][12] ;
wire   [8:0] \level_4_sums[15][13] ;
wire   [8:0] \level_4_sums[15][14] ;
wire   [8:0] \level_4_sums[15][15] ;
wire   [8:0] \level_4_sums[16][0] ;
wire   [8:0] \level_4_sums[16][1] ;
wire   [8:0] \level_4_sums[16][2] ;
wire   [8:0] \level_4_sums[16][3] ;
wire   [8:0] \level_4_sums[16][4] ;
wire   [8:0] \level_4_sums[16][5] ;
wire   [8:0] \level_4_sums[16][6] ;
wire   [8:0] \level_4_sums[16][7] ;
wire   [8:0] \level_4_sums[16][8] ;
wire   [8:0] \level_4_sums[16][9] ;
wire   [8:0] \level_4_sums[16][10] ;
wire   [8:0] \level_4_sums[16][11] ;
wire   [8:0] \level_4_sums[16][12] ;
wire   [8:0] \level_4_sums[16][13] ;
wire   [8:0] \level_4_sums[16][14] ;
wire   [8:0] \level_4_sums[16][15] ;
wire   [8:0] \level_4_sums[17][0] ;
wire   [8:0] \level_4_sums[17][1] ;
wire   [8:0] \level_4_sums[17][2] ;
wire   [8:0] \level_4_sums[17][3] ;
wire   [8:0] \level_4_sums[17][4] ;
wire   [8:0] \level_4_sums[17][5] ;
wire   [8:0] \level_4_sums[17][6] ;
wire   [8:0] \level_4_sums[17][7] ;
wire   [8:0] \level_4_sums[17][8] ;
wire   [8:0] \level_4_sums[17][9] ;
wire   [8:0] \level_4_sums[17][10] ;
wire   [8:0] \level_4_sums[17][11] ;
wire   [8:0] \level_4_sums[17][12] ;
wire   [8:0] \level_4_sums[17][13] ;
wire   [8:0] \level_4_sums[17][14] ;
wire   [8:0] \level_4_sums[17][15] ;
wire   [8:0] \level_4_sums[18][0] ;
wire   [8:0] \level_4_sums[18][1] ;
wire   [8:0] \level_4_sums[18][2] ;
wire   [8:0] \level_4_sums[18][3] ;
wire   [8:0] \level_4_sums[18][4] ;
wire   [8:0] \level_4_sums[18][5] ;
wire   [8:0] \level_4_sums[18][6] ;
wire   [8:0] \level_4_sums[18][7] ;
wire   [8:0] \level_4_sums[18][8] ;
wire   [8:0] \level_4_sums[18][9] ;
wire   [8:0] \level_4_sums[18][10] ;
wire   [8:0] \level_4_sums[18][11] ;
wire   [8:0] \level_4_sums[18][12] ;
wire   [8:0] \level_4_sums[18][13] ;
wire   [8:0] \level_4_sums[18][14] ;
wire   [8:0] \level_4_sums[18][15] ;
wire   [8:0] \level_4_sums[19][0] ;
wire   [8:0] \level_4_sums[19][1] ;
wire   [8:0] \level_4_sums[19][2] ;
wire   [8:0] \level_4_sums[19][3] ;
wire   [8:0] \level_4_sums[19][4] ;
wire   [8:0] \level_4_sums[19][5] ;
wire   [8:0] \level_4_sums[19][6] ;
wire   [8:0] \level_4_sums[19][7] ;
wire   [8:0] \level_4_sums[19][8] ;
wire   [8:0] \level_4_sums[19][9] ;
wire   [8:0] \level_4_sums[19][10] ;
wire   [8:0] \level_4_sums[19][11] ;
wire   [8:0] \level_4_sums[19][12] ;
wire   [8:0] \level_4_sums[19][13] ;
wire   [8:0] \level_4_sums[19][14] ;
wire   [8:0] \level_4_sums[19][15] ;
wire   [7:0] \level_3_sums[0][0] ;
wire   [7:0] \level_3_sums[0][1] ;
wire   [7:0] \level_3_sums[0][2] ;
wire   [7:0] \level_3_sums[0][3] ;
wire   [7:0] \level_3_sums[0][4] ;
wire   [7:0] \level_3_sums[0][5] ;
wire   [7:0] \level_3_sums[0][6] ;
wire   [7:0] \level_3_sums[0][7] ;
wire   [7:0] \level_3_sums[0][8] ;
wire   [7:0] \level_3_sums[0][9] ;
wire   [7:0] \level_3_sums[0][10] ;
wire   [7:0] \level_3_sums[0][11] ;
wire   [7:0] \level_3_sums[0][12] ;
wire   [7:0] \level_3_sums[0][13] ;
wire   [7:0] \level_3_sums[0][14] ;
wire   [7:0] \level_3_sums[0][15] ;
wire   [7:0] \level_3_sums[0][16] ;
wire   [7:0] \level_3_sums[0][17] ;
wire   [7:0] \level_3_sums[0][18] ;
wire   [7:0] \level_3_sums[0][19] ;
wire   [7:0] \level_3_sums[0][20] ;
wire   [7:0] \level_3_sums[0][21] ;
wire   [7:0] \level_3_sums[0][22] ;
wire   [7:0] \level_3_sums[0][23] ;
wire   [7:0] \level_3_sums[0][24] ;
wire   [7:0] \level_3_sums[0][25] ;
wire   [7:0] \level_3_sums[0][26] ;
wire   [7:0] \level_3_sums[0][27] ;
wire   [7:0] \level_3_sums[0][28] ;
wire   [7:0] \level_3_sums[0][29] ;
wire   [7:0] \level_3_sums[0][30] ;
wire   [7:0] \level_3_sums[0][31] ;
wire   [7:0] \level_3_sums[1][0] ;
wire   [7:0] \level_3_sums[1][1] ;
wire   [7:0] \level_3_sums[1][2] ;
wire   [7:0] \level_3_sums[1][3] ;
wire   [7:0] \level_3_sums[1][4] ;
wire   [7:0] \level_3_sums[1][5] ;
wire   [7:0] \level_3_sums[1][6] ;
wire   [7:0] \level_3_sums[1][7] ;
wire   [7:0] \level_3_sums[1][8] ;
wire   [7:0] \level_3_sums[1][9] ;
wire   [7:0] \level_3_sums[1][10] ;
wire   [7:0] \level_3_sums[1][11] ;
wire   [7:0] \level_3_sums[1][12] ;
wire   [7:0] \level_3_sums[1][13] ;
wire   [7:0] \level_3_sums[1][14] ;
wire   [7:0] \level_3_sums[1][15] ;
wire   [7:0] \level_3_sums[1][16] ;
wire   [7:0] \level_3_sums[1][17] ;
wire   [7:0] \level_3_sums[1][18] ;
wire   [7:0] \level_3_sums[1][19] ;
wire   [7:0] \level_3_sums[1][20] ;
wire   [7:0] \level_3_sums[1][21] ;
wire   [7:0] \level_3_sums[1][22] ;
wire   [7:0] \level_3_sums[1][23] ;
wire   [7:0] \level_3_sums[1][24] ;
wire   [7:0] \level_3_sums[1][25] ;
wire   [7:0] \level_3_sums[1][26] ;
wire   [7:0] \level_3_sums[1][27] ;
wire   [7:0] \level_3_sums[1][28] ;
wire   [7:0] \level_3_sums[1][29] ;
wire   [7:0] \level_3_sums[1][30] ;
wire   [7:0] \level_3_sums[1][31] ;
wire   [7:0] \level_3_sums[2][0] ;
wire   [7:0] \level_3_sums[2][1] ;
wire   [7:0] \level_3_sums[2][2] ;
wire   [7:0] \level_3_sums[2][3] ;
wire   [7:0] \level_3_sums[2][4] ;
wire   [7:0] \level_3_sums[2][5] ;
wire   [7:0] \level_3_sums[2][6] ;
wire   [7:0] \level_3_sums[2][7] ;
wire   [7:0] \level_3_sums[2][8] ;
wire   [7:0] \level_3_sums[2][9] ;
wire   [7:0] \level_3_sums[2][10] ;
wire   [7:0] \level_3_sums[2][11] ;
wire   [7:0] \level_3_sums[2][12] ;
wire   [7:0] \level_3_sums[2][13] ;
wire   [7:0] \level_3_sums[2][14] ;
wire   [7:0] \level_3_sums[2][15] ;
wire   [7:0] \level_3_sums[2][16] ;
wire   [7:0] \level_3_sums[2][17] ;
wire   [7:0] \level_3_sums[2][18] ;
wire   [7:0] \level_3_sums[2][19] ;
wire   [7:0] \level_3_sums[2][20] ;
wire   [7:0] \level_3_sums[2][21] ;
wire   [7:0] \level_3_sums[2][22] ;
wire   [7:0] \level_3_sums[2][23] ;
wire   [7:0] \level_3_sums[2][24] ;
wire   [7:0] \level_3_sums[2][25] ;
wire   [7:0] \level_3_sums[2][26] ;
wire   [7:0] \level_3_sums[2][27] ;
wire   [7:0] \level_3_sums[2][28] ;
wire   [7:0] \level_3_sums[2][29] ;
wire   [7:0] \level_3_sums[2][30] ;
wire   [7:0] \level_3_sums[2][31] ;
wire   [7:0] \level_3_sums[3][0] ;
wire   [7:0] \level_3_sums[3][1] ;
wire   [7:0] \level_3_sums[3][2] ;
wire   [7:0] \level_3_sums[3][3] ;
wire   [7:0] \level_3_sums[3][4] ;
wire   [7:0] \level_3_sums[3][5] ;
wire   [7:0] \level_3_sums[3][6] ;
wire   [7:0] \level_3_sums[3][7] ;
wire   [7:0] \level_3_sums[3][8] ;
wire   [7:0] \level_3_sums[3][9] ;
wire   [7:0] \level_3_sums[3][10] ;
wire   [7:0] \level_3_sums[3][11] ;
wire   [7:0] \level_3_sums[3][12] ;
wire   [7:0] \level_3_sums[3][13] ;
wire   [7:0] \level_3_sums[3][14] ;
wire   [7:0] \level_3_sums[3][15] ;
wire   [7:0] \level_3_sums[3][16] ;
wire   [7:0] \level_3_sums[3][17] ;
wire   [7:0] \level_3_sums[3][18] ;
wire   [7:0] \level_3_sums[3][19] ;
wire   [7:0] \level_3_sums[3][20] ;
wire   [7:0] \level_3_sums[3][21] ;
wire   [7:0] \level_3_sums[3][22] ;
wire   [7:0] \level_3_sums[3][23] ;
wire   [7:0] \level_3_sums[3][24] ;
wire   [7:0] \level_3_sums[3][25] ;
wire   [7:0] \level_3_sums[3][26] ;
wire   [7:0] \level_3_sums[3][27] ;
wire   [7:0] \level_3_sums[3][28] ;
wire   [7:0] \level_3_sums[3][29] ;
wire   [7:0] \level_3_sums[3][30] ;
wire   [7:0] \level_3_sums[3][31] ;
wire   [7:0] \level_3_sums[4][0] ;
wire   [7:0] \level_3_sums[4][1] ;
wire   [7:0] \level_3_sums[4][2] ;
wire   [7:0] \level_3_sums[4][3] ;
wire   [7:0] \level_3_sums[4][4] ;
wire   [7:0] \level_3_sums[4][5] ;
wire   [7:0] \level_3_sums[4][6] ;
wire   [7:0] \level_3_sums[4][7] ;
wire   [7:0] \level_3_sums[4][8] ;
wire   [7:0] \level_3_sums[4][9] ;
wire   [7:0] \level_3_sums[4][10] ;
wire   [7:0] \level_3_sums[4][11] ;
wire   [7:0] \level_3_sums[4][12] ;
wire   [7:0] \level_3_sums[4][13] ;
wire   [7:0] \level_3_sums[4][14] ;
wire   [7:0] \level_3_sums[4][15] ;
wire   [7:0] \level_3_sums[4][16] ;
wire   [7:0] \level_3_sums[4][17] ;
wire   [7:0] \level_3_sums[4][18] ;
wire   [7:0] \level_3_sums[4][19] ;
wire   [7:0] \level_3_sums[4][20] ;
wire   [7:0] \level_3_sums[4][21] ;
wire   [7:0] \level_3_sums[4][22] ;
wire   [7:0] \level_3_sums[4][23] ;
wire   [7:0] \level_3_sums[4][24] ;
wire   [7:0] \level_3_sums[4][25] ;
wire   [7:0] \level_3_sums[4][26] ;
wire   [7:0] \level_3_sums[4][27] ;
wire   [7:0] \level_3_sums[4][28] ;
wire   [7:0] \level_3_sums[4][29] ;
wire   [7:0] \level_3_sums[4][30] ;
wire   [7:0] \level_3_sums[4][31] ;
wire   [7:0] \level_3_sums[5][0] ;
wire   [7:0] \level_3_sums[5][1] ;
wire   [7:0] \level_3_sums[5][2] ;
wire   [7:0] \level_3_sums[5][3] ;
wire   [7:0] \level_3_sums[5][4] ;
wire   [7:0] \level_3_sums[5][5] ;
wire   [7:0] \level_3_sums[5][6] ;
wire   [7:0] \level_3_sums[5][7] ;
wire   [7:0] \level_3_sums[5][8] ;
wire   [7:0] \level_3_sums[5][9] ;
wire   [7:0] \level_3_sums[5][10] ;
wire   [7:0] \level_3_sums[5][11] ;
wire   [7:0] \level_3_sums[5][12] ;
wire   [7:0] \level_3_sums[5][13] ;
wire   [7:0] \level_3_sums[5][14] ;
wire   [7:0] \level_3_sums[5][15] ;
wire   [7:0] \level_3_sums[5][16] ;
wire   [7:0] \level_3_sums[5][17] ;
wire   [7:0] \level_3_sums[5][18] ;
wire   [7:0] \level_3_sums[5][19] ;
wire   [7:0] \level_3_sums[5][20] ;
wire   [7:0] \level_3_sums[5][21] ;
wire   [7:0] \level_3_sums[5][22] ;
wire   [7:0] \level_3_sums[5][23] ;
wire   [7:0] \level_3_sums[5][24] ;
wire   [7:0] \level_3_sums[5][25] ;
wire   [7:0] \level_3_sums[5][26] ;
wire   [7:0] \level_3_sums[5][27] ;
wire   [7:0] \level_3_sums[5][28] ;
wire   [7:0] \level_3_sums[5][29] ;
wire   [7:0] \level_3_sums[5][30] ;
wire   [7:0] \level_3_sums[5][31] ;
wire   [7:0] \level_3_sums[6][0] ;
wire   [7:0] \level_3_sums[6][1] ;
wire   [7:0] \level_3_sums[6][2] ;
wire   [7:0] \level_3_sums[6][3] ;
wire   [7:0] \level_3_sums[6][4] ;
wire   [7:0] \level_3_sums[6][5] ;
wire   [7:0] \level_3_sums[6][6] ;
wire   [7:0] \level_3_sums[6][7] ;
wire   [7:0] \level_3_sums[6][8] ;
wire   [7:0] \level_3_sums[6][9] ;
wire   [7:0] \level_3_sums[6][10] ;
wire   [7:0] \level_3_sums[6][11] ;
wire   [7:0] \level_3_sums[6][12] ;
wire   [7:0] \level_3_sums[6][13] ;
wire   [7:0] \level_3_sums[6][14] ;
wire   [7:0] \level_3_sums[6][15] ;
wire   [7:0] \level_3_sums[6][16] ;
wire   [7:0] \level_3_sums[6][17] ;
wire   [7:0] \level_3_sums[6][18] ;
wire   [7:0] \level_3_sums[6][19] ;
wire   [7:0] \level_3_sums[6][20] ;
wire   [7:0] \level_3_sums[6][21] ;
wire   [7:0] \level_3_sums[6][22] ;
wire   [7:0] \level_3_sums[6][23] ;
wire   [7:0] \level_3_sums[6][24] ;
wire   [7:0] \level_3_sums[6][25] ;
wire   [7:0] \level_3_sums[6][26] ;
wire   [7:0] \level_3_sums[6][27] ;
wire   [7:0] \level_3_sums[6][28] ;
wire   [7:0] \level_3_sums[6][29] ;
wire   [7:0] \level_3_sums[6][30] ;
wire   [7:0] \level_3_sums[6][31] ;
wire   [7:0] \level_3_sums[7][0] ;
wire   [7:0] \level_3_sums[7][1] ;
wire   [7:0] \level_3_sums[7][2] ;
wire   [7:0] \level_3_sums[7][3] ;
wire   [7:0] \level_3_sums[7][4] ;
wire   [7:0] \level_3_sums[7][5] ;
wire   [7:0] \level_3_sums[7][6] ;
wire   [7:0] \level_3_sums[7][7] ;
wire   [7:0] \level_3_sums[7][8] ;
wire   [7:0] \level_3_sums[7][9] ;
wire   [7:0] \level_3_sums[7][10] ;
wire   [7:0] \level_3_sums[7][11] ;
wire   [7:0] \level_3_sums[7][12] ;
wire   [7:0] \level_3_sums[7][13] ;
wire   [7:0] \level_3_sums[7][14] ;
wire   [7:0] \level_3_sums[7][15] ;
wire   [7:0] \level_3_sums[7][16] ;
wire   [7:0] \level_3_sums[7][17] ;
wire   [7:0] \level_3_sums[7][18] ;
wire   [7:0] \level_3_sums[7][19] ;
wire   [7:0] \level_3_sums[7][20] ;
wire   [7:0] \level_3_sums[7][21] ;
wire   [7:0] \level_3_sums[7][22] ;
wire   [7:0] \level_3_sums[7][23] ;
wire   [7:0] \level_3_sums[7][24] ;
wire   [7:0] \level_3_sums[7][25] ;
wire   [7:0] \level_3_sums[7][26] ;
wire   [7:0] \level_3_sums[7][27] ;
wire   [7:0] \level_3_sums[7][28] ;
wire   [7:0] \level_3_sums[7][29] ;
wire   [7:0] \level_3_sums[7][30] ;
wire   [7:0] \level_3_sums[7][31] ;
wire   [7:0] \level_3_sums[8][0] ;
wire   [7:0] \level_3_sums[8][1] ;
wire   [7:0] \level_3_sums[8][2] ;
wire   [7:0] \level_3_sums[8][3] ;
wire   [7:0] \level_3_sums[8][4] ;
wire   [7:0] \level_3_sums[8][5] ;
wire   [7:0] \level_3_sums[8][6] ;
wire   [7:0] \level_3_sums[8][7] ;
wire   [7:0] \level_3_sums[8][8] ;
wire   [7:0] \level_3_sums[8][9] ;
wire   [7:0] \level_3_sums[8][10] ;
wire   [7:0] \level_3_sums[8][11] ;
wire   [7:0] \level_3_sums[8][12] ;
wire   [7:0] \level_3_sums[8][13] ;
wire   [7:0] \level_3_sums[8][14] ;
wire   [7:0] \level_3_sums[8][15] ;
wire   [7:0] \level_3_sums[8][16] ;
wire   [7:0] \level_3_sums[8][17] ;
wire   [7:0] \level_3_sums[8][18] ;
wire   [7:0] \level_3_sums[8][19] ;
wire   [7:0] \level_3_sums[8][20] ;
wire   [7:0] \level_3_sums[8][21] ;
wire   [7:0] \level_3_sums[8][22] ;
wire   [7:0] \level_3_sums[8][23] ;
wire   [7:0] \level_3_sums[8][24] ;
wire   [7:0] \level_3_sums[8][25] ;
wire   [7:0] \level_3_sums[8][26] ;
wire   [7:0] \level_3_sums[8][27] ;
wire   [7:0] \level_3_sums[8][28] ;
wire   [7:0] \level_3_sums[8][29] ;
wire   [7:0] \level_3_sums[8][30] ;
wire   [7:0] \level_3_sums[8][31] ;
wire   [7:0] \level_3_sums[9][0] ;
wire   [7:0] \level_3_sums[9][1] ;
wire   [7:0] \level_3_sums[9][2] ;
wire   [7:0] \level_3_sums[9][3] ;
wire   [7:0] \level_3_sums[9][4] ;
wire   [7:0] \level_3_sums[9][5] ;
wire   [7:0] \level_3_sums[9][6] ;
wire   [7:0] \level_3_sums[9][7] ;
wire   [7:0] \level_3_sums[9][8] ;
wire   [7:0] \level_3_sums[9][9] ;
wire   [7:0] \level_3_sums[9][10] ;
wire   [7:0] \level_3_sums[9][11] ;
wire   [7:0] \level_3_sums[9][12] ;
wire   [7:0] \level_3_sums[9][13] ;
wire   [7:0] \level_3_sums[9][14] ;
wire   [7:0] \level_3_sums[9][15] ;
wire   [7:0] \level_3_sums[9][16] ;
wire   [7:0] \level_3_sums[9][17] ;
wire   [7:0] \level_3_sums[9][18] ;
wire   [7:0] \level_3_sums[9][19] ;
wire   [7:0] \level_3_sums[9][20] ;
wire   [7:0] \level_3_sums[9][21] ;
wire   [7:0] \level_3_sums[9][22] ;
wire   [7:0] \level_3_sums[9][23] ;
wire   [7:0] \level_3_sums[9][24] ;
wire   [7:0] \level_3_sums[9][25] ;
wire   [7:0] \level_3_sums[9][26] ;
wire   [7:0] \level_3_sums[9][27] ;
wire   [7:0] \level_3_sums[9][28] ;
wire   [7:0] \level_3_sums[9][29] ;
wire   [7:0] \level_3_sums[9][30] ;
wire   [7:0] \level_3_sums[9][31] ;
wire   [7:0] \level_3_sums[10][0] ;
wire   [7:0] \level_3_sums[10][1] ;
wire   [7:0] \level_3_sums[10][2] ;
wire   [7:0] \level_3_sums[10][3] ;
wire   [7:0] \level_3_sums[10][4] ;
wire   [7:0] \level_3_sums[10][5] ;
wire   [7:0] \level_3_sums[10][6] ;
wire   [7:0] \level_3_sums[10][7] ;
wire   [7:0] \level_3_sums[10][8] ;
wire   [7:0] \level_3_sums[10][9] ;
wire   [7:0] \level_3_sums[10][10] ;
wire   [7:0] \level_3_sums[10][11] ;
wire   [7:0] \level_3_sums[10][12] ;
wire   [7:0] \level_3_sums[10][13] ;
wire   [7:0] \level_3_sums[10][14] ;
wire   [7:0] \level_3_sums[10][15] ;
wire   [7:0] \level_3_sums[10][16] ;
wire   [7:0] \level_3_sums[10][17] ;
wire   [7:0] \level_3_sums[10][18] ;
wire   [7:0] \level_3_sums[10][19] ;
wire   [7:0] \level_3_sums[10][20] ;
wire   [7:0] \level_3_sums[10][21] ;
wire   [7:0] \level_3_sums[10][22] ;
wire   [7:0] \level_3_sums[10][23] ;
wire   [7:0] \level_3_sums[10][24] ;
wire   [7:0] \level_3_sums[10][25] ;
wire   [7:0] \level_3_sums[10][26] ;
wire   [7:0] \level_3_sums[10][27] ;
wire   [7:0] \level_3_sums[10][28] ;
wire   [7:0] \level_3_sums[10][29] ;
wire   [7:0] \level_3_sums[10][30] ;
wire   [7:0] \level_3_sums[10][31] ;
wire   [7:0] \level_3_sums[11][0] ;
wire   [7:0] \level_3_sums[11][1] ;
wire   [7:0] \level_3_sums[11][2] ;
wire   [7:0] \level_3_sums[11][3] ;
wire   [7:0] \level_3_sums[11][4] ;
wire   [7:0] \level_3_sums[11][5] ;
wire   [7:0] \level_3_sums[11][6] ;
wire   [7:0] \level_3_sums[11][7] ;
wire   [7:0] \level_3_sums[11][8] ;
wire   [7:0] \level_3_sums[11][9] ;
wire   [7:0] \level_3_sums[11][10] ;
wire   [7:0] \level_3_sums[11][11] ;
wire   [7:0] \level_3_sums[11][12] ;
wire   [7:0] \level_3_sums[11][13] ;
wire   [7:0] \level_3_sums[11][14] ;
wire   [7:0] \level_3_sums[11][15] ;
wire   [7:0] \level_3_sums[11][16] ;
wire   [7:0] \level_3_sums[11][17] ;
wire   [7:0] \level_3_sums[11][18] ;
wire   [7:0] \level_3_sums[11][19] ;
wire   [7:0] \level_3_sums[11][20] ;
wire   [7:0] \level_3_sums[11][21] ;
wire   [7:0] \level_3_sums[11][22] ;
wire   [7:0] \level_3_sums[11][23] ;
wire   [7:0] \level_3_sums[11][24] ;
wire   [7:0] \level_3_sums[11][25] ;
wire   [7:0] \level_3_sums[11][26] ;
wire   [7:0] \level_3_sums[11][27] ;
wire   [7:0] \level_3_sums[11][28] ;
wire   [7:0] \level_3_sums[11][29] ;
wire   [7:0] \level_3_sums[11][30] ;
wire   [7:0] \level_3_sums[11][31] ;
wire   [7:0] \level_3_sums[12][0] ;
wire   [7:0] \level_3_sums[12][1] ;
wire   [7:0] \level_3_sums[12][2] ;
wire   [7:0] \level_3_sums[12][3] ;
wire   [7:0] \level_3_sums[12][4] ;
wire   [7:0] \level_3_sums[12][5] ;
wire   [7:0] \level_3_sums[12][6] ;
wire   [7:0] \level_3_sums[12][7] ;
wire   [7:0] \level_3_sums[12][8] ;
wire   [7:0] \level_3_sums[12][9] ;
wire   [7:0] \level_3_sums[12][10] ;
wire   [7:0] \level_3_sums[12][11] ;
wire   [7:0] \level_3_sums[12][12] ;
wire   [7:0] \level_3_sums[12][13] ;
wire   [7:0] \level_3_sums[12][14] ;
wire   [7:0] \level_3_sums[12][15] ;
wire   [7:0] \level_3_sums[12][16] ;
wire   [7:0] \level_3_sums[12][17] ;
wire   [7:0] \level_3_sums[12][18] ;
wire   [7:0] \level_3_sums[12][19] ;
wire   [7:0] \level_3_sums[12][20] ;
wire   [7:0] \level_3_sums[12][21] ;
wire   [7:0] \level_3_sums[12][22] ;
wire   [7:0] \level_3_sums[12][23] ;
wire   [7:0] \level_3_sums[12][24] ;
wire   [7:0] \level_3_sums[12][25] ;
wire   [7:0] \level_3_sums[12][26] ;
wire   [7:0] \level_3_sums[12][27] ;
wire   [7:0] \level_3_sums[12][28] ;
wire   [7:0] \level_3_sums[12][29] ;
wire   [7:0] \level_3_sums[12][30] ;
wire   [7:0] \level_3_sums[12][31] ;
wire   [7:0] \level_3_sums[13][0] ;
wire   [7:0] \level_3_sums[13][1] ;
wire   [7:0] \level_3_sums[13][2] ;
wire   [7:0] \level_3_sums[13][3] ;
wire   [7:0] \level_3_sums[13][4] ;
wire   [7:0] \level_3_sums[13][5] ;
wire   [7:0] \level_3_sums[13][6] ;
wire   [7:0] \level_3_sums[13][7] ;
wire   [7:0] \level_3_sums[13][8] ;
wire   [7:0] \level_3_sums[13][9] ;
wire   [7:0] \level_3_sums[13][10] ;
wire   [7:0] \level_3_sums[13][11] ;
wire   [7:0] \level_3_sums[13][12] ;
wire   [7:0] \level_3_sums[13][13] ;
wire   [7:0] \level_3_sums[13][14] ;
wire   [7:0] \level_3_sums[13][15] ;
wire   [7:0] \level_3_sums[13][16] ;
wire   [7:0] \level_3_sums[13][17] ;
wire   [7:0] \level_3_sums[13][18] ;
wire   [7:0] \level_3_sums[13][19] ;
wire   [7:0] \level_3_sums[13][20] ;
wire   [7:0] \level_3_sums[13][21] ;
wire   [7:0] \level_3_sums[13][22] ;
wire   [7:0] \level_3_sums[13][23] ;
wire   [7:0] \level_3_sums[13][24] ;
wire   [7:0] \level_3_sums[13][25] ;
wire   [7:0] \level_3_sums[13][26] ;
wire   [7:0] \level_3_sums[13][27] ;
wire   [7:0] \level_3_sums[13][28] ;
wire   [7:0] \level_3_sums[13][29] ;
wire   [7:0] \level_3_sums[13][30] ;
wire   [7:0] \level_3_sums[13][31] ;
wire   [7:0] \level_3_sums[14][0] ;
wire   [7:0] \level_3_sums[14][1] ;
wire   [7:0] \level_3_sums[14][2] ;
wire   [7:0] \level_3_sums[14][3] ;
wire   [7:0] \level_3_sums[14][4] ;
wire   [7:0] \level_3_sums[14][5] ;
wire   [7:0] \level_3_sums[14][6] ;
wire   [7:0] \level_3_sums[14][7] ;
wire   [7:0] \level_3_sums[14][8] ;
wire   [7:0] \level_3_sums[14][9] ;
wire   [7:0] \level_3_sums[14][10] ;
wire   [7:0] \level_3_sums[14][11] ;
wire   [7:0] \level_3_sums[14][12] ;
wire   [7:0] \level_3_sums[14][13] ;
wire   [7:0] \level_3_sums[14][14] ;
wire   [7:0] \level_3_sums[14][15] ;
wire   [7:0] \level_3_sums[14][16] ;
wire   [7:0] \level_3_sums[14][17] ;
wire   [7:0] \level_3_sums[14][18] ;
wire   [7:0] \level_3_sums[14][19] ;
wire   [7:0] \level_3_sums[14][20] ;
wire   [7:0] \level_3_sums[14][21] ;
wire   [7:0] \level_3_sums[14][22] ;
wire   [7:0] \level_3_sums[14][23] ;
wire   [7:0] \level_3_sums[14][24] ;
wire   [7:0] \level_3_sums[14][25] ;
wire   [7:0] \level_3_sums[14][26] ;
wire   [7:0] \level_3_sums[14][27] ;
wire   [7:0] \level_3_sums[14][28] ;
wire   [7:0] \level_3_sums[14][29] ;
wire   [7:0] \level_3_sums[14][30] ;
wire   [7:0] \level_3_sums[14][31] ;
wire   [7:0] \level_3_sums[15][0] ;
wire   [7:0] \level_3_sums[15][1] ;
wire   [7:0] \level_3_sums[15][2] ;
wire   [7:0] \level_3_sums[15][3] ;
wire   [7:0] \level_3_sums[15][4] ;
wire   [7:0] \level_3_sums[15][5] ;
wire   [7:0] \level_3_sums[15][6] ;
wire   [7:0] \level_3_sums[15][7] ;
wire   [7:0] \level_3_sums[15][8] ;
wire   [7:0] \level_3_sums[15][9] ;
wire   [7:0] \level_3_sums[15][10] ;
wire   [7:0] \level_3_sums[15][11] ;
wire   [7:0] \level_3_sums[15][12] ;
wire   [7:0] \level_3_sums[15][13] ;
wire   [7:0] \level_3_sums[15][14] ;
wire   [7:0] \level_3_sums[15][15] ;
wire   [7:0] \level_3_sums[15][16] ;
wire   [7:0] \level_3_sums[15][17] ;
wire   [7:0] \level_3_sums[15][18] ;
wire   [7:0] \level_3_sums[15][19] ;
wire   [7:0] \level_3_sums[15][20] ;
wire   [7:0] \level_3_sums[15][21] ;
wire   [7:0] \level_3_sums[15][22] ;
wire   [7:0] \level_3_sums[15][23] ;
wire   [7:0] \level_3_sums[15][24] ;
wire   [7:0] \level_3_sums[15][25] ;
wire   [7:0] \level_3_sums[15][26] ;
wire   [7:0] \level_3_sums[15][27] ;
wire   [7:0] \level_3_sums[15][28] ;
wire   [7:0] \level_3_sums[15][29] ;
wire   [7:0] \level_3_sums[15][30] ;
wire   [7:0] \level_3_sums[15][31] ;
wire   [7:0] \level_3_sums[16][0] ;
wire   [7:0] \level_3_sums[16][1] ;
wire   [7:0] \level_3_sums[16][2] ;
wire   [7:0] \level_3_sums[16][3] ;
wire   [7:0] \level_3_sums[16][4] ;
wire   [7:0] \level_3_sums[16][5] ;
wire   [7:0] \level_3_sums[16][6] ;
wire   [7:0] \level_3_sums[16][7] ;
wire   [7:0] \level_3_sums[16][8] ;
wire   [7:0] \level_3_sums[16][9] ;
wire   [7:0] \level_3_sums[16][10] ;
wire   [7:0] \level_3_sums[16][11] ;
wire   [7:0] \level_3_sums[16][12] ;
wire   [7:0] \level_3_sums[16][13] ;
wire   [7:0] \level_3_sums[16][14] ;
wire   [7:0] \level_3_sums[16][15] ;
wire   [7:0] \level_3_sums[16][16] ;
wire   [7:0] \level_3_sums[16][17] ;
wire   [7:0] \level_3_sums[16][18] ;
wire   [7:0] \level_3_sums[16][19] ;
wire   [7:0] \level_3_sums[16][20] ;
wire   [7:0] \level_3_sums[16][21] ;
wire   [7:0] \level_3_sums[16][22] ;
wire   [7:0] \level_3_sums[16][23] ;
wire   [7:0] \level_3_sums[16][24] ;
wire   [7:0] \level_3_sums[16][25] ;
wire   [7:0] \level_3_sums[16][26] ;
wire   [7:0] \level_3_sums[16][27] ;
wire   [7:0] \level_3_sums[16][28] ;
wire   [7:0] \level_3_sums[16][29] ;
wire   [7:0] \level_3_sums[16][30] ;
wire   [7:0] \level_3_sums[16][31] ;
wire   [7:0] \level_3_sums[17][0] ;
wire   [7:0] \level_3_sums[17][1] ;
wire   [7:0] \level_3_sums[17][2] ;
wire   [7:0] \level_3_sums[17][3] ;
wire   [7:0] \level_3_sums[17][4] ;
wire   [7:0] \level_3_sums[17][5] ;
wire   [7:0] \level_3_sums[17][6] ;
wire   [7:0] \level_3_sums[17][7] ;
wire   [7:0] \level_3_sums[17][8] ;
wire   [7:0] \level_3_sums[17][9] ;
wire   [7:0] \level_3_sums[17][10] ;
wire   [7:0] \level_3_sums[17][11] ;
wire   [7:0] \level_3_sums[17][12] ;
wire   [7:0] \level_3_sums[17][13] ;
wire   [7:0] \level_3_sums[17][14] ;
wire   [7:0] \level_3_sums[17][15] ;
wire   [7:0] \level_3_sums[17][16] ;
wire   [7:0] \level_3_sums[17][17] ;
wire   [7:0] \level_3_sums[17][18] ;
wire   [7:0] \level_3_sums[17][19] ;
wire   [7:0] \level_3_sums[17][20] ;
wire   [7:0] \level_3_sums[17][21] ;
wire   [7:0] \level_3_sums[17][22] ;
wire   [7:0] \level_3_sums[17][23] ;
wire   [7:0] \level_3_sums[17][24] ;
wire   [7:0] \level_3_sums[17][25] ;
wire   [7:0] \level_3_sums[17][26] ;
wire   [7:0] \level_3_sums[17][27] ;
wire   [7:0] \level_3_sums[17][28] ;
wire   [7:0] \level_3_sums[17][29] ;
wire   [7:0] \level_3_sums[17][30] ;
wire   [7:0] \level_3_sums[17][31] ;
wire   [7:0] \level_3_sums[18][0] ;
wire   [7:0] \level_3_sums[18][1] ;
wire   [7:0] \level_3_sums[18][2] ;
wire   [7:0] \level_3_sums[18][3] ;
wire   [7:0] \level_3_sums[18][4] ;
wire   [7:0] \level_3_sums[18][5] ;
wire   [7:0] \level_3_sums[18][6] ;
wire   [7:0] \level_3_sums[18][7] ;
wire   [7:0] \level_3_sums[18][8] ;
wire   [7:0] \level_3_sums[18][9] ;
wire   [7:0] \level_3_sums[18][10] ;
wire   [7:0] \level_3_sums[18][11] ;
wire   [7:0] \level_3_sums[18][12] ;
wire   [7:0] \level_3_sums[18][13] ;
wire   [7:0] \level_3_sums[18][14] ;
wire   [7:0] \level_3_sums[18][15] ;
wire   [7:0] \level_3_sums[18][16] ;
wire   [7:0] \level_3_sums[18][17] ;
wire   [7:0] \level_3_sums[18][18] ;
wire   [7:0] \level_3_sums[18][19] ;
wire   [7:0] \level_3_sums[18][20] ;
wire   [7:0] \level_3_sums[18][21] ;
wire   [7:0] \level_3_sums[18][22] ;
wire   [7:0] \level_3_sums[18][23] ;
wire   [7:0] \level_3_sums[18][24] ;
wire   [7:0] \level_3_sums[18][25] ;
wire   [7:0] \level_3_sums[18][26] ;
wire   [7:0] \level_3_sums[18][27] ;
wire   [7:0] \level_3_sums[18][28] ;
wire   [7:0] \level_3_sums[18][29] ;
wire   [7:0] \level_3_sums[18][30] ;
wire   [7:0] \level_3_sums[18][31] ;
wire   [7:0] \level_3_sums[19][0] ;
wire   [7:0] \level_3_sums[19][1] ;
wire   [7:0] \level_3_sums[19][2] ;
wire   [7:0] \level_3_sums[19][3] ;
wire   [7:0] \level_3_sums[19][4] ;
wire   [7:0] \level_3_sums[19][5] ;
wire   [7:0] \level_3_sums[19][6] ;
wire   [7:0] \level_3_sums[19][7] ;
wire   [7:0] \level_3_sums[19][8] ;
wire   [7:0] \level_3_sums[19][9] ;
wire   [7:0] \level_3_sums[19][10] ;
wire   [7:0] \level_3_sums[19][11] ;
wire   [7:0] \level_3_sums[19][12] ;
wire   [7:0] \level_3_sums[19][13] ;
wire   [7:0] \level_3_sums[19][14] ;
wire   [7:0] \level_3_sums[19][15] ;
wire   [7:0] \level_3_sums[19][16] ;
wire   [7:0] \level_3_sums[19][17] ;
wire   [7:0] \level_3_sums[19][18] ;
wire   [7:0] \level_3_sums[19][19] ;
wire   [7:0] \level_3_sums[19][20] ;
wire   [7:0] \level_3_sums[19][21] ;
wire   [7:0] \level_3_sums[19][22] ;
wire   [7:0] \level_3_sums[19][23] ;
wire   [7:0] \level_3_sums[19][24] ;
wire   [7:0] \level_3_sums[19][25] ;
wire   [7:0] \level_3_sums[19][26] ;
wire   [7:0] \level_3_sums[19][27] ;
wire   [7:0] \level_3_sums[19][28] ;
wire   [7:0] \level_3_sums[19][29] ;
wire   [7:0] \level_3_sums[19][30] ;
wire   [7:0] \level_3_sums[19][31] ;
wire   [6:0] \level_2_sums[0][0] ;
wire   [6:0] \level_2_sums[0][1] ;
wire   [6:0] \level_2_sums[0][2] ;
wire   [6:0] \level_2_sums[0][3] ;
wire   [6:0] \level_2_sums[0][4] ;
wire   [6:0] \level_2_sums[0][5] ;
wire   [6:0] \level_2_sums[0][6] ;
wire   [6:0] \level_2_sums[0][7] ;
wire   [6:0] \level_2_sums[0][8] ;
wire   [6:0] \level_2_sums[0][9] ;
wire   [6:0] \level_2_sums[0][10] ;
wire   [6:0] \level_2_sums[0][11] ;
wire   [6:0] \level_2_sums[0][12] ;
wire   [6:0] \level_2_sums[0][13] ;
wire   [6:0] \level_2_sums[0][14] ;
wire   [6:0] \level_2_sums[0][15] ;
wire   [6:0] \level_2_sums[0][16] ;
wire   [6:0] \level_2_sums[0][17] ;
wire   [6:0] \level_2_sums[0][18] ;
wire   [6:0] \level_2_sums[0][19] ;
wire   [6:0] \level_2_sums[0][20] ;
wire   [6:0] \level_2_sums[0][21] ;
wire   [6:0] \level_2_sums[0][22] ;
wire   [6:0] \level_2_sums[0][23] ;
wire   [6:0] \level_2_sums[0][24] ;
wire   [6:0] \level_2_sums[0][25] ;
wire   [6:0] \level_2_sums[0][26] ;
wire   [6:0] \level_2_sums[0][27] ;
wire   [6:0] \level_2_sums[0][28] ;
wire   [6:0] \level_2_sums[0][29] ;
wire   [6:0] \level_2_sums[0][30] ;
wire   [6:0] \level_2_sums[0][31] ;
wire   [6:0] \level_2_sums[0][32] ;
wire   [6:0] \level_2_sums[0][33] ;
wire   [6:0] \level_2_sums[0][34] ;
wire   [6:0] \level_2_sums[0][35] ;
wire   [6:0] \level_2_sums[0][36] ;
wire   [6:0] \level_2_sums[0][37] ;
wire   [6:0] \level_2_sums[0][38] ;
wire   [6:0] \level_2_sums[0][39] ;
wire   [6:0] \level_2_sums[0][40] ;
wire   [6:0] \level_2_sums[0][41] ;
wire   [6:0] \level_2_sums[0][42] ;
wire   [6:0] \level_2_sums[0][43] ;
wire   [6:0] \level_2_sums[0][44] ;
wire   [6:0] \level_2_sums[0][45] ;
wire   [6:0] \level_2_sums[0][46] ;
wire   [6:0] \level_2_sums[0][47] ;
wire   [6:0] \level_2_sums[0][48] ;
wire   [6:0] \level_2_sums[0][49] ;
wire   [6:0] \level_2_sums[0][50] ;
wire   [6:0] \level_2_sums[0][51] ;
wire   [6:0] \level_2_sums[0][52] ;
wire   [6:0] \level_2_sums[0][53] ;
wire   [6:0] \level_2_sums[0][54] ;
wire   [6:0] \level_2_sums[0][55] ;
wire   [6:0] \level_2_sums[0][56] ;
wire   [6:0] \level_2_sums[0][57] ;
wire   [6:0] \level_2_sums[0][58] ;
wire   [6:0] \level_2_sums[0][59] ;
wire   [6:0] \level_2_sums[0][60] ;
wire   [6:0] \level_2_sums[0][61] ;
wire   [6:0] \level_2_sums[0][62] ;
wire   [6:0] \level_2_sums[0][63] ;
wire   [6:0] \level_2_sums[1][0] ;
wire   [6:0] \level_2_sums[1][1] ;
wire   [6:0] \level_2_sums[1][2] ;
wire   [6:0] \level_2_sums[1][3] ;
wire   [6:0] \level_2_sums[1][4] ;
wire   [6:0] \level_2_sums[1][5] ;
wire   [6:0] \level_2_sums[1][6] ;
wire   [6:0] \level_2_sums[1][7] ;
wire   [6:0] \level_2_sums[1][8] ;
wire   [6:0] \level_2_sums[1][9] ;
wire   [6:0] \level_2_sums[1][10] ;
wire   [6:0] \level_2_sums[1][11] ;
wire   [6:0] \level_2_sums[1][12] ;
wire   [6:0] \level_2_sums[1][13] ;
wire   [6:0] \level_2_sums[1][14] ;
wire   [6:0] \level_2_sums[1][15] ;
wire   [6:0] \level_2_sums[1][16] ;
wire   [6:0] \level_2_sums[1][17] ;
wire   [6:0] \level_2_sums[1][18] ;
wire   [6:0] \level_2_sums[1][19] ;
wire   [6:0] \level_2_sums[1][20] ;
wire   [6:0] \level_2_sums[1][21] ;
wire   [6:0] \level_2_sums[1][22] ;
wire   [6:0] \level_2_sums[1][23] ;
wire   [6:0] \level_2_sums[1][24] ;
wire   [6:0] \level_2_sums[1][25] ;
wire   [6:0] \level_2_sums[1][26] ;
wire   [6:0] \level_2_sums[1][27] ;
wire   [6:0] \level_2_sums[1][28] ;
wire   [6:0] \level_2_sums[1][29] ;
wire   [6:0] \level_2_sums[1][30] ;
wire   [6:0] \level_2_sums[1][31] ;
wire   [6:0] \level_2_sums[1][32] ;
wire   [6:0] \level_2_sums[1][33] ;
wire   [6:0] \level_2_sums[1][34] ;
wire   [6:0] \level_2_sums[1][35] ;
wire   [6:0] \level_2_sums[1][36] ;
wire   [6:0] \level_2_sums[1][37] ;
wire   [6:0] \level_2_sums[1][38] ;
wire   [6:0] \level_2_sums[1][39] ;
wire   [6:0] \level_2_sums[1][40] ;
wire   [6:0] \level_2_sums[1][41] ;
wire   [6:0] \level_2_sums[1][42] ;
wire   [6:0] \level_2_sums[1][43] ;
wire   [6:0] \level_2_sums[1][44] ;
wire   [6:0] \level_2_sums[1][45] ;
wire   [6:0] \level_2_sums[1][46] ;
wire   [6:0] \level_2_sums[1][47] ;
wire   [6:0] \level_2_sums[1][48] ;
wire   [6:0] \level_2_sums[1][49] ;
wire   [6:0] \level_2_sums[1][50] ;
wire   [6:0] \level_2_sums[1][51] ;
wire   [6:0] \level_2_sums[1][52] ;
wire   [6:0] \level_2_sums[1][53] ;
wire   [6:0] \level_2_sums[1][54] ;
wire   [6:0] \level_2_sums[1][55] ;
wire   [6:0] \level_2_sums[1][56] ;
wire   [6:0] \level_2_sums[1][57] ;
wire   [6:0] \level_2_sums[1][58] ;
wire   [6:0] \level_2_sums[1][59] ;
wire   [6:0] \level_2_sums[1][60] ;
wire   [6:0] \level_2_sums[1][61] ;
wire   [6:0] \level_2_sums[1][62] ;
wire   [6:0] \level_2_sums[1][63] ;
wire   [6:0] \level_2_sums[2][0] ;
wire   [6:0] \level_2_sums[2][1] ;
wire   [6:0] \level_2_sums[2][2] ;
wire   [6:0] \level_2_sums[2][3] ;
wire   [6:0] \level_2_sums[2][4] ;
wire   [6:0] \level_2_sums[2][5] ;
wire   [6:0] \level_2_sums[2][6] ;
wire   [6:0] \level_2_sums[2][7] ;
wire   [6:0] \level_2_sums[2][8] ;
wire   [6:0] \level_2_sums[2][9] ;
wire   [6:0] \level_2_sums[2][10] ;
wire   [6:0] \level_2_sums[2][11] ;
wire   [6:0] \level_2_sums[2][12] ;
wire   [6:0] \level_2_sums[2][13] ;
wire   [6:0] \level_2_sums[2][14] ;
wire   [6:0] \level_2_sums[2][15] ;
wire   [6:0] \level_2_sums[2][16] ;
wire   [6:0] \level_2_sums[2][17] ;
wire   [6:0] \level_2_sums[2][18] ;
wire   [6:0] \level_2_sums[2][19] ;
wire   [6:0] \level_2_sums[2][20] ;
wire   [6:0] \level_2_sums[2][21] ;
wire   [6:0] \level_2_sums[2][22] ;
wire   [6:0] \level_2_sums[2][23] ;
wire   [6:0] \level_2_sums[2][24] ;
wire   [6:0] \level_2_sums[2][25] ;
wire   [6:0] \level_2_sums[2][26] ;
wire   [6:0] \level_2_sums[2][27] ;
wire   [6:0] \level_2_sums[2][28] ;
wire   [6:0] \level_2_sums[2][29] ;
wire   [6:0] \level_2_sums[2][30] ;
wire   [6:0] \level_2_sums[2][31] ;
wire   [6:0] \level_2_sums[2][32] ;
wire   [6:0] \level_2_sums[2][33] ;
wire   [6:0] \level_2_sums[2][34] ;
wire   [6:0] \level_2_sums[2][35] ;
wire   [6:0] \level_2_sums[2][36] ;
wire   [6:0] \level_2_sums[2][37] ;
wire   [6:0] \level_2_sums[2][38] ;
wire   [6:0] \level_2_sums[2][39] ;
wire   [6:0] \level_2_sums[2][40] ;
wire   [6:0] \level_2_sums[2][41] ;
wire   [6:0] \level_2_sums[2][42] ;
wire   [6:0] \level_2_sums[2][43] ;
wire   [6:0] \level_2_sums[2][44] ;
wire   [6:0] \level_2_sums[2][45] ;
wire   [6:0] \level_2_sums[2][46] ;
wire   [6:0] \level_2_sums[2][47] ;
wire   [6:0] \level_2_sums[2][48] ;
wire   [6:0] \level_2_sums[2][49] ;
wire   [6:0] \level_2_sums[2][50] ;
wire   [6:0] \level_2_sums[2][51] ;
wire   [6:0] \level_2_sums[2][52] ;
wire   [6:0] \level_2_sums[2][53] ;
wire   [6:0] \level_2_sums[2][54] ;
wire   [6:0] \level_2_sums[2][55] ;
wire   [6:0] \level_2_sums[2][56] ;
wire   [6:0] \level_2_sums[2][57] ;
wire   [6:0] \level_2_sums[2][58] ;
wire   [6:0] \level_2_sums[2][59] ;
wire   [6:0] \level_2_sums[2][60] ;
wire   [6:0] \level_2_sums[2][61] ;
wire   [6:0] \level_2_sums[2][62] ;
wire   [6:0] \level_2_sums[2][63] ;
wire   [6:0] \level_2_sums[3][0] ;
wire   [6:0] \level_2_sums[3][1] ;
wire   [6:0] \level_2_sums[3][2] ;
wire   [6:0] \level_2_sums[3][3] ;
wire   [6:0] \level_2_sums[3][4] ;
wire   [6:0] \level_2_sums[3][5] ;
wire   [6:0] \level_2_sums[3][6] ;
wire   [6:0] \level_2_sums[3][7] ;
wire   [6:0] \level_2_sums[3][8] ;
wire   [6:0] \level_2_sums[3][9] ;
wire   [6:0] \level_2_sums[3][10] ;
wire   [6:0] \level_2_sums[3][11] ;
wire   [6:0] \level_2_sums[3][12] ;
wire   [6:0] \level_2_sums[3][13] ;
wire   [6:0] \level_2_sums[3][14] ;
wire   [6:0] \level_2_sums[3][15] ;
wire   [6:0] \level_2_sums[3][16] ;
wire   [6:0] \level_2_sums[3][17] ;
wire   [6:0] \level_2_sums[3][18] ;
wire   [6:0] \level_2_sums[3][19] ;
wire   [6:0] \level_2_sums[3][20] ;
wire   [6:0] \level_2_sums[3][21] ;
wire   [6:0] \level_2_sums[3][22] ;
wire   [6:0] \level_2_sums[3][23] ;
wire   [6:0] \level_2_sums[3][24] ;
wire   [6:0] \level_2_sums[3][25] ;
wire   [6:0] \level_2_sums[3][26] ;
wire   [6:0] \level_2_sums[3][27] ;
wire   [6:0] \level_2_sums[3][28] ;
wire   [6:0] \level_2_sums[3][29] ;
wire   [6:0] \level_2_sums[3][30] ;
wire   [6:0] \level_2_sums[3][31] ;
wire   [6:0] \level_2_sums[3][32] ;
wire   [6:0] \level_2_sums[3][33] ;
wire   [6:0] \level_2_sums[3][34] ;
wire   [6:0] \level_2_sums[3][35] ;
wire   [6:0] \level_2_sums[3][36] ;
wire   [6:0] \level_2_sums[3][37] ;
wire   [6:0] \level_2_sums[3][38] ;
wire   [6:0] \level_2_sums[3][39] ;
wire   [6:0] \level_2_sums[3][40] ;
wire   [6:0] \level_2_sums[3][41] ;
wire   [6:0] \level_2_sums[3][42] ;
wire   [6:0] \level_2_sums[3][43] ;
wire   [6:0] \level_2_sums[3][44] ;
wire   [6:0] \level_2_sums[3][45] ;
wire   [6:0] \level_2_sums[3][46] ;
wire   [6:0] \level_2_sums[3][47] ;
wire   [6:0] \level_2_sums[3][48] ;
wire   [6:0] \level_2_sums[3][49] ;
wire   [6:0] \level_2_sums[3][50] ;
wire   [6:0] \level_2_sums[3][51] ;
wire   [6:0] \level_2_sums[3][52] ;
wire   [6:0] \level_2_sums[3][53] ;
wire   [6:0] \level_2_sums[3][54] ;
wire   [6:0] \level_2_sums[3][55] ;
wire   [6:0] \level_2_sums[3][56] ;
wire   [6:0] \level_2_sums[3][57] ;
wire   [6:0] \level_2_sums[3][58] ;
wire   [6:0] \level_2_sums[3][59] ;
wire   [6:0] \level_2_sums[3][60] ;
wire   [6:0] \level_2_sums[3][61] ;
wire   [6:0] \level_2_sums[3][62] ;
wire   [6:0] \level_2_sums[3][63] ;
wire   [6:0] \level_2_sums[4][0] ;
wire   [6:0] \level_2_sums[4][1] ;
wire   [6:0] \level_2_sums[4][2] ;
wire   [6:0] \level_2_sums[4][3] ;
wire   [6:0] \level_2_sums[4][4] ;
wire   [6:0] \level_2_sums[4][5] ;
wire   [6:0] \level_2_sums[4][6] ;
wire   [6:0] \level_2_sums[4][7] ;
wire   [6:0] \level_2_sums[4][8] ;
wire   [6:0] \level_2_sums[4][9] ;
wire   [6:0] \level_2_sums[4][10] ;
wire   [6:0] \level_2_sums[4][11] ;
wire   [6:0] \level_2_sums[4][12] ;
wire   [6:0] \level_2_sums[4][13] ;
wire   [6:0] \level_2_sums[4][14] ;
wire   [6:0] \level_2_sums[4][15] ;
wire   [6:0] \level_2_sums[4][16] ;
wire   [6:0] \level_2_sums[4][17] ;
wire   [6:0] \level_2_sums[4][18] ;
wire   [6:0] \level_2_sums[4][19] ;
wire   [6:0] \level_2_sums[4][20] ;
wire   [6:0] \level_2_sums[4][21] ;
wire   [6:0] \level_2_sums[4][22] ;
wire   [6:0] \level_2_sums[4][23] ;
wire   [6:0] \level_2_sums[4][24] ;
wire   [6:0] \level_2_sums[4][25] ;
wire   [6:0] \level_2_sums[4][26] ;
wire   [6:0] \level_2_sums[4][27] ;
wire   [6:0] \level_2_sums[4][28] ;
wire   [6:0] \level_2_sums[4][29] ;
wire   [6:0] \level_2_sums[4][30] ;
wire   [6:0] \level_2_sums[4][31] ;
wire   [6:0] \level_2_sums[4][32] ;
wire   [6:0] \level_2_sums[4][33] ;
wire   [6:0] \level_2_sums[4][34] ;
wire   [6:0] \level_2_sums[4][35] ;
wire   [6:0] \level_2_sums[4][36] ;
wire   [6:0] \level_2_sums[4][37] ;
wire   [6:0] \level_2_sums[4][38] ;
wire   [6:0] \level_2_sums[4][39] ;
wire   [6:0] \level_2_sums[4][40] ;
wire   [6:0] \level_2_sums[4][41] ;
wire   [6:0] \level_2_sums[4][42] ;
wire   [6:0] \level_2_sums[4][43] ;
wire   [6:0] \level_2_sums[4][44] ;
wire   [6:0] \level_2_sums[4][45] ;
wire   [6:0] \level_2_sums[4][46] ;
wire   [6:0] \level_2_sums[4][47] ;
wire   [6:0] \level_2_sums[4][48] ;
wire   [6:0] \level_2_sums[4][49] ;
wire   [6:0] \level_2_sums[4][50] ;
wire   [6:0] \level_2_sums[4][51] ;
wire   [6:0] \level_2_sums[4][52] ;
wire   [6:0] \level_2_sums[4][53] ;
wire   [6:0] \level_2_sums[4][54] ;
wire   [6:0] \level_2_sums[4][55] ;
wire   [6:0] \level_2_sums[4][56] ;
wire   [6:0] \level_2_sums[4][57] ;
wire   [6:0] \level_2_sums[4][58] ;
wire   [6:0] \level_2_sums[4][59] ;
wire   [6:0] \level_2_sums[4][60] ;
wire   [6:0] \level_2_sums[4][61] ;
wire   [6:0] \level_2_sums[4][62] ;
wire   [6:0] \level_2_sums[4][63] ;
wire   [6:0] \level_2_sums[5][0] ;
wire   [6:0] \level_2_sums[5][1] ;
wire   [6:0] \level_2_sums[5][2] ;
wire   [6:0] \level_2_sums[5][3] ;
wire   [6:0] \level_2_sums[5][4] ;
wire   [6:0] \level_2_sums[5][5] ;
wire   [6:0] \level_2_sums[5][6] ;
wire   [6:0] \level_2_sums[5][7] ;
wire   [6:0] \level_2_sums[5][8] ;
wire   [6:0] \level_2_sums[5][9] ;
wire   [6:0] \level_2_sums[5][10] ;
wire   [6:0] \level_2_sums[5][11] ;
wire   [6:0] \level_2_sums[5][12] ;
wire   [6:0] \level_2_sums[5][13] ;
wire   [6:0] \level_2_sums[5][14] ;
wire   [6:0] \level_2_sums[5][15] ;
wire   [6:0] \level_2_sums[5][16] ;
wire   [6:0] \level_2_sums[5][17] ;
wire   [6:0] \level_2_sums[5][18] ;
wire   [6:0] \level_2_sums[5][19] ;
wire   [6:0] \level_2_sums[5][20] ;
wire   [6:0] \level_2_sums[5][21] ;
wire   [6:0] \level_2_sums[5][22] ;
wire   [6:0] \level_2_sums[5][23] ;
wire   [6:0] \level_2_sums[5][24] ;
wire   [6:0] \level_2_sums[5][25] ;
wire   [6:0] \level_2_sums[5][26] ;
wire   [6:0] \level_2_sums[5][27] ;
wire   [6:0] \level_2_sums[5][28] ;
wire   [6:0] \level_2_sums[5][29] ;
wire   [6:0] \level_2_sums[5][30] ;
wire   [6:0] \level_2_sums[5][31] ;
wire   [6:0] \level_2_sums[5][32] ;
wire   [6:0] \level_2_sums[5][33] ;
wire   [6:0] \level_2_sums[5][34] ;
wire   [6:0] \level_2_sums[5][35] ;
wire   [6:0] \level_2_sums[5][36] ;
wire   [6:0] \level_2_sums[5][37] ;
wire   [6:0] \level_2_sums[5][38] ;
wire   [6:0] \level_2_sums[5][39] ;
wire   [6:0] \level_2_sums[5][40] ;
wire   [6:0] \level_2_sums[5][41] ;
wire   [6:0] \level_2_sums[5][42] ;
wire   [6:0] \level_2_sums[5][43] ;
wire   [6:0] \level_2_sums[5][44] ;
wire   [6:0] \level_2_sums[5][45] ;
wire   [6:0] \level_2_sums[5][46] ;
wire   [6:0] \level_2_sums[5][47] ;
wire   [6:0] \level_2_sums[5][48] ;
wire   [6:0] \level_2_sums[5][49] ;
wire   [6:0] \level_2_sums[5][50] ;
wire   [6:0] \level_2_sums[5][51] ;
wire   [6:0] \level_2_sums[5][52] ;
wire   [6:0] \level_2_sums[5][53] ;
wire   [6:0] \level_2_sums[5][54] ;
wire   [6:0] \level_2_sums[5][55] ;
wire   [6:0] \level_2_sums[5][56] ;
wire   [6:0] \level_2_sums[5][57] ;
wire   [6:0] \level_2_sums[5][58] ;
wire   [6:0] \level_2_sums[5][59] ;
wire   [6:0] \level_2_sums[5][60] ;
wire   [6:0] \level_2_sums[5][61] ;
wire   [6:0] \level_2_sums[5][62] ;
wire   [6:0] \level_2_sums[5][63] ;
wire   [6:0] \level_2_sums[6][0] ;
wire   [6:0] \level_2_sums[6][1] ;
wire   [6:0] \level_2_sums[6][2] ;
wire   [6:0] \level_2_sums[6][3] ;
wire   [6:0] \level_2_sums[6][4] ;
wire   [6:0] \level_2_sums[6][5] ;
wire   [6:0] \level_2_sums[6][6] ;
wire   [6:0] \level_2_sums[6][7] ;
wire   [6:0] \level_2_sums[6][8] ;
wire   [6:0] \level_2_sums[6][9] ;
wire   [6:0] \level_2_sums[6][10] ;
wire   [6:0] \level_2_sums[6][11] ;
wire   [6:0] \level_2_sums[6][12] ;
wire   [6:0] \level_2_sums[6][13] ;
wire   [6:0] \level_2_sums[6][14] ;
wire   [6:0] \level_2_sums[6][15] ;
wire   [6:0] \level_2_sums[6][16] ;
wire   [6:0] \level_2_sums[6][17] ;
wire   [6:0] \level_2_sums[6][18] ;
wire   [6:0] \level_2_sums[6][19] ;
wire   [6:0] \level_2_sums[6][20] ;
wire   [6:0] \level_2_sums[6][21] ;
wire   [6:0] \level_2_sums[6][22] ;
wire   [6:0] \level_2_sums[6][23] ;
wire   [6:0] \level_2_sums[6][24] ;
wire   [6:0] \level_2_sums[6][25] ;
wire   [6:0] \level_2_sums[6][26] ;
wire   [6:0] \level_2_sums[6][27] ;
wire   [6:0] \level_2_sums[6][28] ;
wire   [6:0] \level_2_sums[6][29] ;
wire   [6:0] \level_2_sums[6][30] ;
wire   [6:0] \level_2_sums[6][31] ;
wire   [6:0] \level_2_sums[6][32] ;
wire   [6:0] \level_2_sums[6][33] ;
wire   [6:0] \level_2_sums[6][34] ;
wire   [6:0] \level_2_sums[6][35] ;
wire   [6:0] \level_2_sums[6][36] ;
wire   [6:0] \level_2_sums[6][37] ;
wire   [6:0] \level_2_sums[6][38] ;
wire   [6:0] \level_2_sums[6][39] ;
wire   [6:0] \level_2_sums[6][40] ;
wire   [6:0] \level_2_sums[6][41] ;
wire   [6:0] \level_2_sums[6][42] ;
wire   [6:0] \level_2_sums[6][43] ;
wire   [6:0] \level_2_sums[6][44] ;
wire   [6:0] \level_2_sums[6][45] ;
wire   [6:0] \level_2_sums[6][46] ;
wire   [6:0] \level_2_sums[6][47] ;
wire   [6:0] \level_2_sums[6][48] ;
wire   [6:0] \level_2_sums[6][49] ;
wire   [6:0] \level_2_sums[6][50] ;
wire   [6:0] \level_2_sums[6][51] ;
wire   [6:0] \level_2_sums[6][52] ;
wire   [6:0] \level_2_sums[6][53] ;
wire   [6:0] \level_2_sums[6][54] ;
wire   [6:0] \level_2_sums[6][55] ;
wire   [6:0] \level_2_sums[6][56] ;
wire   [6:0] \level_2_sums[6][57] ;
wire   [6:0] \level_2_sums[6][58] ;
wire   [6:0] \level_2_sums[6][59] ;
wire   [6:0] \level_2_sums[6][60] ;
wire   [6:0] \level_2_sums[6][61] ;
wire   [6:0] \level_2_sums[6][62] ;
wire   [6:0] \level_2_sums[6][63] ;
wire   [6:0] \level_2_sums[7][0] ;
wire   [6:0] \level_2_sums[7][1] ;
wire   [6:0] \level_2_sums[7][2] ;
wire   [6:0] \level_2_sums[7][3] ;
wire   [6:0] \level_2_sums[7][4] ;
wire   [6:0] \level_2_sums[7][5] ;
wire   [6:0] \level_2_sums[7][6] ;
wire   [6:0] \level_2_sums[7][7] ;
wire   [6:0] \level_2_sums[7][8] ;
wire   [6:0] \level_2_sums[7][9] ;
wire   [6:0] \level_2_sums[7][10] ;
wire   [6:0] \level_2_sums[7][11] ;
wire   [6:0] \level_2_sums[7][12] ;
wire   [6:0] \level_2_sums[7][13] ;
wire   [6:0] \level_2_sums[7][14] ;
wire   [6:0] \level_2_sums[7][15] ;
wire   [6:0] \level_2_sums[7][16] ;
wire   [6:0] \level_2_sums[7][17] ;
wire   [6:0] \level_2_sums[7][18] ;
wire   [6:0] \level_2_sums[7][19] ;
wire   [6:0] \level_2_sums[7][20] ;
wire   [6:0] \level_2_sums[7][21] ;
wire   [6:0] \level_2_sums[7][22] ;
wire   [6:0] \level_2_sums[7][23] ;
wire   [6:0] \level_2_sums[7][24] ;
wire   [6:0] \level_2_sums[7][25] ;
wire   [6:0] \level_2_sums[7][26] ;
wire   [6:0] \level_2_sums[7][27] ;
wire   [6:0] \level_2_sums[7][28] ;
wire   [6:0] \level_2_sums[7][29] ;
wire   [6:0] \level_2_sums[7][30] ;
wire   [6:0] \level_2_sums[7][31] ;
wire   [6:0] \level_2_sums[7][32] ;
wire   [6:0] \level_2_sums[7][33] ;
wire   [6:0] \level_2_sums[7][34] ;
wire   [6:0] \level_2_sums[7][35] ;
wire   [6:0] \level_2_sums[7][36] ;
wire   [6:0] \level_2_sums[7][37] ;
wire   [6:0] \level_2_sums[7][38] ;
wire   [6:0] \level_2_sums[7][39] ;
wire   [6:0] \level_2_sums[7][40] ;
wire   [6:0] \level_2_sums[7][41] ;
wire   [6:0] \level_2_sums[7][42] ;
wire   [6:0] \level_2_sums[7][43] ;
wire   [6:0] \level_2_sums[7][44] ;
wire   [6:0] \level_2_sums[7][45] ;
wire   [6:0] \level_2_sums[7][46] ;
wire   [6:0] \level_2_sums[7][47] ;
wire   [6:0] \level_2_sums[7][48] ;
wire   [6:0] \level_2_sums[7][49] ;
wire   [6:0] \level_2_sums[7][50] ;
wire   [6:0] \level_2_sums[7][51] ;
wire   [6:0] \level_2_sums[7][52] ;
wire   [6:0] \level_2_sums[7][53] ;
wire   [6:0] \level_2_sums[7][54] ;
wire   [6:0] \level_2_sums[7][55] ;
wire   [6:0] \level_2_sums[7][56] ;
wire   [6:0] \level_2_sums[7][57] ;
wire   [6:0] \level_2_sums[7][58] ;
wire   [6:0] \level_2_sums[7][59] ;
wire   [6:0] \level_2_sums[7][60] ;
wire   [6:0] \level_2_sums[7][61] ;
wire   [6:0] \level_2_sums[7][62] ;
wire   [6:0] \level_2_sums[7][63] ;
wire   [6:0] \level_2_sums[8][0] ;
wire   [6:0] \level_2_sums[8][1] ;
wire   [6:0] \level_2_sums[8][2] ;
wire   [6:0] \level_2_sums[8][3] ;
wire   [6:0] \level_2_sums[8][4] ;
wire   [6:0] \level_2_sums[8][5] ;
wire   [6:0] \level_2_sums[8][6] ;
wire   [6:0] \level_2_sums[8][7] ;
wire   [6:0] \level_2_sums[8][8] ;
wire   [6:0] \level_2_sums[8][9] ;
wire   [6:0] \level_2_sums[8][10] ;
wire   [6:0] \level_2_sums[8][11] ;
wire   [6:0] \level_2_sums[8][12] ;
wire   [6:0] \level_2_sums[8][13] ;
wire   [6:0] \level_2_sums[8][14] ;
wire   [6:0] \level_2_sums[8][15] ;
wire   [6:0] \level_2_sums[8][16] ;
wire   [6:0] \level_2_sums[8][17] ;
wire   [6:0] \level_2_sums[8][18] ;
wire   [6:0] \level_2_sums[8][19] ;
wire   [6:0] \level_2_sums[8][20] ;
wire   [6:0] \level_2_sums[8][21] ;
wire   [6:0] \level_2_sums[8][22] ;
wire   [6:0] \level_2_sums[8][23] ;
wire   [6:0] \level_2_sums[8][24] ;
wire   [6:0] \level_2_sums[8][25] ;
wire   [6:0] \level_2_sums[8][26] ;
wire   [6:0] \level_2_sums[8][27] ;
wire   [6:0] \level_2_sums[8][28] ;
wire   [6:0] \level_2_sums[8][29] ;
wire   [6:0] \level_2_sums[8][30] ;
wire   [6:0] \level_2_sums[8][31] ;
wire   [6:0] \level_2_sums[8][32] ;
wire   [6:0] \level_2_sums[8][33] ;
wire   [6:0] \level_2_sums[8][34] ;
wire   [6:0] \level_2_sums[8][35] ;
wire   [6:0] \level_2_sums[8][36] ;
wire   [6:0] \level_2_sums[8][37] ;
wire   [6:0] \level_2_sums[8][38] ;
wire   [6:0] \level_2_sums[8][39] ;
wire   [6:0] \level_2_sums[8][40] ;
wire   [6:0] \level_2_sums[8][41] ;
wire   [6:0] \level_2_sums[8][42] ;
wire   [6:0] \level_2_sums[8][43] ;
wire   [6:0] \level_2_sums[8][44] ;
wire   [6:0] \level_2_sums[8][45] ;
wire   [6:0] \level_2_sums[8][46] ;
wire   [6:0] \level_2_sums[8][47] ;
wire   [6:0] \level_2_sums[8][48] ;
wire   [6:0] \level_2_sums[8][49] ;
wire   [6:0] \level_2_sums[8][50] ;
wire   [6:0] \level_2_sums[8][51] ;
wire   [6:0] \level_2_sums[8][52] ;
wire   [6:0] \level_2_sums[8][53] ;
wire   [6:0] \level_2_sums[8][54] ;
wire   [6:0] \level_2_sums[8][55] ;
wire   [6:0] \level_2_sums[8][56] ;
wire   [6:0] \level_2_sums[8][57] ;
wire   [6:0] \level_2_sums[8][58] ;
wire   [6:0] \level_2_sums[8][59] ;
wire   [6:0] \level_2_sums[8][60] ;
wire   [6:0] \level_2_sums[8][61] ;
wire   [6:0] \level_2_sums[8][62] ;
wire   [6:0] \level_2_sums[8][63] ;
wire   [6:0] \level_2_sums[9][0] ;
wire   [6:0] \level_2_sums[9][1] ;
wire   [6:0] \level_2_sums[9][2] ;
wire   [6:0] \level_2_sums[9][3] ;
wire   [6:0] \level_2_sums[9][4] ;
wire   [6:0] \level_2_sums[9][5] ;
wire   [6:0] \level_2_sums[9][6] ;
wire   [6:0] \level_2_sums[9][7] ;
wire   [6:0] \level_2_sums[9][8] ;
wire   [6:0] \level_2_sums[9][9] ;
wire   [6:0] \level_2_sums[9][10] ;
wire   [6:0] \level_2_sums[9][11] ;
wire   [6:0] \level_2_sums[9][12] ;
wire   [6:0] \level_2_sums[9][13] ;
wire   [6:0] \level_2_sums[9][14] ;
wire   [6:0] \level_2_sums[9][15] ;
wire   [6:0] \level_2_sums[9][16] ;
wire   [6:0] \level_2_sums[9][17] ;
wire   [6:0] \level_2_sums[9][18] ;
wire   [6:0] \level_2_sums[9][19] ;
wire   [6:0] \level_2_sums[9][20] ;
wire   [6:0] \level_2_sums[9][21] ;
wire   [6:0] \level_2_sums[9][22] ;
wire   [6:0] \level_2_sums[9][23] ;
wire   [6:0] \level_2_sums[9][24] ;
wire   [6:0] \level_2_sums[9][25] ;
wire   [6:0] \level_2_sums[9][26] ;
wire   [6:0] \level_2_sums[9][27] ;
wire   [6:0] \level_2_sums[9][28] ;
wire   [6:0] \level_2_sums[9][29] ;
wire   [6:0] \level_2_sums[9][30] ;
wire   [6:0] \level_2_sums[9][31] ;
wire   [6:0] \level_2_sums[9][32] ;
wire   [6:0] \level_2_sums[9][33] ;
wire   [6:0] \level_2_sums[9][34] ;
wire   [6:0] \level_2_sums[9][35] ;
wire   [6:0] \level_2_sums[9][36] ;
wire   [6:0] \level_2_sums[9][37] ;
wire   [6:0] \level_2_sums[9][38] ;
wire   [6:0] \level_2_sums[9][39] ;
wire   [6:0] \level_2_sums[9][40] ;
wire   [6:0] \level_2_sums[9][41] ;
wire   [6:0] \level_2_sums[9][42] ;
wire   [6:0] \level_2_sums[9][43] ;
wire   [6:0] \level_2_sums[9][44] ;
wire   [6:0] \level_2_sums[9][45] ;
wire   [6:0] \level_2_sums[9][46] ;
wire   [6:0] \level_2_sums[9][47] ;
wire   [6:0] \level_2_sums[9][48] ;
wire   [6:0] \level_2_sums[9][49] ;
wire   [6:0] \level_2_sums[9][50] ;
wire   [6:0] \level_2_sums[9][51] ;
wire   [6:0] \level_2_sums[9][52] ;
wire   [6:0] \level_2_sums[9][53] ;
wire   [6:0] \level_2_sums[9][54] ;
wire   [6:0] \level_2_sums[9][55] ;
wire   [6:0] \level_2_sums[9][56] ;
wire   [6:0] \level_2_sums[9][57] ;
wire   [6:0] \level_2_sums[9][58] ;
wire   [6:0] \level_2_sums[9][59] ;
wire   [6:0] \level_2_sums[9][60] ;
wire   [6:0] \level_2_sums[9][61] ;
wire   [6:0] \level_2_sums[9][62] ;
wire   [6:0] \level_2_sums[9][63] ;
wire   [6:0] \level_2_sums[10][0] ;
wire   [6:0] \level_2_sums[10][1] ;
wire   [6:0] \level_2_sums[10][2] ;
wire   [6:0] \level_2_sums[10][3] ;
wire   [6:0] \level_2_sums[10][4] ;
wire   [6:0] \level_2_sums[10][5] ;
wire   [6:0] \level_2_sums[10][6] ;
wire   [6:0] \level_2_sums[10][7] ;
wire   [6:0] \level_2_sums[10][8] ;
wire   [6:0] \level_2_sums[10][9] ;
wire   [6:0] \level_2_sums[10][10] ;
wire   [6:0] \level_2_sums[10][11] ;
wire   [6:0] \level_2_sums[10][12] ;
wire   [6:0] \level_2_sums[10][13] ;
wire   [6:0] \level_2_sums[10][14] ;
wire   [6:0] \level_2_sums[10][15] ;
wire   [6:0] \level_2_sums[10][16] ;
wire   [6:0] \level_2_sums[10][17] ;
wire   [6:0] \level_2_sums[10][18] ;
wire   [6:0] \level_2_sums[10][19] ;
wire   [6:0] \level_2_sums[10][20] ;
wire   [6:0] \level_2_sums[10][21] ;
wire   [6:0] \level_2_sums[10][22] ;
wire   [6:0] \level_2_sums[10][23] ;
wire   [6:0] \level_2_sums[10][24] ;
wire   [6:0] \level_2_sums[10][25] ;
wire   [6:0] \level_2_sums[10][26] ;
wire   [6:0] \level_2_sums[10][27] ;
wire   [6:0] \level_2_sums[10][28] ;
wire   [6:0] \level_2_sums[10][29] ;
wire   [6:0] \level_2_sums[10][30] ;
wire   [6:0] \level_2_sums[10][31] ;
wire   [6:0] \level_2_sums[10][32] ;
wire   [6:0] \level_2_sums[10][33] ;
wire   [6:0] \level_2_sums[10][34] ;
wire   [6:0] \level_2_sums[10][35] ;
wire   [6:0] \level_2_sums[10][36] ;
wire   [6:0] \level_2_sums[10][37] ;
wire   [6:0] \level_2_sums[10][38] ;
wire   [6:0] \level_2_sums[10][39] ;
wire   [6:0] \level_2_sums[10][40] ;
wire   [6:0] \level_2_sums[10][41] ;
wire   [6:0] \level_2_sums[10][42] ;
wire   [6:0] \level_2_sums[10][43] ;
wire   [6:0] \level_2_sums[10][44] ;
wire   [6:0] \level_2_sums[10][45] ;
wire   [6:0] \level_2_sums[10][46] ;
wire   [6:0] \level_2_sums[10][47] ;
wire   [6:0] \level_2_sums[10][48] ;
wire   [6:0] \level_2_sums[10][49] ;
wire   [6:0] \level_2_sums[10][50] ;
wire   [6:0] \level_2_sums[10][51] ;
wire   [6:0] \level_2_sums[10][52] ;
wire   [6:0] \level_2_sums[10][53] ;
wire   [6:0] \level_2_sums[10][54] ;
wire   [6:0] \level_2_sums[10][55] ;
wire   [6:0] \level_2_sums[10][56] ;
wire   [6:0] \level_2_sums[10][57] ;
wire   [6:0] \level_2_sums[10][58] ;
wire   [6:0] \level_2_sums[10][59] ;
wire   [6:0] \level_2_sums[10][60] ;
wire   [6:0] \level_2_sums[10][61] ;
wire   [6:0] \level_2_sums[10][62] ;
wire   [6:0] \level_2_sums[10][63] ;
wire   [6:0] \level_2_sums[11][0] ;
wire   [6:0] \level_2_sums[11][1] ;
wire   [6:0] \level_2_sums[11][2] ;
wire   [6:0] \level_2_sums[11][3] ;
wire   [6:0] \level_2_sums[11][4] ;
wire   [6:0] \level_2_sums[11][5] ;
wire   [6:0] \level_2_sums[11][6] ;
wire   [6:0] \level_2_sums[11][7] ;
wire   [6:0] \level_2_sums[11][8] ;
wire   [6:0] \level_2_sums[11][9] ;
wire   [6:0] \level_2_sums[11][10] ;
wire   [6:0] \level_2_sums[11][11] ;
wire   [6:0] \level_2_sums[11][12] ;
wire   [6:0] \level_2_sums[11][13] ;
wire   [6:0] \level_2_sums[11][14] ;
wire   [6:0] \level_2_sums[11][15] ;
wire   [6:0] \level_2_sums[11][16] ;
wire   [6:0] \level_2_sums[11][17] ;
wire   [6:0] \level_2_sums[11][18] ;
wire   [6:0] \level_2_sums[11][19] ;
wire   [6:0] \level_2_sums[11][20] ;
wire   [6:0] \level_2_sums[11][21] ;
wire   [6:0] \level_2_sums[11][22] ;
wire   [6:0] \level_2_sums[11][23] ;
wire   [6:0] \level_2_sums[11][24] ;
wire   [6:0] \level_2_sums[11][25] ;
wire   [6:0] \level_2_sums[11][26] ;
wire   [6:0] \level_2_sums[11][27] ;
wire   [6:0] \level_2_sums[11][28] ;
wire   [6:0] \level_2_sums[11][29] ;
wire   [6:0] \level_2_sums[11][30] ;
wire   [6:0] \level_2_sums[11][31] ;
wire   [6:0] \level_2_sums[11][32] ;
wire   [6:0] \level_2_sums[11][33] ;
wire   [6:0] \level_2_sums[11][34] ;
wire   [6:0] \level_2_sums[11][35] ;
wire   [6:0] \level_2_sums[11][36] ;
wire   [6:0] \level_2_sums[11][37] ;
wire   [6:0] \level_2_sums[11][38] ;
wire   [6:0] \level_2_sums[11][39] ;
wire   [6:0] \level_2_sums[11][40] ;
wire   [6:0] \level_2_sums[11][41] ;
wire   [6:0] \level_2_sums[11][42] ;
wire   [6:0] \level_2_sums[11][43] ;
wire   [6:0] \level_2_sums[11][44] ;
wire   [6:0] \level_2_sums[11][45] ;
wire   [6:0] \level_2_sums[11][46] ;
wire   [6:0] \level_2_sums[11][47] ;
wire   [6:0] \level_2_sums[11][48] ;
wire   [6:0] \level_2_sums[11][49] ;
wire   [6:0] \level_2_sums[11][50] ;
wire   [6:0] \level_2_sums[11][51] ;
wire   [6:0] \level_2_sums[11][52] ;
wire   [6:0] \level_2_sums[11][53] ;
wire   [6:0] \level_2_sums[11][54] ;
wire   [6:0] \level_2_sums[11][55] ;
wire   [6:0] \level_2_sums[11][56] ;
wire   [6:0] \level_2_sums[11][57] ;
wire   [6:0] \level_2_sums[11][58] ;
wire   [6:0] \level_2_sums[11][59] ;
wire   [6:0] \level_2_sums[11][60] ;
wire   [6:0] \level_2_sums[11][61] ;
wire   [6:0] \level_2_sums[11][62] ;
wire   [6:0] \level_2_sums[11][63] ;
wire   [6:0] \level_2_sums[12][0] ;
wire   [6:0] \level_2_sums[12][1] ;
wire   [6:0] \level_2_sums[12][2] ;
wire   [6:0] \level_2_sums[12][3] ;
wire   [6:0] \level_2_sums[12][4] ;
wire   [6:0] \level_2_sums[12][5] ;
wire   [6:0] \level_2_sums[12][6] ;
wire   [6:0] \level_2_sums[12][7] ;
wire   [6:0] \level_2_sums[12][8] ;
wire   [6:0] \level_2_sums[12][9] ;
wire   [6:0] \level_2_sums[12][10] ;
wire   [6:0] \level_2_sums[12][11] ;
wire   [6:0] \level_2_sums[12][12] ;
wire   [6:0] \level_2_sums[12][13] ;
wire   [6:0] \level_2_sums[12][14] ;
wire   [6:0] \level_2_sums[12][15] ;
wire   [6:0] \level_2_sums[12][16] ;
wire   [6:0] \level_2_sums[12][17] ;
wire   [6:0] \level_2_sums[12][18] ;
wire   [6:0] \level_2_sums[12][19] ;
wire   [6:0] \level_2_sums[12][20] ;
wire   [6:0] \level_2_sums[12][21] ;
wire   [6:0] \level_2_sums[12][22] ;
wire   [6:0] \level_2_sums[12][23] ;
wire   [6:0] \level_2_sums[12][24] ;
wire   [6:0] \level_2_sums[12][25] ;
wire   [6:0] \level_2_sums[12][26] ;
wire   [6:0] \level_2_sums[12][27] ;
wire   [6:0] \level_2_sums[12][28] ;
wire   [6:0] \level_2_sums[12][29] ;
wire   [6:0] \level_2_sums[12][30] ;
wire   [6:0] \level_2_sums[12][31] ;
wire   [6:0] \level_2_sums[12][32] ;
wire   [6:0] \level_2_sums[12][33] ;
wire   [6:0] \level_2_sums[12][34] ;
wire   [6:0] \level_2_sums[12][35] ;
wire   [6:0] \level_2_sums[12][36] ;
wire   [6:0] \level_2_sums[12][37] ;
wire   [6:0] \level_2_sums[12][38] ;
wire   [6:0] \level_2_sums[12][39] ;
wire   [6:0] \level_2_sums[12][40] ;
wire   [6:0] \level_2_sums[12][41] ;
wire   [6:0] \level_2_sums[12][42] ;
wire   [6:0] \level_2_sums[12][43] ;
wire   [6:0] \level_2_sums[12][44] ;
wire   [6:0] \level_2_sums[12][45] ;
wire   [6:0] \level_2_sums[12][46] ;
wire   [6:0] \level_2_sums[12][47] ;
wire   [6:0] \level_2_sums[12][48] ;
wire   [6:0] \level_2_sums[12][49] ;
wire   [6:0] \level_2_sums[12][50] ;
wire   [6:0] \level_2_sums[12][51] ;
wire   [6:0] \level_2_sums[12][52] ;
wire   [6:0] \level_2_sums[12][53] ;
wire   [6:0] \level_2_sums[12][54] ;
wire   [6:0] \level_2_sums[12][55] ;
wire   [6:0] \level_2_sums[12][56] ;
wire   [6:0] \level_2_sums[12][57] ;
wire   [6:0] \level_2_sums[12][58] ;
wire   [6:0] \level_2_sums[12][59] ;
wire   [6:0] \level_2_sums[12][60] ;
wire   [6:0] \level_2_sums[12][61] ;
wire   [6:0] \level_2_sums[12][62] ;
wire   [6:0] \level_2_sums[12][63] ;
wire   [6:0] \level_2_sums[13][0] ;
wire   [6:0] \level_2_sums[13][1] ;
wire   [6:0] \level_2_sums[13][2] ;
wire   [6:0] \level_2_sums[13][3] ;
wire   [6:0] \level_2_sums[13][4] ;
wire   [6:0] \level_2_sums[13][5] ;
wire   [6:0] \level_2_sums[13][6] ;
wire   [6:0] \level_2_sums[13][7] ;
wire   [6:0] \level_2_sums[13][8] ;
wire   [6:0] \level_2_sums[13][9] ;
wire   [6:0] \level_2_sums[13][10] ;
wire   [6:0] \level_2_sums[13][11] ;
wire   [6:0] \level_2_sums[13][12] ;
wire   [6:0] \level_2_sums[13][13] ;
wire   [6:0] \level_2_sums[13][14] ;
wire   [6:0] \level_2_sums[13][15] ;
wire   [6:0] \level_2_sums[13][16] ;
wire   [6:0] \level_2_sums[13][17] ;
wire   [6:0] \level_2_sums[13][18] ;
wire   [6:0] \level_2_sums[13][19] ;
wire   [6:0] \level_2_sums[13][20] ;
wire   [6:0] \level_2_sums[13][21] ;
wire   [6:0] \level_2_sums[13][22] ;
wire   [6:0] \level_2_sums[13][23] ;
wire   [6:0] \level_2_sums[13][24] ;
wire   [6:0] \level_2_sums[13][25] ;
wire   [6:0] \level_2_sums[13][26] ;
wire   [6:0] \level_2_sums[13][27] ;
wire   [6:0] \level_2_sums[13][28] ;
wire   [6:0] \level_2_sums[13][29] ;
wire   [6:0] \level_2_sums[13][30] ;
wire   [6:0] \level_2_sums[13][31] ;
wire   [6:0] \level_2_sums[13][32] ;
wire   [6:0] \level_2_sums[13][33] ;
wire   [6:0] \level_2_sums[13][34] ;
wire   [6:0] \level_2_sums[13][35] ;
wire   [6:0] \level_2_sums[13][36] ;
wire   [6:0] \level_2_sums[13][37] ;
wire   [6:0] \level_2_sums[13][38] ;
wire   [6:0] \level_2_sums[13][39] ;
wire   [6:0] \level_2_sums[13][40] ;
wire   [6:0] \level_2_sums[13][41] ;
wire   [6:0] \level_2_sums[13][42] ;
wire   [6:0] \level_2_sums[13][43] ;
wire   [6:0] \level_2_sums[13][44] ;
wire   [6:0] \level_2_sums[13][45] ;
wire   [6:0] \level_2_sums[13][46] ;
wire   [6:0] \level_2_sums[13][47] ;
wire   [6:0] \level_2_sums[13][48] ;
wire   [6:0] \level_2_sums[13][49] ;
wire   [6:0] \level_2_sums[13][50] ;
wire   [6:0] \level_2_sums[13][51] ;
wire   [6:0] \level_2_sums[13][52] ;
wire   [6:0] \level_2_sums[13][53] ;
wire   [6:0] \level_2_sums[13][54] ;
wire   [6:0] \level_2_sums[13][55] ;
wire   [6:0] \level_2_sums[13][56] ;
wire   [6:0] \level_2_sums[13][57] ;
wire   [6:0] \level_2_sums[13][58] ;
wire   [6:0] \level_2_sums[13][59] ;
wire   [6:0] \level_2_sums[13][60] ;
wire   [6:0] \level_2_sums[13][61] ;
wire   [6:0] \level_2_sums[13][62] ;
wire   [6:0] \level_2_sums[13][63] ;
wire   [6:0] \level_2_sums[14][0] ;
wire   [6:0] \level_2_sums[14][1] ;
wire   [6:0] \level_2_sums[14][2] ;
wire   [6:0] \level_2_sums[14][3] ;
wire   [6:0] \level_2_sums[14][4] ;
wire   [6:0] \level_2_sums[14][5] ;
wire   [6:0] \level_2_sums[14][6] ;
wire   [6:0] \level_2_sums[14][7] ;
wire   [6:0] \level_2_sums[14][8] ;
wire   [6:0] \level_2_sums[14][9] ;
wire   [6:0] \level_2_sums[14][10] ;
wire   [6:0] \level_2_sums[14][11] ;
wire   [6:0] \level_2_sums[14][12] ;
wire   [6:0] \level_2_sums[14][13] ;
wire   [6:0] \level_2_sums[14][14] ;
wire   [6:0] \level_2_sums[14][15] ;
wire   [6:0] \level_2_sums[14][16] ;
wire   [6:0] \level_2_sums[14][17] ;
wire   [6:0] \level_2_sums[14][18] ;
wire   [6:0] \level_2_sums[14][19] ;
wire   [6:0] \level_2_sums[14][20] ;
wire   [6:0] \level_2_sums[14][21] ;
wire   [6:0] \level_2_sums[14][22] ;
wire   [6:0] \level_2_sums[14][23] ;
wire   [6:0] \level_2_sums[14][24] ;
wire   [6:0] \level_2_sums[14][25] ;
wire   [6:0] \level_2_sums[14][26] ;
wire   [6:0] \level_2_sums[14][27] ;
wire   [6:0] \level_2_sums[14][28] ;
wire   [6:0] \level_2_sums[14][29] ;
wire   [6:0] \level_2_sums[14][30] ;
wire   [6:0] \level_2_sums[14][31] ;
wire   [6:0] \level_2_sums[14][32] ;
wire   [6:0] \level_2_sums[14][33] ;
wire   [6:0] \level_2_sums[14][34] ;
wire   [6:0] \level_2_sums[14][35] ;
wire   [6:0] \level_2_sums[14][36] ;
wire   [6:0] \level_2_sums[14][37] ;
wire   [6:0] \level_2_sums[14][38] ;
wire   [6:0] \level_2_sums[14][39] ;
wire   [6:0] \level_2_sums[14][40] ;
wire   [6:0] \level_2_sums[14][41] ;
wire   [6:0] \level_2_sums[14][42] ;
wire   [6:0] \level_2_sums[14][43] ;
wire   [6:0] \level_2_sums[14][44] ;
wire   [6:0] \level_2_sums[14][45] ;
wire   [6:0] \level_2_sums[14][46] ;
wire   [6:0] \level_2_sums[14][47] ;
wire   [6:0] \level_2_sums[14][48] ;
wire   [6:0] \level_2_sums[14][49] ;
wire   [6:0] \level_2_sums[14][50] ;
wire   [6:0] \level_2_sums[14][51] ;
wire   [6:0] \level_2_sums[14][52] ;
wire   [6:0] \level_2_sums[14][53] ;
wire   [6:0] \level_2_sums[14][54] ;
wire   [6:0] \level_2_sums[14][55] ;
wire   [6:0] \level_2_sums[14][56] ;
wire   [6:0] \level_2_sums[14][57] ;
wire   [6:0] \level_2_sums[14][58] ;
wire   [6:0] \level_2_sums[14][59] ;
wire   [6:0] \level_2_sums[14][60] ;
wire   [6:0] \level_2_sums[14][61] ;
wire   [6:0] \level_2_sums[14][62] ;
wire   [6:0] \level_2_sums[14][63] ;
wire   [6:0] \level_2_sums[15][0] ;
wire   [6:0] \level_2_sums[15][1] ;
wire   [6:0] \level_2_sums[15][2] ;
wire   [6:0] \level_2_sums[15][3] ;
wire   [6:0] \level_2_sums[15][4] ;
wire   [6:0] \level_2_sums[15][5] ;
wire   [6:0] \level_2_sums[15][6] ;
wire   [6:0] \level_2_sums[15][7] ;
wire   [6:0] \level_2_sums[15][8] ;
wire   [6:0] \level_2_sums[15][9] ;
wire   [6:0] \level_2_sums[15][10] ;
wire   [6:0] \level_2_sums[15][11] ;
wire   [6:0] \level_2_sums[15][12] ;
wire   [6:0] \level_2_sums[15][13] ;
wire   [6:0] \level_2_sums[15][14] ;
wire   [6:0] \level_2_sums[15][15] ;
wire   [6:0] \level_2_sums[15][16] ;
wire   [6:0] \level_2_sums[15][17] ;
wire   [6:0] \level_2_sums[15][18] ;
wire   [6:0] \level_2_sums[15][19] ;
wire   [6:0] \level_2_sums[15][20] ;
wire   [6:0] \level_2_sums[15][21] ;
wire   [6:0] \level_2_sums[15][22] ;
wire   [6:0] \level_2_sums[15][23] ;
wire   [6:0] \level_2_sums[15][24] ;
wire   [6:0] \level_2_sums[15][25] ;
wire   [6:0] \level_2_sums[15][26] ;
wire   [6:0] \level_2_sums[15][27] ;
wire   [6:0] \level_2_sums[15][28] ;
wire   [6:0] \level_2_sums[15][29] ;
wire   [6:0] \level_2_sums[15][30] ;
wire   [6:0] \level_2_sums[15][31] ;
wire   [6:0] \level_2_sums[15][32] ;
wire   [6:0] \level_2_sums[15][33] ;
wire   [6:0] \level_2_sums[15][34] ;
wire   [6:0] \level_2_sums[15][35] ;
wire   [6:0] \level_2_sums[15][36] ;
wire   [6:0] \level_2_sums[15][37] ;
wire   [6:0] \level_2_sums[15][38] ;
wire   [6:0] \level_2_sums[15][39] ;
wire   [6:0] \level_2_sums[15][40] ;
wire   [6:0] \level_2_sums[15][41] ;
wire   [6:0] \level_2_sums[15][42] ;
wire   [6:0] \level_2_sums[15][43] ;
wire   [6:0] \level_2_sums[15][44] ;
wire   [6:0] \level_2_sums[15][45] ;
wire   [6:0] \level_2_sums[15][46] ;
wire   [6:0] \level_2_sums[15][47] ;
wire   [6:0] \level_2_sums[15][48] ;
wire   [6:0] \level_2_sums[15][49] ;
wire   [6:0] \level_2_sums[15][50] ;
wire   [6:0] \level_2_sums[15][51] ;
wire   [6:0] \level_2_sums[15][52] ;
wire   [6:0] \level_2_sums[15][53] ;
wire   [6:0] \level_2_sums[15][54] ;
wire   [6:0] \level_2_sums[15][55] ;
wire   [6:0] \level_2_sums[15][56] ;
wire   [6:0] \level_2_sums[15][57] ;
wire   [6:0] \level_2_sums[15][58] ;
wire   [6:0] \level_2_sums[15][59] ;
wire   [6:0] \level_2_sums[15][60] ;
wire   [6:0] \level_2_sums[15][61] ;
wire   [6:0] \level_2_sums[15][62] ;
wire   [6:0] \level_2_sums[15][63] ;
wire   [6:0] \level_2_sums[16][0] ;
wire   [6:0] \level_2_sums[16][1] ;
wire   [6:0] \level_2_sums[16][2] ;
wire   [6:0] \level_2_sums[16][3] ;
wire   [6:0] \level_2_sums[16][4] ;
wire   [6:0] \level_2_sums[16][5] ;
wire   [6:0] \level_2_sums[16][6] ;
wire   [6:0] \level_2_sums[16][7] ;
wire   [6:0] \level_2_sums[16][8] ;
wire   [6:0] \level_2_sums[16][9] ;
wire   [6:0] \level_2_sums[16][10] ;
wire   [6:0] \level_2_sums[16][11] ;
wire   [6:0] \level_2_sums[16][12] ;
wire   [6:0] \level_2_sums[16][13] ;
wire   [6:0] \level_2_sums[16][14] ;
wire   [6:0] \level_2_sums[16][15] ;
wire   [6:0] \level_2_sums[16][16] ;
wire   [6:0] \level_2_sums[16][17] ;
wire   [6:0] \level_2_sums[16][18] ;
wire   [6:0] \level_2_sums[16][19] ;
wire   [6:0] \level_2_sums[16][20] ;
wire   [6:0] \level_2_sums[16][21] ;
wire   [6:0] \level_2_sums[16][22] ;
wire   [6:0] \level_2_sums[16][23] ;
wire   [6:0] \level_2_sums[16][24] ;
wire   [6:0] \level_2_sums[16][25] ;
wire   [6:0] \level_2_sums[16][26] ;
wire   [6:0] \level_2_sums[16][27] ;
wire   [6:0] \level_2_sums[16][28] ;
wire   [6:0] \level_2_sums[16][29] ;
wire   [6:0] \level_2_sums[16][30] ;
wire   [6:0] \level_2_sums[16][31] ;
wire   [6:0] \level_2_sums[16][32] ;
wire   [6:0] \level_2_sums[16][33] ;
wire   [6:0] \level_2_sums[16][34] ;
wire   [6:0] \level_2_sums[16][35] ;
wire   [6:0] \level_2_sums[16][36] ;
wire   [6:0] \level_2_sums[16][37] ;
wire   [6:0] \level_2_sums[16][38] ;
wire   [6:0] \level_2_sums[16][39] ;
wire   [6:0] \level_2_sums[16][40] ;
wire   [6:0] \level_2_sums[16][41] ;
wire   [6:0] \level_2_sums[16][42] ;
wire   [6:0] \level_2_sums[16][43] ;
wire   [6:0] \level_2_sums[16][44] ;
wire   [6:0] \level_2_sums[16][45] ;
wire   [6:0] \level_2_sums[16][46] ;
wire   [6:0] \level_2_sums[16][47] ;
wire   [6:0] \level_2_sums[16][48] ;
wire   [6:0] \level_2_sums[16][49] ;
wire   [6:0] \level_2_sums[16][50] ;
wire   [6:0] \level_2_sums[16][51] ;
wire   [6:0] \level_2_sums[16][52] ;
wire   [6:0] \level_2_sums[16][53] ;
wire   [6:0] \level_2_sums[16][54] ;
wire   [6:0] \level_2_sums[16][55] ;
wire   [6:0] \level_2_sums[16][56] ;
wire   [6:0] \level_2_sums[16][57] ;
wire   [6:0] \level_2_sums[16][58] ;
wire   [6:0] \level_2_sums[16][59] ;
wire   [6:0] \level_2_sums[16][60] ;
wire   [6:0] \level_2_sums[16][61] ;
wire   [6:0] \level_2_sums[16][62] ;
wire   [6:0] \level_2_sums[16][63] ;
wire   [6:0] \level_2_sums[17][0] ;
wire   [6:0] \level_2_sums[17][1] ;
wire   [6:0] \level_2_sums[17][2] ;
wire   [6:0] \level_2_sums[17][3] ;
wire   [6:0] \level_2_sums[17][4] ;
wire   [6:0] \level_2_sums[17][5] ;
wire   [6:0] \level_2_sums[17][6] ;
wire   [6:0] \level_2_sums[17][7] ;
wire   [6:0] \level_2_sums[17][8] ;
wire   [6:0] \level_2_sums[17][9] ;
wire   [6:0] \level_2_sums[17][10] ;
wire   [6:0] \level_2_sums[17][11] ;
wire   [6:0] \level_2_sums[17][12] ;
wire   [6:0] \level_2_sums[17][13] ;
wire   [6:0] \level_2_sums[17][14] ;
wire   [6:0] \level_2_sums[17][15] ;
wire   [6:0] \level_2_sums[17][16] ;
wire   [6:0] \level_2_sums[17][17] ;
wire   [6:0] \level_2_sums[17][18] ;
wire   [6:0] \level_2_sums[17][19] ;
wire   [6:0] \level_2_sums[17][20] ;
wire   [6:0] \level_2_sums[17][21] ;
wire   [6:0] \level_2_sums[17][22] ;
wire   [6:0] \level_2_sums[17][23] ;
wire   [6:0] \level_2_sums[17][24] ;
wire   [6:0] \level_2_sums[17][25] ;
wire   [6:0] \level_2_sums[17][26] ;
wire   [6:0] \level_2_sums[17][27] ;
wire   [6:0] \level_2_sums[17][28] ;
wire   [6:0] \level_2_sums[17][29] ;
wire   [6:0] \level_2_sums[17][30] ;
wire   [6:0] \level_2_sums[17][31] ;
wire   [6:0] \level_2_sums[17][32] ;
wire   [6:0] \level_2_sums[17][33] ;
wire   [6:0] \level_2_sums[17][34] ;
wire   [6:0] \level_2_sums[17][35] ;
wire   [6:0] \level_2_sums[17][36] ;
wire   [6:0] \level_2_sums[17][37] ;
wire   [6:0] \level_2_sums[17][38] ;
wire   [6:0] \level_2_sums[17][39] ;
wire   [6:0] \level_2_sums[17][40] ;
wire   [6:0] \level_2_sums[17][41] ;
wire   [6:0] \level_2_sums[17][42] ;
wire   [6:0] \level_2_sums[17][43] ;
wire   [6:0] \level_2_sums[17][44] ;
wire   [6:0] \level_2_sums[17][45] ;
wire   [6:0] \level_2_sums[17][46] ;
wire   [6:0] \level_2_sums[17][47] ;
wire   [6:0] \level_2_sums[17][48] ;
wire   [6:0] \level_2_sums[17][49] ;
wire   [6:0] \level_2_sums[17][50] ;
wire   [6:0] \level_2_sums[17][51] ;
wire   [6:0] \level_2_sums[17][52] ;
wire   [6:0] \level_2_sums[17][53] ;
wire   [6:0] \level_2_sums[17][54] ;
wire   [6:0] \level_2_sums[17][55] ;
wire   [6:0] \level_2_sums[17][56] ;
wire   [6:0] \level_2_sums[17][57] ;
wire   [6:0] \level_2_sums[17][58] ;
wire   [6:0] \level_2_sums[17][59] ;
wire   [6:0] \level_2_sums[17][60] ;
wire   [6:0] \level_2_sums[17][61] ;
wire   [6:0] \level_2_sums[17][62] ;
wire   [6:0] \level_2_sums[17][63] ;
wire   [6:0] \level_2_sums[18][0] ;
wire   [6:0] \level_2_sums[18][1] ;
wire   [6:0] \level_2_sums[18][2] ;
wire   [6:0] \level_2_sums[18][3] ;
wire   [6:0] \level_2_sums[18][4] ;
wire   [6:0] \level_2_sums[18][5] ;
wire   [6:0] \level_2_sums[18][6] ;
wire   [6:0] \level_2_sums[18][7] ;
wire   [6:0] \level_2_sums[18][8] ;
wire   [6:0] \level_2_sums[18][9] ;
wire   [6:0] \level_2_sums[18][10] ;
wire   [6:0] \level_2_sums[18][11] ;
wire   [6:0] \level_2_sums[18][12] ;
wire   [6:0] \level_2_sums[18][13] ;
wire   [6:0] \level_2_sums[18][14] ;
wire   [6:0] \level_2_sums[18][15] ;
wire   [6:0] \level_2_sums[18][16] ;
wire   [6:0] \level_2_sums[18][17] ;
wire   [6:0] \level_2_sums[18][18] ;
wire   [6:0] \level_2_sums[18][19] ;
wire   [6:0] \level_2_sums[18][20] ;
wire   [6:0] \level_2_sums[18][21] ;
wire   [6:0] \level_2_sums[18][22] ;
wire   [6:0] \level_2_sums[18][23] ;
wire   [6:0] \level_2_sums[18][24] ;
wire   [6:0] \level_2_sums[18][25] ;
wire   [6:0] \level_2_sums[18][26] ;
wire   [6:0] \level_2_sums[18][27] ;
wire   [6:0] \level_2_sums[18][28] ;
wire   [6:0] \level_2_sums[18][29] ;
wire   [6:0] \level_2_sums[18][30] ;
wire   [6:0] \level_2_sums[18][31] ;
wire   [6:0] \level_2_sums[18][32] ;
wire   [6:0] \level_2_sums[18][33] ;
wire   [6:0] \level_2_sums[18][34] ;
wire   [6:0] \level_2_sums[18][35] ;
wire   [6:0] \level_2_sums[18][36] ;
wire   [6:0] \level_2_sums[18][37] ;
wire   [6:0] \level_2_sums[18][38] ;
wire   [6:0] \level_2_sums[18][39] ;
wire   [6:0] \level_2_sums[18][40] ;
wire   [6:0] \level_2_sums[18][41] ;
wire   [6:0] \level_2_sums[18][42] ;
wire   [6:0] \level_2_sums[18][43] ;
wire   [6:0] \level_2_sums[18][44] ;
wire   [6:0] \level_2_sums[18][45] ;
wire   [6:0] \level_2_sums[18][46] ;
wire   [6:0] \level_2_sums[18][47] ;
wire   [6:0] \level_2_sums[18][48] ;
wire   [6:0] \level_2_sums[18][49] ;
wire   [6:0] \level_2_sums[18][50] ;
wire   [6:0] \level_2_sums[18][51] ;
wire   [6:0] \level_2_sums[18][52] ;
wire   [6:0] \level_2_sums[18][53] ;
wire   [6:0] \level_2_sums[18][54] ;
wire   [6:0] \level_2_sums[18][55] ;
wire   [6:0] \level_2_sums[18][56] ;
wire   [6:0] \level_2_sums[18][57] ;
wire   [6:0] \level_2_sums[18][58] ;
wire   [6:0] \level_2_sums[18][59] ;
wire   [6:0] \level_2_sums[18][60] ;
wire   [6:0] \level_2_sums[18][61] ;
wire   [6:0] \level_2_sums[18][62] ;
wire   [6:0] \level_2_sums[18][63] ;
wire   [6:0] \level_2_sums[19][0] ;
wire   [6:0] \level_2_sums[19][1] ;
wire   [6:0] \level_2_sums[19][2] ;
wire   [6:0] \level_2_sums[19][3] ;
wire   [6:0] \level_2_sums[19][4] ;
wire   [6:0] \level_2_sums[19][5] ;
wire   [6:0] \level_2_sums[19][6] ;
wire   [6:0] \level_2_sums[19][7] ;
wire   [6:0] \level_2_sums[19][8] ;
wire   [6:0] \level_2_sums[19][9] ;
wire   [6:0] \level_2_sums[19][10] ;
wire   [6:0] \level_2_sums[19][11] ;
wire   [6:0] \level_2_sums[19][12] ;
wire   [6:0] \level_2_sums[19][13] ;
wire   [6:0] \level_2_sums[19][14] ;
wire   [6:0] \level_2_sums[19][15] ;
wire   [6:0] \level_2_sums[19][16] ;
wire   [6:0] \level_2_sums[19][17] ;
wire   [6:0] \level_2_sums[19][18] ;
wire   [6:0] \level_2_sums[19][19] ;
wire   [6:0] \level_2_sums[19][20] ;
wire   [6:0] \level_2_sums[19][21] ;
wire   [6:0] \level_2_sums[19][22] ;
wire   [6:0] \level_2_sums[19][23] ;
wire   [6:0] \level_2_sums[19][24] ;
wire   [6:0] \level_2_sums[19][25] ;
wire   [6:0] \level_2_sums[19][26] ;
wire   [6:0] \level_2_sums[19][27] ;
wire   [6:0] \level_2_sums[19][28] ;
wire   [6:0] \level_2_sums[19][29] ;
wire   [6:0] \level_2_sums[19][30] ;
wire   [6:0] \level_2_sums[19][31] ;
wire   [6:0] \level_2_sums[19][32] ;
wire   [6:0] \level_2_sums[19][33] ;
wire   [6:0] \level_2_sums[19][34] ;
wire   [6:0] \level_2_sums[19][35] ;
wire   [6:0] \level_2_sums[19][36] ;
wire   [6:0] \level_2_sums[19][37] ;
wire   [6:0] \level_2_sums[19][38] ;
wire   [6:0] \level_2_sums[19][39] ;
wire   [6:0] \level_2_sums[19][40] ;
wire   [6:0] \level_2_sums[19][41] ;
wire   [6:0] \level_2_sums[19][42] ;
wire   [6:0] \level_2_sums[19][43] ;
wire   [6:0] \level_2_sums[19][44] ;
wire   [6:0] \level_2_sums[19][45] ;
wire   [6:0] \level_2_sums[19][46] ;
wire   [6:0] \level_2_sums[19][47] ;
wire   [6:0] \level_2_sums[19][48] ;
wire   [6:0] \level_2_sums[19][49] ;
wire   [6:0] \level_2_sums[19][50] ;
wire   [6:0] \level_2_sums[19][51] ;
wire   [6:0] \level_2_sums[19][52] ;
wire   [6:0] \level_2_sums[19][53] ;
wire   [6:0] \level_2_sums[19][54] ;
wire   [6:0] \level_2_sums[19][55] ;
wire   [6:0] \level_2_sums[19][56] ;
wire   [6:0] \level_2_sums[19][57] ;
wire   [6:0] \level_2_sums[19][58] ;
wire   [6:0] \level_2_sums[19][59] ;
wire   [6:0] \level_2_sums[19][60] ;
wire   [6:0] \level_2_sums[19][61] ;
wire   [6:0] \level_2_sums[19][62] ;
wire   [6:0] \level_2_sums[19][63] ;
wire   [5:0] \level_1_sums[0][0] ;
wire   [5:0] \level_1_sums[0][1] ;
wire   [5:0] \level_1_sums[0][2] ;
wire   [5:0] \level_1_sums[0][3] ;
wire   [5:0] \level_1_sums[0][4] ;
wire   [5:0] \level_1_sums[0][5] ;
wire   [5:0] \level_1_sums[0][6] ;
wire   [5:0] \level_1_sums[0][7] ;
wire   [5:0] \level_1_sums[0][8] ;
wire   [5:0] \level_1_sums[0][9] ;
wire   [5:0] \level_1_sums[0][10] ;
wire   [5:0] \level_1_sums[0][11] ;
wire   [5:0] \level_1_sums[0][12] ;
wire   [5:0] \level_1_sums[0][13] ;
wire   [5:0] \level_1_sums[0][14] ;
wire   [5:0] \level_1_sums[0][15] ;
wire   [5:0] \level_1_sums[0][16] ;
wire   [5:0] \level_1_sums[0][17] ;
wire   [5:0] \level_1_sums[0][18] ;
wire   [5:0] \level_1_sums[0][19] ;
wire   [5:0] \level_1_sums[0][20] ;
wire   [5:0] \level_1_sums[0][21] ;
wire   [5:0] \level_1_sums[0][22] ;
wire   [5:0] \level_1_sums[0][23] ;
wire   [5:0] \level_1_sums[0][24] ;
wire   [5:0] \level_1_sums[0][25] ;
wire   [5:0] \level_1_sums[0][26] ;
wire   [5:0] \level_1_sums[0][27] ;
wire   [5:0] \level_1_sums[0][28] ;
wire   [5:0] \level_1_sums[0][29] ;
wire   [5:0] \level_1_sums[0][30] ;
wire   [5:0] \level_1_sums[0][31] ;
wire   [5:0] \level_1_sums[0][32] ;
wire   [5:0] \level_1_sums[0][33] ;
wire   [5:0] \level_1_sums[0][34] ;
wire   [5:0] \level_1_sums[0][35] ;
wire   [5:0] \level_1_sums[0][36] ;
wire   [5:0] \level_1_sums[0][37] ;
wire   [5:0] \level_1_sums[0][38] ;
wire   [5:0] \level_1_sums[0][39] ;
wire   [5:0] \level_1_sums[0][40] ;
wire   [5:0] \level_1_sums[0][41] ;
wire   [5:0] \level_1_sums[0][42] ;
wire   [5:0] \level_1_sums[0][43] ;
wire   [5:0] \level_1_sums[0][44] ;
wire   [5:0] \level_1_sums[0][45] ;
wire   [5:0] \level_1_sums[0][46] ;
wire   [5:0] \level_1_sums[0][47] ;
wire   [5:0] \level_1_sums[0][48] ;
wire   [5:0] \level_1_sums[0][49] ;
wire   [5:0] \level_1_sums[0][50] ;
wire   [5:0] \level_1_sums[0][51] ;
wire   [5:0] \level_1_sums[0][52] ;
wire   [5:0] \level_1_sums[0][53] ;
wire   [5:0] \level_1_sums[0][54] ;
wire   [5:0] \level_1_sums[0][55] ;
wire   [5:0] \level_1_sums[0][56] ;
wire   [5:0] \level_1_sums[0][57] ;
wire   [5:0] \level_1_sums[0][58] ;
wire   [5:0] \level_1_sums[0][59] ;
wire   [5:0] \level_1_sums[0][60] ;
wire   [5:0] \level_1_sums[0][61] ;
wire   [5:0] \level_1_sums[0][62] ;
wire   [5:0] \level_1_sums[0][63] ;
wire   [5:0] \level_1_sums[0][64] ;
wire   [5:0] \level_1_sums[0][65] ;
wire   [5:0] \level_1_sums[0][66] ;
wire   [5:0] \level_1_sums[0][67] ;
wire   [5:0] \level_1_sums[0][68] ;
wire   [5:0] \level_1_sums[0][69] ;
wire   [5:0] \level_1_sums[0][70] ;
wire   [5:0] \level_1_sums[0][71] ;
wire   [5:0] \level_1_sums[0][72] ;
wire   [5:0] \level_1_sums[0][73] ;
wire   [5:0] \level_1_sums[0][74] ;
wire   [5:0] \level_1_sums[0][75] ;
wire   [5:0] \level_1_sums[0][76] ;
wire   [5:0] \level_1_sums[0][77] ;
wire   [5:0] \level_1_sums[0][78] ;
wire   [5:0] \level_1_sums[0][79] ;
wire   [5:0] \level_1_sums[0][80] ;
wire   [5:0] \level_1_sums[0][81] ;
wire   [5:0] \level_1_sums[0][82] ;
wire   [5:0] \level_1_sums[0][83] ;
wire   [5:0] \level_1_sums[0][84] ;
wire   [5:0] \level_1_sums[0][85] ;
wire   [5:0] \level_1_sums[0][86] ;
wire   [5:0] \level_1_sums[0][87] ;
wire   [5:0] \level_1_sums[0][88] ;
wire   [5:0] \level_1_sums[0][89] ;
wire   [5:0] \level_1_sums[0][90] ;
wire   [5:0] \level_1_sums[0][91] ;
wire   [5:0] \level_1_sums[0][92] ;
wire   [5:0] \level_1_sums[0][93] ;
wire   [5:0] \level_1_sums[0][94] ;
wire   [5:0] \level_1_sums[0][95] ;
wire   [5:0] \level_1_sums[0][96] ;
wire   [5:0] \level_1_sums[0][97] ;
wire   [5:0] \level_1_sums[0][98] ;
wire   [5:0] \level_1_sums[0][99] ;
wire   [5:0] \level_1_sums[0][100] ;
wire   [5:0] \level_1_sums[0][101] ;
wire   [5:0] \level_1_sums[0][102] ;
wire   [5:0] \level_1_sums[0][103] ;
wire   [5:0] \level_1_sums[0][104] ;
wire   [5:0] \level_1_sums[0][105] ;
wire   [5:0] \level_1_sums[0][106] ;
wire   [5:0] \level_1_sums[0][107] ;
wire   [5:0] \level_1_sums[0][108] ;
wire   [5:0] \level_1_sums[0][109] ;
wire   [5:0] \level_1_sums[0][110] ;
wire   [5:0] \level_1_sums[0][111] ;
wire   [5:0] \level_1_sums[0][112] ;
wire   [5:0] \level_1_sums[0][113] ;
wire   [5:0] \level_1_sums[0][114] ;
wire   [5:0] \level_1_sums[0][115] ;
wire   [5:0] \level_1_sums[0][116] ;
wire   [5:0] \level_1_sums[0][117] ;
wire   [5:0] \level_1_sums[0][118] ;
wire   [5:0] \level_1_sums[0][119] ;
wire   [5:0] \level_1_sums[0][120] ;
wire   [5:0] \level_1_sums[0][121] ;
wire   [5:0] \level_1_sums[0][122] ;
wire   [5:0] \level_1_sums[0][123] ;
wire   [5:0] \level_1_sums[0][124] ;
wire   [5:0] \level_1_sums[0][125] ;
wire   [5:0] \level_1_sums[0][126] ;
wire   [5:0] \level_1_sums[0][127] ;
wire   [5:0] \level_1_sums[1][0] ;
wire   [5:0] \level_1_sums[1][1] ;
wire   [5:0] \level_1_sums[1][2] ;
wire   [5:0] \level_1_sums[1][3] ;
wire   [5:0] \level_1_sums[1][4] ;
wire   [5:0] \level_1_sums[1][5] ;
wire   [5:0] \level_1_sums[1][6] ;
wire   [5:0] \level_1_sums[1][7] ;
wire   [5:0] \level_1_sums[1][8] ;
wire   [5:0] \level_1_sums[1][9] ;
wire   [5:0] \level_1_sums[1][10] ;
wire   [5:0] \level_1_sums[1][11] ;
wire   [5:0] \level_1_sums[1][12] ;
wire   [5:0] \level_1_sums[1][13] ;
wire   [5:0] \level_1_sums[1][14] ;
wire   [5:0] \level_1_sums[1][15] ;
wire   [5:0] \level_1_sums[1][16] ;
wire   [5:0] \level_1_sums[1][17] ;
wire   [5:0] \level_1_sums[1][18] ;
wire   [5:0] \level_1_sums[1][19] ;
wire   [5:0] \level_1_sums[1][20] ;
wire   [5:0] \level_1_sums[1][21] ;
wire   [5:0] \level_1_sums[1][22] ;
wire   [5:0] \level_1_sums[1][23] ;
wire   [5:0] \level_1_sums[1][24] ;
wire   [5:0] \level_1_sums[1][25] ;
wire   [5:0] \level_1_sums[1][26] ;
wire   [5:0] \level_1_sums[1][27] ;
wire   [5:0] \level_1_sums[1][28] ;
wire   [5:0] \level_1_sums[1][29] ;
wire   [5:0] \level_1_sums[1][30] ;
wire   [5:0] \level_1_sums[1][31] ;
wire   [5:0] \level_1_sums[1][32] ;
wire   [5:0] \level_1_sums[1][33] ;
wire   [5:0] \level_1_sums[1][34] ;
wire   [5:0] \level_1_sums[1][35] ;
wire   [5:0] \level_1_sums[1][36] ;
wire   [5:0] \level_1_sums[1][37] ;
wire   [5:0] \level_1_sums[1][38] ;
wire   [5:0] \level_1_sums[1][39] ;
wire   [5:0] \level_1_sums[1][40] ;
wire   [5:0] \level_1_sums[1][41] ;
wire   [5:0] \level_1_sums[1][42] ;
wire   [5:0] \level_1_sums[1][43] ;
wire   [5:0] \level_1_sums[1][44] ;
wire   [5:0] \level_1_sums[1][45] ;
wire   [5:0] \level_1_sums[1][46] ;
wire   [5:0] \level_1_sums[1][47] ;
wire   [5:0] \level_1_sums[1][48] ;
wire   [5:0] \level_1_sums[1][49] ;
wire   [5:0] \level_1_sums[1][50] ;
wire   [5:0] \level_1_sums[1][51] ;
wire   [5:0] \level_1_sums[1][52] ;
wire   [5:0] \level_1_sums[1][53] ;
wire   [5:0] \level_1_sums[1][54] ;
wire   [5:0] \level_1_sums[1][55] ;
wire   [5:0] \level_1_sums[1][56] ;
wire   [5:0] \level_1_sums[1][57] ;
wire   [5:0] \level_1_sums[1][58] ;
wire   [5:0] \level_1_sums[1][59] ;
wire   [5:0] \level_1_sums[1][60] ;
wire   [5:0] \level_1_sums[1][61] ;
wire   [5:0] \level_1_sums[1][62] ;
wire   [5:0] \level_1_sums[1][63] ;
wire   [5:0] \level_1_sums[1][64] ;
wire   [5:0] \level_1_sums[1][65] ;
wire   [5:0] \level_1_sums[1][66] ;
wire   [5:0] \level_1_sums[1][67] ;
wire   [5:0] \level_1_sums[1][68] ;
wire   [5:0] \level_1_sums[1][69] ;
wire   [5:0] \level_1_sums[1][70] ;
wire   [5:0] \level_1_sums[1][71] ;
wire   [5:0] \level_1_sums[1][72] ;
wire   [5:0] \level_1_sums[1][73] ;
wire   [5:0] \level_1_sums[1][74] ;
wire   [5:0] \level_1_sums[1][75] ;
wire   [5:0] \level_1_sums[1][76] ;
wire   [5:0] \level_1_sums[1][77] ;
wire   [5:0] \level_1_sums[1][78] ;
wire   [5:0] \level_1_sums[1][79] ;
wire   [5:0] \level_1_sums[1][80] ;
wire   [5:0] \level_1_sums[1][81] ;
wire   [5:0] \level_1_sums[1][82] ;
wire   [5:0] \level_1_sums[1][83] ;
wire   [5:0] \level_1_sums[1][84] ;
wire   [5:0] \level_1_sums[1][85] ;
wire   [5:0] \level_1_sums[1][86] ;
wire   [5:0] \level_1_sums[1][87] ;
wire   [5:0] \level_1_sums[1][88] ;
wire   [5:0] \level_1_sums[1][89] ;
wire   [5:0] \level_1_sums[1][90] ;
wire   [5:0] \level_1_sums[1][91] ;
wire   [5:0] \level_1_sums[1][92] ;
wire   [5:0] \level_1_sums[1][93] ;
wire   [5:0] \level_1_sums[1][94] ;
wire   [5:0] \level_1_sums[1][95] ;
wire   [5:0] \level_1_sums[1][96] ;
wire   [5:0] \level_1_sums[1][97] ;
wire   [5:0] \level_1_sums[1][98] ;
wire   [5:0] \level_1_sums[1][99] ;
wire   [5:0] \level_1_sums[1][100] ;
wire   [5:0] \level_1_sums[1][101] ;
wire   [5:0] \level_1_sums[1][102] ;
wire   [5:0] \level_1_sums[1][103] ;
wire   [5:0] \level_1_sums[1][104] ;
wire   [5:0] \level_1_sums[1][105] ;
wire   [5:0] \level_1_sums[1][106] ;
wire   [5:0] \level_1_sums[1][107] ;
wire   [5:0] \level_1_sums[1][108] ;
wire   [5:0] \level_1_sums[1][109] ;
wire   [5:0] \level_1_sums[1][110] ;
wire   [5:0] \level_1_sums[1][111] ;
wire   [5:0] \level_1_sums[1][112] ;
wire   [5:0] \level_1_sums[1][113] ;
wire   [5:0] \level_1_sums[1][114] ;
wire   [5:0] \level_1_sums[1][115] ;
wire   [5:0] \level_1_sums[1][116] ;
wire   [5:0] \level_1_sums[1][117] ;
wire   [5:0] \level_1_sums[1][118] ;
wire   [5:0] \level_1_sums[1][119] ;
wire   [5:0] \level_1_sums[1][120] ;
wire   [5:0] \level_1_sums[1][121] ;
wire   [5:0] \level_1_sums[1][122] ;
wire   [5:0] \level_1_sums[1][123] ;
wire   [5:0] \level_1_sums[1][124] ;
wire   [5:0] \level_1_sums[1][125] ;
wire   [5:0] \level_1_sums[1][126] ;
wire   [5:0] \level_1_sums[1][127] ;
wire   [5:0] \level_1_sums[2][0] ;
wire   [5:0] \level_1_sums[2][1] ;
wire   [5:0] \level_1_sums[2][2] ;
wire   [5:0] \level_1_sums[2][3] ;
wire   [5:0] \level_1_sums[2][4] ;
wire   [5:0] \level_1_sums[2][5] ;
wire   [5:0] \level_1_sums[2][6] ;
wire   [5:0] \level_1_sums[2][7] ;
wire   [5:0] \level_1_sums[2][8] ;
wire   [5:0] \level_1_sums[2][9] ;
wire   [5:0] \level_1_sums[2][10] ;
wire   [5:0] \level_1_sums[2][11] ;
wire   [5:0] \level_1_sums[2][12] ;
wire   [5:0] \level_1_sums[2][13] ;
wire   [5:0] \level_1_sums[2][14] ;
wire   [5:0] \level_1_sums[2][15] ;
wire   [5:0] \level_1_sums[2][16] ;
wire   [5:0] \level_1_sums[2][17] ;
wire   [5:0] \level_1_sums[2][18] ;
wire   [5:0] \level_1_sums[2][19] ;
wire   [5:0] \level_1_sums[2][20] ;
wire   [5:0] \level_1_sums[2][21] ;
wire   [5:0] \level_1_sums[2][22] ;
wire   [5:0] \level_1_sums[2][23] ;
wire   [5:0] \level_1_sums[2][24] ;
wire   [5:0] \level_1_sums[2][25] ;
wire   [5:0] \level_1_sums[2][26] ;
wire   [5:0] \level_1_sums[2][27] ;
wire   [5:0] \level_1_sums[2][28] ;
wire   [5:0] \level_1_sums[2][29] ;
wire   [5:0] \level_1_sums[2][30] ;
wire   [5:0] \level_1_sums[2][31] ;
wire   [5:0] \level_1_sums[2][32] ;
wire   [5:0] \level_1_sums[2][33] ;
wire   [5:0] \level_1_sums[2][34] ;
wire   [5:0] \level_1_sums[2][35] ;
wire   [5:0] \level_1_sums[2][36] ;
wire   [5:0] \level_1_sums[2][37] ;
wire   [5:0] \level_1_sums[2][38] ;
wire   [5:0] \level_1_sums[2][39] ;
wire   [5:0] \level_1_sums[2][40] ;
wire   [5:0] \level_1_sums[2][41] ;
wire   [5:0] \level_1_sums[2][42] ;
wire   [5:0] \level_1_sums[2][43] ;
wire   [5:0] \level_1_sums[2][44] ;
wire   [5:0] \level_1_sums[2][45] ;
wire   [5:0] \level_1_sums[2][46] ;
wire   [5:0] \level_1_sums[2][47] ;
wire   [5:0] \level_1_sums[2][48] ;
wire   [5:0] \level_1_sums[2][49] ;
wire   [5:0] \level_1_sums[2][50] ;
wire   [5:0] \level_1_sums[2][51] ;
wire   [5:0] \level_1_sums[2][52] ;
wire   [5:0] \level_1_sums[2][53] ;
wire   [5:0] \level_1_sums[2][54] ;
wire   [5:0] \level_1_sums[2][55] ;
wire   [5:0] \level_1_sums[2][56] ;
wire   [5:0] \level_1_sums[2][57] ;
wire   [5:0] \level_1_sums[2][58] ;
wire   [5:0] \level_1_sums[2][59] ;
wire   [5:0] \level_1_sums[2][60] ;
wire   [5:0] \level_1_sums[2][61] ;
wire   [5:0] \level_1_sums[2][62] ;
wire   [5:0] \level_1_sums[2][63] ;
wire   [5:0] \level_1_sums[2][64] ;
wire   [5:0] \level_1_sums[2][65] ;
wire   [5:0] \level_1_sums[2][66] ;
wire   [5:0] \level_1_sums[2][67] ;
wire   [5:0] \level_1_sums[2][68] ;
wire   [5:0] \level_1_sums[2][69] ;
wire   [5:0] \level_1_sums[2][70] ;
wire   [5:0] \level_1_sums[2][71] ;
wire   [5:0] \level_1_sums[2][72] ;
wire   [5:0] \level_1_sums[2][73] ;
wire   [5:0] \level_1_sums[2][74] ;
wire   [5:0] \level_1_sums[2][75] ;
wire   [5:0] \level_1_sums[2][76] ;
wire   [5:0] \level_1_sums[2][77] ;
wire   [5:0] \level_1_sums[2][78] ;
wire   [5:0] \level_1_sums[2][79] ;
wire   [5:0] \level_1_sums[2][80] ;
wire   [5:0] \level_1_sums[2][81] ;
wire   [5:0] \level_1_sums[2][82] ;
wire   [5:0] \level_1_sums[2][83] ;
wire   [5:0] \level_1_sums[2][84] ;
wire   [5:0] \level_1_sums[2][85] ;
wire   [5:0] \level_1_sums[2][86] ;
wire   [5:0] \level_1_sums[2][87] ;
wire   [5:0] \level_1_sums[2][88] ;
wire   [5:0] \level_1_sums[2][89] ;
wire   [5:0] \level_1_sums[2][90] ;
wire   [5:0] \level_1_sums[2][91] ;
wire   [5:0] \level_1_sums[2][92] ;
wire   [5:0] \level_1_sums[2][93] ;
wire   [5:0] \level_1_sums[2][94] ;
wire   [5:0] \level_1_sums[2][95] ;
wire   [5:0] \level_1_sums[2][96] ;
wire   [5:0] \level_1_sums[2][97] ;
wire   [5:0] \level_1_sums[2][98] ;
wire   [5:0] \level_1_sums[2][99] ;
wire   [5:0] \level_1_sums[2][100] ;
wire   [5:0] \level_1_sums[2][101] ;
wire   [5:0] \level_1_sums[2][102] ;
wire   [5:0] \level_1_sums[2][103] ;
wire   [5:0] \level_1_sums[2][104] ;
wire   [5:0] \level_1_sums[2][105] ;
wire   [5:0] \level_1_sums[2][106] ;
wire   [5:0] \level_1_sums[2][107] ;
wire   [5:0] \level_1_sums[2][108] ;
wire   [5:0] \level_1_sums[2][109] ;
wire   [5:0] \level_1_sums[2][110] ;
wire   [5:0] \level_1_sums[2][111] ;
wire   [5:0] \level_1_sums[2][112] ;
wire   [5:0] \level_1_sums[2][113] ;
wire   [5:0] \level_1_sums[2][114] ;
wire   [5:0] \level_1_sums[2][115] ;
wire   [5:0] \level_1_sums[2][116] ;
wire   [5:0] \level_1_sums[2][117] ;
wire   [5:0] \level_1_sums[2][118] ;
wire   [5:0] \level_1_sums[2][119] ;
wire   [5:0] \level_1_sums[2][120] ;
wire   [5:0] \level_1_sums[2][121] ;
wire   [5:0] \level_1_sums[2][122] ;
wire   [5:0] \level_1_sums[2][123] ;
wire   [5:0] \level_1_sums[2][124] ;
wire   [5:0] \level_1_sums[2][125] ;
wire   [5:0] \level_1_sums[2][126] ;
wire   [5:0] \level_1_sums[2][127] ;
wire   [5:0] \level_1_sums[3][0] ;
wire   [5:0] \level_1_sums[3][1] ;
wire   [5:0] \level_1_sums[3][2] ;
wire   [5:0] \level_1_sums[3][3] ;
wire   [5:0] \level_1_sums[3][4] ;
wire   [5:0] \level_1_sums[3][5] ;
wire   [5:0] \level_1_sums[3][6] ;
wire   [5:0] \level_1_sums[3][7] ;
wire   [5:0] \level_1_sums[3][8] ;
wire   [5:0] \level_1_sums[3][9] ;
wire   [5:0] \level_1_sums[3][10] ;
wire   [5:0] \level_1_sums[3][11] ;
wire   [5:0] \level_1_sums[3][12] ;
wire   [5:0] \level_1_sums[3][13] ;
wire   [5:0] \level_1_sums[3][14] ;
wire   [5:0] \level_1_sums[3][15] ;
wire   [5:0] \level_1_sums[3][16] ;
wire   [5:0] \level_1_sums[3][17] ;
wire   [5:0] \level_1_sums[3][18] ;
wire   [5:0] \level_1_sums[3][19] ;
wire   [5:0] \level_1_sums[3][20] ;
wire   [5:0] \level_1_sums[3][21] ;
wire   [5:0] \level_1_sums[3][22] ;
wire   [5:0] \level_1_sums[3][23] ;
wire   [5:0] \level_1_sums[3][24] ;
wire   [5:0] \level_1_sums[3][25] ;
wire   [5:0] \level_1_sums[3][26] ;
wire   [5:0] \level_1_sums[3][27] ;
wire   [5:0] \level_1_sums[3][28] ;
wire   [5:0] \level_1_sums[3][29] ;
wire   [5:0] \level_1_sums[3][30] ;
wire   [5:0] \level_1_sums[3][31] ;
wire   [5:0] \level_1_sums[3][32] ;
wire   [5:0] \level_1_sums[3][33] ;
wire   [5:0] \level_1_sums[3][34] ;
wire   [5:0] \level_1_sums[3][35] ;
wire   [5:0] \level_1_sums[3][36] ;
wire   [5:0] \level_1_sums[3][37] ;
wire   [5:0] \level_1_sums[3][38] ;
wire   [5:0] \level_1_sums[3][39] ;
wire   [5:0] \level_1_sums[3][40] ;
wire   [5:0] \level_1_sums[3][41] ;
wire   [5:0] \level_1_sums[3][42] ;
wire   [5:0] \level_1_sums[3][43] ;
wire   [5:0] \level_1_sums[3][44] ;
wire   [5:0] \level_1_sums[3][45] ;
wire   [5:0] \level_1_sums[3][46] ;
wire   [5:0] \level_1_sums[3][47] ;
wire   [5:0] \level_1_sums[3][48] ;
wire   [5:0] \level_1_sums[3][49] ;
wire   [5:0] \level_1_sums[3][50] ;
wire   [5:0] \level_1_sums[3][51] ;
wire   [5:0] \level_1_sums[3][52] ;
wire   [5:0] \level_1_sums[3][53] ;
wire   [5:0] \level_1_sums[3][54] ;
wire   [5:0] \level_1_sums[3][55] ;
wire   [5:0] \level_1_sums[3][56] ;
wire   [5:0] \level_1_sums[3][57] ;
wire   [5:0] \level_1_sums[3][58] ;
wire   [5:0] \level_1_sums[3][59] ;
wire   [5:0] \level_1_sums[3][60] ;
wire   [5:0] \level_1_sums[3][61] ;
wire   [5:0] \level_1_sums[3][62] ;
wire   [5:0] \level_1_sums[3][63] ;
wire   [5:0] \level_1_sums[3][64] ;
wire   [5:0] \level_1_sums[3][65] ;
wire   [5:0] \level_1_sums[3][66] ;
wire   [5:0] \level_1_sums[3][67] ;
wire   [5:0] \level_1_sums[3][68] ;
wire   [5:0] \level_1_sums[3][69] ;
wire   [5:0] \level_1_sums[3][70] ;
wire   [5:0] \level_1_sums[3][71] ;
wire   [5:0] \level_1_sums[3][72] ;
wire   [5:0] \level_1_sums[3][73] ;
wire   [5:0] \level_1_sums[3][74] ;
wire   [5:0] \level_1_sums[3][75] ;
wire   [5:0] \level_1_sums[3][76] ;
wire   [5:0] \level_1_sums[3][77] ;
wire   [5:0] \level_1_sums[3][78] ;
wire   [5:0] \level_1_sums[3][79] ;
wire   [5:0] \level_1_sums[3][80] ;
wire   [5:0] \level_1_sums[3][81] ;
wire   [5:0] \level_1_sums[3][82] ;
wire   [5:0] \level_1_sums[3][83] ;
wire   [5:0] \level_1_sums[3][84] ;
wire   [5:0] \level_1_sums[3][85] ;
wire   [5:0] \level_1_sums[3][86] ;
wire   [5:0] \level_1_sums[3][87] ;
wire   [5:0] \level_1_sums[3][88] ;
wire   [5:0] \level_1_sums[3][89] ;
wire   [5:0] \level_1_sums[3][90] ;
wire   [5:0] \level_1_sums[3][91] ;
wire   [5:0] \level_1_sums[3][92] ;
wire   [5:0] \level_1_sums[3][93] ;
wire   [5:0] \level_1_sums[3][94] ;
wire   [5:0] \level_1_sums[3][95] ;
wire   [5:0] \level_1_sums[3][96] ;
wire   [5:0] \level_1_sums[3][97] ;
wire   [5:0] \level_1_sums[3][98] ;
wire   [5:0] \level_1_sums[3][99] ;
wire   [5:0] \level_1_sums[3][100] ;
wire   [5:0] \level_1_sums[3][101] ;
wire   [5:0] \level_1_sums[3][102] ;
wire   [5:0] \level_1_sums[3][103] ;
wire   [5:0] \level_1_sums[3][104] ;
wire   [5:0] \level_1_sums[3][105] ;
wire   [5:0] \level_1_sums[3][106] ;
wire   [5:0] \level_1_sums[3][107] ;
wire   [5:0] \level_1_sums[3][108] ;
wire   [5:0] \level_1_sums[3][109] ;
wire   [5:0] \level_1_sums[3][110] ;
wire   [5:0] \level_1_sums[3][111] ;
wire   [5:0] \level_1_sums[3][112] ;
wire   [5:0] \level_1_sums[3][113] ;
wire   [5:0] \level_1_sums[3][114] ;
wire   [5:0] \level_1_sums[3][115] ;
wire   [5:0] \level_1_sums[3][116] ;
wire   [5:0] \level_1_sums[3][117] ;
wire   [5:0] \level_1_sums[3][118] ;
wire   [5:0] \level_1_sums[3][119] ;
wire   [5:0] \level_1_sums[3][120] ;
wire   [5:0] \level_1_sums[3][121] ;
wire   [5:0] \level_1_sums[3][122] ;
wire   [5:0] \level_1_sums[3][123] ;
wire   [5:0] \level_1_sums[3][124] ;
wire   [5:0] \level_1_sums[3][125] ;
wire   [5:0] \level_1_sums[3][126] ;
wire   [5:0] \level_1_sums[3][127] ;
wire   [5:0] \level_1_sums[4][0] ;
wire   [5:0] \level_1_sums[4][1] ;
wire   [5:0] \level_1_sums[4][2] ;
wire   [5:0] \level_1_sums[4][3] ;
wire   [5:0] \level_1_sums[4][4] ;
wire   [5:0] \level_1_sums[4][5] ;
wire   [5:0] \level_1_sums[4][6] ;
wire   [5:0] \level_1_sums[4][7] ;
wire   [5:0] \level_1_sums[4][8] ;
wire   [5:0] \level_1_sums[4][9] ;
wire   [5:0] \level_1_sums[4][10] ;
wire   [5:0] \level_1_sums[4][11] ;
wire   [5:0] \level_1_sums[4][12] ;
wire   [5:0] \level_1_sums[4][13] ;
wire   [5:0] \level_1_sums[4][14] ;
wire   [5:0] \level_1_sums[4][15] ;
wire   [5:0] \level_1_sums[4][16] ;
wire   [5:0] \level_1_sums[4][17] ;
wire   [5:0] \level_1_sums[4][18] ;
wire   [5:0] \level_1_sums[4][19] ;
wire   [5:0] \level_1_sums[4][20] ;
wire   [5:0] \level_1_sums[4][21] ;
wire   [5:0] \level_1_sums[4][22] ;
wire   [5:0] \level_1_sums[4][23] ;
wire   [5:0] \level_1_sums[4][24] ;
wire   [5:0] \level_1_sums[4][25] ;
wire   [5:0] \level_1_sums[4][26] ;
wire   [5:0] \level_1_sums[4][27] ;
wire   [5:0] \level_1_sums[4][28] ;
wire   [5:0] \level_1_sums[4][29] ;
wire   [5:0] \level_1_sums[4][30] ;
wire   [5:0] \level_1_sums[4][31] ;
wire   [5:0] \level_1_sums[4][32] ;
wire   [5:0] \level_1_sums[4][33] ;
wire   [5:0] \level_1_sums[4][34] ;
wire   [5:0] \level_1_sums[4][35] ;
wire   [5:0] \level_1_sums[4][36] ;
wire   [5:0] \level_1_sums[4][37] ;
wire   [5:0] \level_1_sums[4][38] ;
wire   [5:0] \level_1_sums[4][39] ;
wire   [5:0] \level_1_sums[4][40] ;
wire   [5:0] \level_1_sums[4][41] ;
wire   [5:0] \level_1_sums[4][42] ;
wire   [5:0] \level_1_sums[4][43] ;
wire   [5:0] \level_1_sums[4][44] ;
wire   [5:0] \level_1_sums[4][45] ;
wire   [5:0] \level_1_sums[4][46] ;
wire   [5:0] \level_1_sums[4][47] ;
wire   [5:0] \level_1_sums[4][48] ;
wire   [5:0] \level_1_sums[4][49] ;
wire   [5:0] \level_1_sums[4][50] ;
wire   [5:0] \level_1_sums[4][51] ;
wire   [5:0] \level_1_sums[4][52] ;
wire   [5:0] \level_1_sums[4][53] ;
wire   [5:0] \level_1_sums[4][54] ;
wire   [5:0] \level_1_sums[4][55] ;
wire   [5:0] \level_1_sums[4][56] ;
wire   [5:0] \level_1_sums[4][57] ;
wire   [5:0] \level_1_sums[4][58] ;
wire   [5:0] \level_1_sums[4][59] ;
wire   [5:0] \level_1_sums[4][60] ;
wire   [5:0] \level_1_sums[4][61] ;
wire   [5:0] \level_1_sums[4][62] ;
wire   [5:0] \level_1_sums[4][63] ;
wire   [5:0] \level_1_sums[4][64] ;
wire   [5:0] \level_1_sums[4][65] ;
wire   [5:0] \level_1_sums[4][66] ;
wire   [5:0] \level_1_sums[4][67] ;
wire   [5:0] \level_1_sums[4][68] ;
wire   [5:0] \level_1_sums[4][69] ;
wire   [5:0] \level_1_sums[4][70] ;
wire   [5:0] \level_1_sums[4][71] ;
wire   [5:0] \level_1_sums[4][72] ;
wire   [5:0] \level_1_sums[4][73] ;
wire   [5:0] \level_1_sums[4][74] ;
wire   [5:0] \level_1_sums[4][75] ;
wire   [5:0] \level_1_sums[4][76] ;
wire   [5:0] \level_1_sums[4][77] ;
wire   [5:0] \level_1_sums[4][78] ;
wire   [5:0] \level_1_sums[4][79] ;
wire   [5:0] \level_1_sums[4][80] ;
wire   [5:0] \level_1_sums[4][81] ;
wire   [5:0] \level_1_sums[4][82] ;
wire   [5:0] \level_1_sums[4][83] ;
wire   [5:0] \level_1_sums[4][84] ;
wire   [5:0] \level_1_sums[4][85] ;
wire   [5:0] \level_1_sums[4][86] ;
wire   [5:0] \level_1_sums[4][87] ;
wire   [5:0] \level_1_sums[4][88] ;
wire   [5:0] \level_1_sums[4][89] ;
wire   [5:0] \level_1_sums[4][90] ;
wire   [5:0] \level_1_sums[4][91] ;
wire   [5:0] \level_1_sums[4][92] ;
wire   [5:0] \level_1_sums[4][93] ;
wire   [5:0] \level_1_sums[4][94] ;
wire   [5:0] \level_1_sums[4][95] ;
wire   [5:0] \level_1_sums[4][96] ;
wire   [5:0] \level_1_sums[4][97] ;
wire   [5:0] \level_1_sums[4][98] ;
wire   [5:0] \level_1_sums[4][99] ;
wire   [5:0] \level_1_sums[4][100] ;
wire   [5:0] \level_1_sums[4][101] ;
wire   [5:0] \level_1_sums[4][102] ;
wire   [5:0] \level_1_sums[4][103] ;
wire   [5:0] \level_1_sums[4][104] ;
wire   [5:0] \level_1_sums[4][105] ;
wire   [5:0] \level_1_sums[4][106] ;
wire   [5:0] \level_1_sums[4][107] ;
wire   [5:0] \level_1_sums[4][108] ;
wire   [5:0] \level_1_sums[4][109] ;
wire   [5:0] \level_1_sums[4][110] ;
wire   [5:0] \level_1_sums[4][111] ;
wire   [5:0] \level_1_sums[4][112] ;
wire   [5:0] \level_1_sums[4][113] ;
wire   [5:0] \level_1_sums[4][114] ;
wire   [5:0] \level_1_sums[4][115] ;
wire   [5:0] \level_1_sums[4][116] ;
wire   [5:0] \level_1_sums[4][117] ;
wire   [5:0] \level_1_sums[4][118] ;
wire   [5:0] \level_1_sums[4][119] ;
wire   [5:0] \level_1_sums[4][120] ;
wire   [5:0] \level_1_sums[4][121] ;
wire   [5:0] \level_1_sums[4][122] ;
wire   [5:0] \level_1_sums[4][123] ;
wire   [5:0] \level_1_sums[4][124] ;
wire   [5:0] \level_1_sums[4][125] ;
wire   [5:0] \level_1_sums[4][126] ;
wire   [5:0] \level_1_sums[4][127] ;
wire   [5:0] \level_1_sums[5][0] ;
wire   [5:0] \level_1_sums[5][1] ;
wire   [5:0] \level_1_sums[5][2] ;
wire   [5:0] \level_1_sums[5][3] ;
wire   [5:0] \level_1_sums[5][4] ;
wire   [5:0] \level_1_sums[5][5] ;
wire   [5:0] \level_1_sums[5][6] ;
wire   [5:0] \level_1_sums[5][7] ;
wire   [5:0] \level_1_sums[5][8] ;
wire   [5:0] \level_1_sums[5][9] ;
wire   [5:0] \level_1_sums[5][10] ;
wire   [5:0] \level_1_sums[5][11] ;
wire   [5:0] \level_1_sums[5][12] ;
wire   [5:0] \level_1_sums[5][13] ;
wire   [5:0] \level_1_sums[5][14] ;
wire   [5:0] \level_1_sums[5][15] ;
wire   [5:0] \level_1_sums[5][16] ;
wire   [5:0] \level_1_sums[5][17] ;
wire   [5:0] \level_1_sums[5][18] ;
wire   [5:0] \level_1_sums[5][19] ;
wire   [5:0] \level_1_sums[5][20] ;
wire   [5:0] \level_1_sums[5][21] ;
wire   [5:0] \level_1_sums[5][22] ;
wire   [5:0] \level_1_sums[5][23] ;
wire   [5:0] \level_1_sums[5][24] ;
wire   [5:0] \level_1_sums[5][25] ;
wire   [5:0] \level_1_sums[5][26] ;
wire   [5:0] \level_1_sums[5][27] ;
wire   [5:0] \level_1_sums[5][28] ;
wire   [5:0] \level_1_sums[5][29] ;
wire   [5:0] \level_1_sums[5][30] ;
wire   [5:0] \level_1_sums[5][31] ;
wire   [5:0] \level_1_sums[5][32] ;
wire   [5:0] \level_1_sums[5][33] ;
wire   [5:0] \level_1_sums[5][34] ;
wire   [5:0] \level_1_sums[5][35] ;
wire   [5:0] \level_1_sums[5][36] ;
wire   [5:0] \level_1_sums[5][37] ;
wire   [5:0] \level_1_sums[5][38] ;
wire   [5:0] \level_1_sums[5][39] ;
wire   [5:0] \level_1_sums[5][40] ;
wire   [5:0] \level_1_sums[5][41] ;
wire   [5:0] \level_1_sums[5][42] ;
wire   [5:0] \level_1_sums[5][43] ;
wire   [5:0] \level_1_sums[5][44] ;
wire   [5:0] \level_1_sums[5][45] ;
wire   [5:0] \level_1_sums[5][46] ;
wire   [5:0] \level_1_sums[5][47] ;
wire   [5:0] \level_1_sums[5][48] ;
wire   [5:0] \level_1_sums[5][49] ;
wire   [5:0] \level_1_sums[5][50] ;
wire   [5:0] \level_1_sums[5][51] ;
wire   [5:0] \level_1_sums[5][52] ;
wire   [5:0] \level_1_sums[5][53] ;
wire   [5:0] \level_1_sums[5][54] ;
wire   [5:0] \level_1_sums[5][55] ;
wire   [5:0] \level_1_sums[5][56] ;
wire   [5:0] \level_1_sums[5][57] ;
wire   [5:0] \level_1_sums[5][58] ;
wire   [5:0] \level_1_sums[5][59] ;
wire   [5:0] \level_1_sums[5][60] ;
wire   [5:0] \level_1_sums[5][61] ;
wire   [5:0] \level_1_sums[5][62] ;
wire   [5:0] \level_1_sums[5][63] ;
wire   [5:0] \level_1_sums[5][64] ;
wire   [5:0] \level_1_sums[5][65] ;
wire   [5:0] \level_1_sums[5][66] ;
wire   [5:0] \level_1_sums[5][67] ;
wire   [5:0] \level_1_sums[5][68] ;
wire   [5:0] \level_1_sums[5][69] ;
wire   [5:0] \level_1_sums[5][70] ;
wire   [5:0] \level_1_sums[5][71] ;
wire   [5:0] \level_1_sums[5][72] ;
wire   [5:0] \level_1_sums[5][73] ;
wire   [5:0] \level_1_sums[5][74] ;
wire   [5:0] \level_1_sums[5][75] ;
wire   [5:0] \level_1_sums[5][76] ;
wire   [5:0] \level_1_sums[5][77] ;
wire   [5:0] \level_1_sums[5][78] ;
wire   [5:0] \level_1_sums[5][79] ;
wire   [5:0] \level_1_sums[5][80] ;
wire   [5:0] \level_1_sums[5][81] ;
wire   [5:0] \level_1_sums[5][82] ;
wire   [5:0] \level_1_sums[5][83] ;
wire   [5:0] \level_1_sums[5][84] ;
wire   [5:0] \level_1_sums[5][85] ;
wire   [5:0] \level_1_sums[5][86] ;
wire   [5:0] \level_1_sums[5][87] ;
wire   [5:0] \level_1_sums[5][88] ;
wire   [5:0] \level_1_sums[5][89] ;
wire   [5:0] \level_1_sums[5][90] ;
wire   [5:0] \level_1_sums[5][91] ;
wire   [5:0] \level_1_sums[5][92] ;
wire   [5:0] \level_1_sums[5][93] ;
wire   [5:0] \level_1_sums[5][94] ;
wire   [5:0] \level_1_sums[5][95] ;
wire   [5:0] \level_1_sums[5][96] ;
wire   [5:0] \level_1_sums[5][97] ;
wire   [5:0] \level_1_sums[5][98] ;
wire   [5:0] \level_1_sums[5][99] ;
wire   [5:0] \level_1_sums[5][100] ;
wire   [5:0] \level_1_sums[5][101] ;
wire   [5:0] \level_1_sums[5][102] ;
wire   [5:0] \level_1_sums[5][103] ;
wire   [5:0] \level_1_sums[5][104] ;
wire   [5:0] \level_1_sums[5][105] ;
wire   [5:0] \level_1_sums[5][106] ;
wire   [5:0] \level_1_sums[5][107] ;
wire   [5:0] \level_1_sums[5][108] ;
wire   [5:0] \level_1_sums[5][109] ;
wire   [5:0] \level_1_sums[5][110] ;
wire   [5:0] \level_1_sums[5][111] ;
wire   [5:0] \level_1_sums[5][112] ;
wire   [5:0] \level_1_sums[5][113] ;
wire   [5:0] \level_1_sums[5][114] ;
wire   [5:0] \level_1_sums[5][115] ;
wire   [5:0] \level_1_sums[5][116] ;
wire   [5:0] \level_1_sums[5][117] ;
wire   [5:0] \level_1_sums[5][118] ;
wire   [5:0] \level_1_sums[5][119] ;
wire   [5:0] \level_1_sums[5][120] ;
wire   [5:0] \level_1_sums[5][121] ;
wire   [5:0] \level_1_sums[5][122] ;
wire   [5:0] \level_1_sums[5][123] ;
wire   [5:0] \level_1_sums[5][124] ;
wire   [5:0] \level_1_sums[5][125] ;
wire   [5:0] \level_1_sums[5][126] ;
wire   [5:0] \level_1_sums[5][127] ;
wire   [5:0] \level_1_sums[6][0] ;
wire   [5:0] \level_1_sums[6][1] ;
wire   [5:0] \level_1_sums[6][2] ;
wire   [5:0] \level_1_sums[6][3] ;
wire   [5:0] \level_1_sums[6][4] ;
wire   [5:0] \level_1_sums[6][5] ;
wire   [5:0] \level_1_sums[6][6] ;
wire   [5:0] \level_1_sums[6][7] ;
wire   [5:0] \level_1_sums[6][8] ;
wire   [5:0] \level_1_sums[6][9] ;
wire   [5:0] \level_1_sums[6][10] ;
wire   [5:0] \level_1_sums[6][11] ;
wire   [5:0] \level_1_sums[6][12] ;
wire   [5:0] \level_1_sums[6][13] ;
wire   [5:0] \level_1_sums[6][14] ;
wire   [5:0] \level_1_sums[6][15] ;
wire   [5:0] \level_1_sums[6][16] ;
wire   [5:0] \level_1_sums[6][17] ;
wire   [5:0] \level_1_sums[6][18] ;
wire   [5:0] \level_1_sums[6][19] ;
wire   [5:0] \level_1_sums[6][20] ;
wire   [5:0] \level_1_sums[6][21] ;
wire   [5:0] \level_1_sums[6][22] ;
wire   [5:0] \level_1_sums[6][23] ;
wire   [5:0] \level_1_sums[6][24] ;
wire   [5:0] \level_1_sums[6][25] ;
wire   [5:0] \level_1_sums[6][26] ;
wire   [5:0] \level_1_sums[6][27] ;
wire   [5:0] \level_1_sums[6][28] ;
wire   [5:0] \level_1_sums[6][29] ;
wire   [5:0] \level_1_sums[6][30] ;
wire   [5:0] \level_1_sums[6][31] ;
wire   [5:0] \level_1_sums[6][32] ;
wire   [5:0] \level_1_sums[6][33] ;
wire   [5:0] \level_1_sums[6][34] ;
wire   [5:0] \level_1_sums[6][35] ;
wire   [5:0] \level_1_sums[6][36] ;
wire   [5:0] \level_1_sums[6][37] ;
wire   [5:0] \level_1_sums[6][38] ;
wire   [5:0] \level_1_sums[6][39] ;
wire   [5:0] \level_1_sums[6][40] ;
wire   [5:0] \level_1_sums[6][41] ;
wire   [5:0] \level_1_sums[6][42] ;
wire   [5:0] \level_1_sums[6][43] ;
wire   [5:0] \level_1_sums[6][44] ;
wire   [5:0] \level_1_sums[6][45] ;
wire   [5:0] \level_1_sums[6][46] ;
wire   [5:0] \level_1_sums[6][47] ;
wire   [5:0] \level_1_sums[6][48] ;
wire   [5:0] \level_1_sums[6][49] ;
wire   [5:0] \level_1_sums[6][50] ;
wire   [5:0] \level_1_sums[6][51] ;
wire   [5:0] \level_1_sums[6][52] ;
wire   [5:0] \level_1_sums[6][53] ;
wire   [5:0] \level_1_sums[6][54] ;
wire   [5:0] \level_1_sums[6][55] ;
wire   [5:0] \level_1_sums[6][56] ;
wire   [5:0] \level_1_sums[6][57] ;
wire   [5:0] \level_1_sums[6][58] ;
wire   [5:0] \level_1_sums[6][59] ;
wire   [5:0] \level_1_sums[6][60] ;
wire   [5:0] \level_1_sums[6][61] ;
wire   [5:0] \level_1_sums[6][62] ;
wire   [5:0] \level_1_sums[6][63] ;
wire   [5:0] \level_1_sums[6][64] ;
wire   [5:0] \level_1_sums[6][65] ;
wire   [5:0] \level_1_sums[6][66] ;
wire   [5:0] \level_1_sums[6][67] ;
wire   [5:0] \level_1_sums[6][68] ;
wire   [5:0] \level_1_sums[6][69] ;
wire   [5:0] \level_1_sums[6][70] ;
wire   [5:0] \level_1_sums[6][71] ;
wire   [5:0] \level_1_sums[6][72] ;
wire   [5:0] \level_1_sums[6][73] ;
wire   [5:0] \level_1_sums[6][74] ;
wire   [5:0] \level_1_sums[6][75] ;
wire   [5:0] \level_1_sums[6][76] ;
wire   [5:0] \level_1_sums[6][77] ;
wire   [5:0] \level_1_sums[6][78] ;
wire   [5:0] \level_1_sums[6][79] ;
wire   [5:0] \level_1_sums[6][80] ;
wire   [5:0] \level_1_sums[6][81] ;
wire   [5:0] \level_1_sums[6][82] ;
wire   [5:0] \level_1_sums[6][83] ;
wire   [5:0] \level_1_sums[6][84] ;
wire   [5:0] \level_1_sums[6][85] ;
wire   [5:0] \level_1_sums[6][86] ;
wire   [5:0] \level_1_sums[6][87] ;
wire   [5:0] \level_1_sums[6][88] ;
wire   [5:0] \level_1_sums[6][89] ;
wire   [5:0] \level_1_sums[6][90] ;
wire   [5:0] \level_1_sums[6][91] ;
wire   [5:0] \level_1_sums[6][92] ;
wire   [5:0] \level_1_sums[6][93] ;
wire   [5:0] \level_1_sums[6][94] ;
wire   [5:0] \level_1_sums[6][95] ;
wire   [5:0] \level_1_sums[6][96] ;
wire   [5:0] \level_1_sums[6][97] ;
wire   [5:0] \level_1_sums[6][98] ;
wire   [5:0] \level_1_sums[6][99] ;
wire   [5:0] \level_1_sums[6][100] ;
wire   [5:0] \level_1_sums[6][101] ;
wire   [5:0] \level_1_sums[6][102] ;
wire   [5:0] \level_1_sums[6][103] ;
wire   [5:0] \level_1_sums[6][104] ;
wire   [5:0] \level_1_sums[6][105] ;
wire   [5:0] \level_1_sums[6][106] ;
wire   [5:0] \level_1_sums[6][107] ;
wire   [5:0] \level_1_sums[6][108] ;
wire   [5:0] \level_1_sums[6][109] ;
wire   [5:0] \level_1_sums[6][110] ;
wire   [5:0] \level_1_sums[6][111] ;
wire   [5:0] \level_1_sums[6][112] ;
wire   [5:0] \level_1_sums[6][113] ;
wire   [5:0] \level_1_sums[6][114] ;
wire   [5:0] \level_1_sums[6][115] ;
wire   [5:0] \level_1_sums[6][116] ;
wire   [5:0] \level_1_sums[6][117] ;
wire   [5:0] \level_1_sums[6][118] ;
wire   [5:0] \level_1_sums[6][119] ;
wire   [5:0] \level_1_sums[6][120] ;
wire   [5:0] \level_1_sums[6][121] ;
wire   [5:0] \level_1_sums[6][122] ;
wire   [5:0] \level_1_sums[6][123] ;
wire   [5:0] \level_1_sums[6][124] ;
wire   [5:0] \level_1_sums[6][125] ;
wire   [5:0] \level_1_sums[6][126] ;
wire   [5:0] \level_1_sums[6][127] ;
wire   [5:0] \level_1_sums[7][0] ;
wire   [5:0] \level_1_sums[7][1] ;
wire   [5:0] \level_1_sums[7][2] ;
wire   [5:0] \level_1_sums[7][3] ;
wire   [5:0] \level_1_sums[7][4] ;
wire   [5:0] \level_1_sums[7][5] ;
wire   [5:0] \level_1_sums[7][6] ;
wire   [5:0] \level_1_sums[7][7] ;
wire   [5:0] \level_1_sums[7][8] ;
wire   [5:0] \level_1_sums[7][9] ;
wire   [5:0] \level_1_sums[7][10] ;
wire   [5:0] \level_1_sums[7][11] ;
wire   [5:0] \level_1_sums[7][12] ;
wire   [5:0] \level_1_sums[7][13] ;
wire   [5:0] \level_1_sums[7][14] ;
wire   [5:0] \level_1_sums[7][15] ;
wire   [5:0] \level_1_sums[7][16] ;
wire   [5:0] \level_1_sums[7][17] ;
wire   [5:0] \level_1_sums[7][18] ;
wire   [5:0] \level_1_sums[7][19] ;
wire   [5:0] \level_1_sums[7][20] ;
wire   [5:0] \level_1_sums[7][21] ;
wire   [5:0] \level_1_sums[7][22] ;
wire   [5:0] \level_1_sums[7][23] ;
wire   [5:0] \level_1_sums[7][24] ;
wire   [5:0] \level_1_sums[7][25] ;
wire   [5:0] \level_1_sums[7][26] ;
wire   [5:0] \level_1_sums[7][27] ;
wire   [5:0] \level_1_sums[7][28] ;
wire   [5:0] \level_1_sums[7][29] ;
wire   [5:0] \level_1_sums[7][30] ;
wire   [5:0] \level_1_sums[7][31] ;
wire   [5:0] \level_1_sums[7][32] ;
wire   [5:0] \level_1_sums[7][33] ;
wire   [5:0] \level_1_sums[7][34] ;
wire   [5:0] \level_1_sums[7][35] ;
wire   [5:0] \level_1_sums[7][36] ;
wire   [5:0] \level_1_sums[7][37] ;
wire   [5:0] \level_1_sums[7][38] ;
wire   [5:0] \level_1_sums[7][39] ;
wire   [5:0] \level_1_sums[7][40] ;
wire   [5:0] \level_1_sums[7][41] ;
wire   [5:0] \level_1_sums[7][42] ;
wire   [5:0] \level_1_sums[7][43] ;
wire   [5:0] \level_1_sums[7][44] ;
wire   [5:0] \level_1_sums[7][45] ;
wire   [5:0] \level_1_sums[7][46] ;
wire   [5:0] \level_1_sums[7][47] ;
wire   [5:0] \level_1_sums[7][48] ;
wire   [5:0] \level_1_sums[7][49] ;
wire   [5:0] \level_1_sums[7][50] ;
wire   [5:0] \level_1_sums[7][51] ;
wire   [5:0] \level_1_sums[7][52] ;
wire   [5:0] \level_1_sums[7][53] ;
wire   [5:0] \level_1_sums[7][54] ;
wire   [5:0] \level_1_sums[7][55] ;
wire   [5:0] \level_1_sums[7][56] ;
wire   [5:0] \level_1_sums[7][57] ;
wire   [5:0] \level_1_sums[7][58] ;
wire   [5:0] \level_1_sums[7][59] ;
wire   [5:0] \level_1_sums[7][60] ;
wire   [5:0] \level_1_sums[7][61] ;
wire   [5:0] \level_1_sums[7][62] ;
wire   [5:0] \level_1_sums[7][63] ;
wire   [5:0] \level_1_sums[7][64] ;
wire   [5:0] \level_1_sums[7][65] ;
wire   [5:0] \level_1_sums[7][66] ;
wire   [5:0] \level_1_sums[7][67] ;
wire   [5:0] \level_1_sums[7][68] ;
wire   [5:0] \level_1_sums[7][69] ;
wire   [5:0] \level_1_sums[7][70] ;
wire   [5:0] \level_1_sums[7][71] ;
wire   [5:0] \level_1_sums[7][72] ;
wire   [5:0] \level_1_sums[7][73] ;
wire   [5:0] \level_1_sums[7][74] ;
wire   [5:0] \level_1_sums[7][75] ;
wire   [5:0] \level_1_sums[7][76] ;
wire   [5:0] \level_1_sums[7][77] ;
wire   [5:0] \level_1_sums[7][78] ;
wire   [5:0] \level_1_sums[7][79] ;
wire   [5:0] \level_1_sums[7][80] ;
wire   [5:0] \level_1_sums[7][81] ;
wire   [5:0] \level_1_sums[7][82] ;
wire   [5:0] \level_1_sums[7][83] ;
wire   [5:0] \level_1_sums[7][84] ;
wire   [5:0] \level_1_sums[7][85] ;
wire   [5:0] \level_1_sums[7][86] ;
wire   [5:0] \level_1_sums[7][87] ;
wire   [5:0] \level_1_sums[7][88] ;
wire   [5:0] \level_1_sums[7][89] ;
wire   [5:0] \level_1_sums[7][90] ;
wire   [5:0] \level_1_sums[7][91] ;
wire   [5:0] \level_1_sums[7][92] ;
wire   [5:0] \level_1_sums[7][93] ;
wire   [5:0] \level_1_sums[7][94] ;
wire   [5:0] \level_1_sums[7][95] ;
wire   [5:0] \level_1_sums[7][96] ;
wire   [5:0] \level_1_sums[7][97] ;
wire   [5:0] \level_1_sums[7][98] ;
wire   [5:0] \level_1_sums[7][99] ;
wire   [5:0] \level_1_sums[7][100] ;
wire   [5:0] \level_1_sums[7][101] ;
wire   [5:0] \level_1_sums[7][102] ;
wire   [5:0] \level_1_sums[7][103] ;
wire   [5:0] \level_1_sums[7][104] ;
wire   [5:0] \level_1_sums[7][105] ;
wire   [5:0] \level_1_sums[7][106] ;
wire   [5:0] \level_1_sums[7][107] ;
wire   [5:0] \level_1_sums[7][108] ;
wire   [5:0] \level_1_sums[7][109] ;
wire   [5:0] \level_1_sums[7][110] ;
wire   [5:0] \level_1_sums[7][111] ;
wire   [5:0] \level_1_sums[7][112] ;
wire   [5:0] \level_1_sums[7][113] ;
wire   [5:0] \level_1_sums[7][114] ;
wire   [5:0] \level_1_sums[7][115] ;
wire   [5:0] \level_1_sums[7][116] ;
wire   [5:0] \level_1_sums[7][117] ;
wire   [5:0] \level_1_sums[7][118] ;
wire   [5:0] \level_1_sums[7][119] ;
wire   [5:0] \level_1_sums[7][120] ;
wire   [5:0] \level_1_sums[7][121] ;
wire   [5:0] \level_1_sums[7][122] ;
wire   [5:0] \level_1_sums[7][123] ;
wire   [5:0] \level_1_sums[7][124] ;
wire   [5:0] \level_1_sums[7][125] ;
wire   [5:0] \level_1_sums[7][126] ;
wire   [5:0] \level_1_sums[7][127] ;
wire   [5:0] \level_1_sums[8][0] ;
wire   [5:0] \level_1_sums[8][1] ;
wire   [5:0] \level_1_sums[8][2] ;
wire   [5:0] \level_1_sums[8][3] ;
wire   [5:0] \level_1_sums[8][4] ;
wire   [5:0] \level_1_sums[8][5] ;
wire   [5:0] \level_1_sums[8][6] ;
wire   [5:0] \level_1_sums[8][7] ;
wire   [5:0] \level_1_sums[8][8] ;
wire   [5:0] \level_1_sums[8][9] ;
wire   [5:0] \level_1_sums[8][10] ;
wire   [5:0] \level_1_sums[8][11] ;
wire   [5:0] \level_1_sums[8][12] ;
wire   [5:0] \level_1_sums[8][13] ;
wire   [5:0] \level_1_sums[8][14] ;
wire   [5:0] \level_1_sums[8][15] ;
wire   [5:0] \level_1_sums[8][16] ;
wire   [5:0] \level_1_sums[8][17] ;
wire   [5:0] \level_1_sums[8][18] ;
wire   [5:0] \level_1_sums[8][19] ;
wire   [5:0] \level_1_sums[8][20] ;
wire   [5:0] \level_1_sums[8][21] ;
wire   [5:0] \level_1_sums[8][22] ;
wire   [5:0] \level_1_sums[8][23] ;
wire   [5:0] \level_1_sums[8][24] ;
wire   [5:0] \level_1_sums[8][25] ;
wire   [5:0] \level_1_sums[8][26] ;
wire   [5:0] \level_1_sums[8][27] ;
wire   [5:0] \level_1_sums[8][28] ;
wire   [5:0] \level_1_sums[8][29] ;
wire   [5:0] \level_1_sums[8][30] ;
wire   [5:0] \level_1_sums[8][31] ;
wire   [5:0] \level_1_sums[8][32] ;
wire   [5:0] \level_1_sums[8][33] ;
wire   [5:0] \level_1_sums[8][34] ;
wire   [5:0] \level_1_sums[8][35] ;
wire   [5:0] \level_1_sums[8][36] ;
wire   [5:0] \level_1_sums[8][37] ;
wire   [5:0] \level_1_sums[8][38] ;
wire   [5:0] \level_1_sums[8][39] ;
wire   [5:0] \level_1_sums[8][40] ;
wire   [5:0] \level_1_sums[8][41] ;
wire   [5:0] \level_1_sums[8][42] ;
wire   [5:0] \level_1_sums[8][43] ;
wire   [5:0] \level_1_sums[8][44] ;
wire   [5:0] \level_1_sums[8][45] ;
wire   [5:0] \level_1_sums[8][46] ;
wire   [5:0] \level_1_sums[8][47] ;
wire   [5:0] \level_1_sums[8][48] ;
wire   [5:0] \level_1_sums[8][49] ;
wire   [5:0] \level_1_sums[8][50] ;
wire   [5:0] \level_1_sums[8][51] ;
wire   [5:0] \level_1_sums[8][52] ;
wire   [5:0] \level_1_sums[8][53] ;
wire   [5:0] \level_1_sums[8][54] ;
wire   [5:0] \level_1_sums[8][55] ;
wire   [5:0] \level_1_sums[8][56] ;
wire   [5:0] \level_1_sums[8][57] ;
wire   [5:0] \level_1_sums[8][58] ;
wire   [5:0] \level_1_sums[8][59] ;
wire   [5:0] \level_1_sums[8][60] ;
wire   [5:0] \level_1_sums[8][61] ;
wire   [5:0] \level_1_sums[8][62] ;
wire   [5:0] \level_1_sums[8][63] ;
wire   [5:0] \level_1_sums[8][64] ;
wire   [5:0] \level_1_sums[8][65] ;
wire   [5:0] \level_1_sums[8][66] ;
wire   [5:0] \level_1_sums[8][67] ;
wire   [5:0] \level_1_sums[8][68] ;
wire   [5:0] \level_1_sums[8][69] ;
wire   [5:0] \level_1_sums[8][70] ;
wire   [5:0] \level_1_sums[8][71] ;
wire   [5:0] \level_1_sums[8][72] ;
wire   [5:0] \level_1_sums[8][73] ;
wire   [5:0] \level_1_sums[8][74] ;
wire   [5:0] \level_1_sums[8][75] ;
wire   [5:0] \level_1_sums[8][76] ;
wire   [5:0] \level_1_sums[8][77] ;
wire   [5:0] \level_1_sums[8][78] ;
wire   [5:0] \level_1_sums[8][79] ;
wire   [5:0] \level_1_sums[8][80] ;
wire   [5:0] \level_1_sums[8][81] ;
wire   [5:0] \level_1_sums[8][82] ;
wire   [5:0] \level_1_sums[8][83] ;
wire   [5:0] \level_1_sums[8][84] ;
wire   [5:0] \level_1_sums[8][85] ;
wire   [5:0] \level_1_sums[8][86] ;
wire   [5:0] \level_1_sums[8][87] ;
wire   [5:0] \level_1_sums[8][88] ;
wire   [5:0] \level_1_sums[8][89] ;
wire   [5:0] \level_1_sums[8][90] ;
wire   [5:0] \level_1_sums[8][91] ;
wire   [5:0] \level_1_sums[8][92] ;
wire   [5:0] \level_1_sums[8][93] ;
wire   [5:0] \level_1_sums[8][94] ;
wire   [5:0] \level_1_sums[8][95] ;
wire   [5:0] \level_1_sums[8][96] ;
wire   [5:0] \level_1_sums[8][97] ;
wire   [5:0] \level_1_sums[8][98] ;
wire   [5:0] \level_1_sums[8][99] ;
wire   [5:0] \level_1_sums[8][100] ;
wire   [5:0] \level_1_sums[8][101] ;
wire   [5:0] \level_1_sums[8][102] ;
wire   [5:0] \level_1_sums[8][103] ;
wire   [5:0] \level_1_sums[8][104] ;
wire   [5:0] \level_1_sums[8][105] ;
wire   [5:0] \level_1_sums[8][106] ;
wire   [5:0] \level_1_sums[8][107] ;
wire   [5:0] \level_1_sums[8][108] ;
wire   [5:0] \level_1_sums[8][109] ;
wire   [5:0] \level_1_sums[8][110] ;
wire   [5:0] \level_1_sums[8][111] ;
wire   [5:0] \level_1_sums[8][112] ;
wire   [5:0] \level_1_sums[8][113] ;
wire   [5:0] \level_1_sums[8][114] ;
wire   [5:0] \level_1_sums[8][115] ;
wire   [5:0] \level_1_sums[8][116] ;
wire   [5:0] \level_1_sums[8][117] ;
wire   [5:0] \level_1_sums[8][118] ;
wire   [5:0] \level_1_sums[8][119] ;
wire   [5:0] \level_1_sums[8][120] ;
wire   [5:0] \level_1_sums[8][121] ;
wire   [5:0] \level_1_sums[8][122] ;
wire   [5:0] \level_1_sums[8][123] ;
wire   [5:0] \level_1_sums[8][124] ;
wire   [5:0] \level_1_sums[8][125] ;
wire   [5:0] \level_1_sums[8][126] ;
wire   [5:0] \level_1_sums[8][127] ;
wire   [5:0] \level_1_sums[9][0] ;
wire   [5:0] \level_1_sums[9][1] ;
wire   [5:0] \level_1_sums[9][2] ;
wire   [5:0] \level_1_sums[9][3] ;
wire   [5:0] \level_1_sums[9][4] ;
wire   [5:0] \level_1_sums[9][5] ;
wire   [5:0] \level_1_sums[9][6] ;
wire   [5:0] \level_1_sums[9][7] ;
wire   [5:0] \level_1_sums[9][8] ;
wire   [5:0] \level_1_sums[9][9] ;
wire   [5:0] \level_1_sums[9][10] ;
wire   [5:0] \level_1_sums[9][11] ;
wire   [5:0] \level_1_sums[9][12] ;
wire   [5:0] \level_1_sums[9][13] ;
wire   [5:0] \level_1_sums[9][14] ;
wire   [5:0] \level_1_sums[9][15] ;
wire   [5:0] \level_1_sums[9][16] ;
wire   [5:0] \level_1_sums[9][17] ;
wire   [5:0] \level_1_sums[9][18] ;
wire   [5:0] \level_1_sums[9][19] ;
wire   [5:0] \level_1_sums[9][20] ;
wire   [5:0] \level_1_sums[9][21] ;
wire   [5:0] \level_1_sums[9][22] ;
wire   [5:0] \level_1_sums[9][23] ;
wire   [5:0] \level_1_sums[9][24] ;
wire   [5:0] \level_1_sums[9][25] ;
wire   [5:0] \level_1_sums[9][26] ;
wire   [5:0] \level_1_sums[9][27] ;
wire   [5:0] \level_1_sums[9][28] ;
wire   [5:0] \level_1_sums[9][29] ;
wire   [5:0] \level_1_sums[9][30] ;
wire   [5:0] \level_1_sums[9][31] ;
wire   [5:0] \level_1_sums[9][32] ;
wire   [5:0] \level_1_sums[9][33] ;
wire   [5:0] \level_1_sums[9][34] ;
wire   [5:0] \level_1_sums[9][35] ;
wire   [5:0] \level_1_sums[9][36] ;
wire   [5:0] \level_1_sums[9][37] ;
wire   [5:0] \level_1_sums[9][38] ;
wire   [5:0] \level_1_sums[9][39] ;
wire   [5:0] \level_1_sums[9][40] ;
wire   [5:0] \level_1_sums[9][41] ;
wire   [5:0] \level_1_sums[9][42] ;
wire   [5:0] \level_1_sums[9][43] ;
wire   [5:0] \level_1_sums[9][44] ;
wire   [5:0] \level_1_sums[9][45] ;
wire   [5:0] \level_1_sums[9][46] ;
wire   [5:0] \level_1_sums[9][47] ;
wire   [5:0] \level_1_sums[9][48] ;
wire   [5:0] \level_1_sums[9][49] ;
wire   [5:0] \level_1_sums[9][50] ;
wire   [5:0] \level_1_sums[9][51] ;
wire   [5:0] \level_1_sums[9][52] ;
wire   [5:0] \level_1_sums[9][53] ;
wire   [5:0] \level_1_sums[9][54] ;
wire   [5:0] \level_1_sums[9][55] ;
wire   [5:0] \level_1_sums[9][56] ;
wire   [5:0] \level_1_sums[9][57] ;
wire   [5:0] \level_1_sums[9][58] ;
wire   [5:0] \level_1_sums[9][59] ;
wire   [5:0] \level_1_sums[9][60] ;
wire   [5:0] \level_1_sums[9][61] ;
wire   [5:0] \level_1_sums[9][62] ;
wire   [5:0] \level_1_sums[9][63] ;
wire   [5:0] \level_1_sums[9][64] ;
wire   [5:0] \level_1_sums[9][65] ;
wire   [5:0] \level_1_sums[9][66] ;
wire   [5:0] \level_1_sums[9][67] ;
wire   [5:0] \level_1_sums[9][68] ;
wire   [5:0] \level_1_sums[9][69] ;
wire   [5:0] \level_1_sums[9][70] ;
wire   [5:0] \level_1_sums[9][71] ;
wire   [5:0] \level_1_sums[9][72] ;
wire   [5:0] \level_1_sums[9][73] ;
wire   [5:0] \level_1_sums[9][74] ;
wire   [5:0] \level_1_sums[9][75] ;
wire   [5:0] \level_1_sums[9][76] ;
wire   [5:0] \level_1_sums[9][77] ;
wire   [5:0] \level_1_sums[9][78] ;
wire   [5:0] \level_1_sums[9][79] ;
wire   [5:0] \level_1_sums[9][80] ;
wire   [5:0] \level_1_sums[9][81] ;
wire   [5:0] \level_1_sums[9][82] ;
wire   [5:0] \level_1_sums[9][83] ;
wire   [5:0] \level_1_sums[9][84] ;
wire   [5:0] \level_1_sums[9][85] ;
wire   [5:0] \level_1_sums[9][86] ;
wire   [5:0] \level_1_sums[9][87] ;
wire   [5:0] \level_1_sums[9][88] ;
wire   [5:0] \level_1_sums[9][89] ;
wire   [5:0] \level_1_sums[9][90] ;
wire   [5:0] \level_1_sums[9][91] ;
wire   [5:0] \level_1_sums[9][92] ;
wire   [5:0] \level_1_sums[9][93] ;
wire   [5:0] \level_1_sums[9][94] ;
wire   [5:0] \level_1_sums[9][95] ;
wire   [5:0] \level_1_sums[9][96] ;
wire   [5:0] \level_1_sums[9][97] ;
wire   [5:0] \level_1_sums[9][98] ;
wire   [5:0] \level_1_sums[9][99] ;
wire   [5:0] \level_1_sums[9][100] ;
wire   [5:0] \level_1_sums[9][101] ;
wire   [5:0] \level_1_sums[9][102] ;
wire   [5:0] \level_1_sums[9][103] ;
wire   [5:0] \level_1_sums[9][104] ;
wire   [5:0] \level_1_sums[9][105] ;
wire   [5:0] \level_1_sums[9][106] ;
wire   [5:0] \level_1_sums[9][107] ;
wire   [5:0] \level_1_sums[9][108] ;
wire   [5:0] \level_1_sums[9][109] ;
wire   [5:0] \level_1_sums[9][110] ;
wire   [5:0] \level_1_sums[9][111] ;
wire   [5:0] \level_1_sums[9][112] ;
wire   [5:0] \level_1_sums[9][113] ;
wire   [5:0] \level_1_sums[9][114] ;
wire   [5:0] \level_1_sums[9][115] ;
wire   [5:0] \level_1_sums[9][116] ;
wire   [5:0] \level_1_sums[9][117] ;
wire   [5:0] \level_1_sums[9][118] ;
wire   [5:0] \level_1_sums[9][119] ;
wire   [5:0] \level_1_sums[9][120] ;
wire   [5:0] \level_1_sums[9][121] ;
wire   [5:0] \level_1_sums[9][122] ;
wire   [5:0] \level_1_sums[9][123] ;
wire   [5:0] \level_1_sums[9][124] ;
wire   [5:0] \level_1_sums[9][125] ;
wire   [5:0] \level_1_sums[9][126] ;
wire   [5:0] \level_1_sums[9][127] ;
wire   [5:0] \level_1_sums[10][0] ;
wire   [5:0] \level_1_sums[10][1] ;
wire   [5:0] \level_1_sums[10][2] ;
wire   [5:0] \level_1_sums[10][3] ;
wire   [5:0] \level_1_sums[10][4] ;
wire   [5:0] \level_1_sums[10][5] ;
wire   [5:0] \level_1_sums[10][6] ;
wire   [5:0] \level_1_sums[10][7] ;
wire   [5:0] \level_1_sums[10][8] ;
wire   [5:0] \level_1_sums[10][9] ;
wire   [5:0] \level_1_sums[10][10] ;
wire   [5:0] \level_1_sums[10][11] ;
wire   [5:0] \level_1_sums[10][12] ;
wire   [5:0] \level_1_sums[10][13] ;
wire   [5:0] \level_1_sums[10][14] ;
wire   [5:0] \level_1_sums[10][15] ;
wire   [5:0] \level_1_sums[10][16] ;
wire   [5:0] \level_1_sums[10][17] ;
wire   [5:0] \level_1_sums[10][18] ;
wire   [5:0] \level_1_sums[10][19] ;
wire   [5:0] \level_1_sums[10][20] ;
wire   [5:0] \level_1_sums[10][21] ;
wire   [5:0] \level_1_sums[10][22] ;
wire   [5:0] \level_1_sums[10][23] ;
wire   [5:0] \level_1_sums[10][24] ;
wire   [5:0] \level_1_sums[10][25] ;
wire   [5:0] \level_1_sums[10][26] ;
wire   [5:0] \level_1_sums[10][27] ;
wire   [5:0] \level_1_sums[10][28] ;
wire   [5:0] \level_1_sums[10][29] ;
wire   [5:0] \level_1_sums[10][30] ;
wire   [5:0] \level_1_sums[10][31] ;
wire   [5:0] \level_1_sums[10][32] ;
wire   [5:0] \level_1_sums[10][33] ;
wire   [5:0] \level_1_sums[10][34] ;
wire   [5:0] \level_1_sums[10][35] ;
wire   [5:0] \level_1_sums[10][36] ;
wire   [5:0] \level_1_sums[10][37] ;
wire   [5:0] \level_1_sums[10][38] ;
wire   [5:0] \level_1_sums[10][39] ;
wire   [5:0] \level_1_sums[10][40] ;
wire   [5:0] \level_1_sums[10][41] ;
wire   [5:0] \level_1_sums[10][42] ;
wire   [5:0] \level_1_sums[10][43] ;
wire   [5:0] \level_1_sums[10][44] ;
wire   [5:0] \level_1_sums[10][45] ;
wire   [5:0] \level_1_sums[10][46] ;
wire   [5:0] \level_1_sums[10][47] ;
wire   [5:0] \level_1_sums[10][48] ;
wire   [5:0] \level_1_sums[10][49] ;
wire   [5:0] \level_1_sums[10][50] ;
wire   [5:0] \level_1_sums[10][51] ;
wire   [5:0] \level_1_sums[10][52] ;
wire   [5:0] \level_1_sums[10][53] ;
wire   [5:0] \level_1_sums[10][54] ;
wire   [5:0] \level_1_sums[10][55] ;
wire   [5:0] \level_1_sums[10][56] ;
wire   [5:0] \level_1_sums[10][57] ;
wire   [5:0] \level_1_sums[10][58] ;
wire   [5:0] \level_1_sums[10][59] ;
wire   [5:0] \level_1_sums[10][60] ;
wire   [5:0] \level_1_sums[10][61] ;
wire   [5:0] \level_1_sums[10][62] ;
wire   [5:0] \level_1_sums[10][63] ;
wire   [5:0] \level_1_sums[10][64] ;
wire   [5:0] \level_1_sums[10][65] ;
wire   [5:0] \level_1_sums[10][66] ;
wire   [5:0] \level_1_sums[10][67] ;
wire   [5:0] \level_1_sums[10][68] ;
wire   [5:0] \level_1_sums[10][69] ;
wire   [5:0] \level_1_sums[10][70] ;
wire   [5:0] \level_1_sums[10][71] ;
wire   [5:0] \level_1_sums[10][72] ;
wire   [5:0] \level_1_sums[10][73] ;
wire   [5:0] \level_1_sums[10][74] ;
wire   [5:0] \level_1_sums[10][75] ;
wire   [5:0] \level_1_sums[10][76] ;
wire   [5:0] \level_1_sums[10][77] ;
wire   [5:0] \level_1_sums[10][78] ;
wire   [5:0] \level_1_sums[10][79] ;
wire   [5:0] \level_1_sums[10][80] ;
wire   [5:0] \level_1_sums[10][81] ;
wire   [5:0] \level_1_sums[10][82] ;
wire   [5:0] \level_1_sums[10][83] ;
wire   [5:0] \level_1_sums[10][84] ;
wire   [5:0] \level_1_sums[10][85] ;
wire   [5:0] \level_1_sums[10][86] ;
wire   [5:0] \level_1_sums[10][87] ;
wire   [5:0] \level_1_sums[10][88] ;
wire   [5:0] \level_1_sums[10][89] ;
wire   [5:0] \level_1_sums[10][90] ;
wire   [5:0] \level_1_sums[10][91] ;
wire   [5:0] \level_1_sums[10][92] ;
wire   [5:0] \level_1_sums[10][93] ;
wire   [5:0] \level_1_sums[10][94] ;
wire   [5:0] \level_1_sums[10][95] ;
wire   [5:0] \level_1_sums[10][96] ;
wire   [5:0] \level_1_sums[10][97] ;
wire   [5:0] \level_1_sums[10][98] ;
wire   [5:0] \level_1_sums[10][99] ;
wire   [5:0] \level_1_sums[10][100] ;
wire   [5:0] \level_1_sums[10][101] ;
wire   [5:0] \level_1_sums[10][102] ;
wire   [5:0] \level_1_sums[10][103] ;
wire   [5:0] \level_1_sums[10][104] ;
wire   [5:0] \level_1_sums[10][105] ;
wire   [5:0] \level_1_sums[10][106] ;
wire   [5:0] \level_1_sums[10][107] ;
wire   [5:0] \level_1_sums[10][108] ;
wire   [5:0] \level_1_sums[10][109] ;
wire   [5:0] \level_1_sums[10][110] ;
wire   [5:0] \level_1_sums[10][111] ;
wire   [5:0] \level_1_sums[10][112] ;
wire   [5:0] \level_1_sums[10][113] ;
wire   [5:0] \level_1_sums[10][114] ;
wire   [5:0] \level_1_sums[10][115] ;
wire   [5:0] \level_1_sums[10][116] ;
wire   [5:0] \level_1_sums[10][117] ;
wire   [5:0] \level_1_sums[10][118] ;
wire   [5:0] \level_1_sums[10][119] ;
wire   [5:0] \level_1_sums[10][120] ;
wire   [5:0] \level_1_sums[10][121] ;
wire   [5:0] \level_1_sums[10][122] ;
wire   [5:0] \level_1_sums[10][123] ;
wire   [5:0] \level_1_sums[10][124] ;
wire   [5:0] \level_1_sums[10][125] ;
wire   [5:0] \level_1_sums[10][126] ;
wire   [5:0] \level_1_sums[10][127] ;
wire   [5:0] \level_1_sums[11][0] ;
wire   [5:0] \level_1_sums[11][1] ;
wire   [5:0] \level_1_sums[11][2] ;
wire   [5:0] \level_1_sums[11][3] ;
wire   [5:0] \level_1_sums[11][4] ;
wire   [5:0] \level_1_sums[11][5] ;
wire   [5:0] \level_1_sums[11][6] ;
wire   [5:0] \level_1_sums[11][7] ;
wire   [5:0] \level_1_sums[11][8] ;
wire   [5:0] \level_1_sums[11][9] ;
wire   [5:0] \level_1_sums[11][10] ;
wire   [5:0] \level_1_sums[11][11] ;
wire   [5:0] \level_1_sums[11][12] ;
wire   [5:0] \level_1_sums[11][13] ;
wire   [5:0] \level_1_sums[11][14] ;
wire   [5:0] \level_1_sums[11][15] ;
wire   [5:0] \level_1_sums[11][16] ;
wire   [5:0] \level_1_sums[11][17] ;
wire   [5:0] \level_1_sums[11][18] ;
wire   [5:0] \level_1_sums[11][19] ;
wire   [5:0] \level_1_sums[11][20] ;
wire   [5:0] \level_1_sums[11][21] ;
wire   [5:0] \level_1_sums[11][22] ;
wire   [5:0] \level_1_sums[11][23] ;
wire   [5:0] \level_1_sums[11][24] ;
wire   [5:0] \level_1_sums[11][25] ;
wire   [5:0] \level_1_sums[11][26] ;
wire   [5:0] \level_1_sums[11][27] ;
wire   [5:0] \level_1_sums[11][28] ;
wire   [5:0] \level_1_sums[11][29] ;
wire   [5:0] \level_1_sums[11][30] ;
wire   [5:0] \level_1_sums[11][31] ;
wire   [5:0] \level_1_sums[11][32] ;
wire   [5:0] \level_1_sums[11][33] ;
wire   [5:0] \level_1_sums[11][34] ;
wire   [5:0] \level_1_sums[11][35] ;
wire   [5:0] \level_1_sums[11][36] ;
wire   [5:0] \level_1_sums[11][37] ;
wire   [5:0] \level_1_sums[11][38] ;
wire   [5:0] \level_1_sums[11][39] ;
wire   [5:0] \level_1_sums[11][40] ;
wire   [5:0] \level_1_sums[11][41] ;
wire   [5:0] \level_1_sums[11][42] ;
wire   [5:0] \level_1_sums[11][43] ;
wire   [5:0] \level_1_sums[11][44] ;
wire   [5:0] \level_1_sums[11][45] ;
wire   [5:0] \level_1_sums[11][46] ;
wire   [5:0] \level_1_sums[11][47] ;
wire   [5:0] \level_1_sums[11][48] ;
wire   [5:0] \level_1_sums[11][49] ;
wire   [5:0] \level_1_sums[11][50] ;
wire   [5:0] \level_1_sums[11][51] ;
wire   [5:0] \level_1_sums[11][52] ;
wire   [5:0] \level_1_sums[11][53] ;
wire   [5:0] \level_1_sums[11][54] ;
wire   [5:0] \level_1_sums[11][55] ;
wire   [5:0] \level_1_sums[11][56] ;
wire   [5:0] \level_1_sums[11][57] ;
wire   [5:0] \level_1_sums[11][58] ;
wire   [5:0] \level_1_sums[11][59] ;
wire   [5:0] \level_1_sums[11][60] ;
wire   [5:0] \level_1_sums[11][61] ;
wire   [5:0] \level_1_sums[11][62] ;
wire   [5:0] \level_1_sums[11][63] ;
wire   [5:0] \level_1_sums[11][64] ;
wire   [5:0] \level_1_sums[11][65] ;
wire   [5:0] \level_1_sums[11][66] ;
wire   [5:0] \level_1_sums[11][67] ;
wire   [5:0] \level_1_sums[11][68] ;
wire   [5:0] \level_1_sums[11][69] ;
wire   [5:0] \level_1_sums[11][70] ;
wire   [5:0] \level_1_sums[11][71] ;
wire   [5:0] \level_1_sums[11][72] ;
wire   [5:0] \level_1_sums[11][73] ;
wire   [5:0] \level_1_sums[11][74] ;
wire   [5:0] \level_1_sums[11][75] ;
wire   [5:0] \level_1_sums[11][76] ;
wire   [5:0] \level_1_sums[11][77] ;
wire   [5:0] \level_1_sums[11][78] ;
wire   [5:0] \level_1_sums[11][79] ;
wire   [5:0] \level_1_sums[11][80] ;
wire   [5:0] \level_1_sums[11][81] ;
wire   [5:0] \level_1_sums[11][82] ;
wire   [5:0] \level_1_sums[11][83] ;
wire   [5:0] \level_1_sums[11][84] ;
wire   [5:0] \level_1_sums[11][85] ;
wire   [5:0] \level_1_sums[11][86] ;
wire   [5:0] \level_1_sums[11][87] ;
wire   [5:0] \level_1_sums[11][88] ;
wire   [5:0] \level_1_sums[11][89] ;
wire   [5:0] \level_1_sums[11][90] ;
wire   [5:0] \level_1_sums[11][91] ;
wire   [5:0] \level_1_sums[11][92] ;
wire   [5:0] \level_1_sums[11][93] ;
wire   [5:0] \level_1_sums[11][94] ;
wire   [5:0] \level_1_sums[11][95] ;
wire   [5:0] \level_1_sums[11][96] ;
wire   [5:0] \level_1_sums[11][97] ;
wire   [5:0] \level_1_sums[11][98] ;
wire   [5:0] \level_1_sums[11][99] ;
wire   [5:0] \level_1_sums[11][100] ;
wire   [5:0] \level_1_sums[11][101] ;
wire   [5:0] \level_1_sums[11][102] ;
wire   [5:0] \level_1_sums[11][103] ;
wire   [5:0] \level_1_sums[11][104] ;
wire   [5:0] \level_1_sums[11][105] ;
wire   [5:0] \level_1_sums[11][106] ;
wire   [5:0] \level_1_sums[11][107] ;
wire   [5:0] \level_1_sums[11][108] ;
wire   [5:0] \level_1_sums[11][109] ;
wire   [5:0] \level_1_sums[11][110] ;
wire   [5:0] \level_1_sums[11][111] ;
wire   [5:0] \level_1_sums[11][112] ;
wire   [5:0] \level_1_sums[11][113] ;
wire   [5:0] \level_1_sums[11][114] ;
wire   [5:0] \level_1_sums[11][115] ;
wire   [5:0] \level_1_sums[11][116] ;
wire   [5:0] \level_1_sums[11][117] ;
wire   [5:0] \level_1_sums[11][118] ;
wire   [5:0] \level_1_sums[11][119] ;
wire   [5:0] \level_1_sums[11][120] ;
wire   [5:0] \level_1_sums[11][121] ;
wire   [5:0] \level_1_sums[11][122] ;
wire   [5:0] \level_1_sums[11][123] ;
wire   [5:0] \level_1_sums[11][124] ;
wire   [5:0] \level_1_sums[11][125] ;
wire   [5:0] \level_1_sums[11][126] ;
wire   [5:0] \level_1_sums[11][127] ;
wire   [5:0] \level_1_sums[12][0] ;
wire   [5:0] \level_1_sums[12][1] ;
wire   [5:0] \level_1_sums[12][2] ;
wire   [5:0] \level_1_sums[12][3] ;
wire   [5:0] \level_1_sums[12][4] ;
wire   [5:0] \level_1_sums[12][5] ;
wire   [5:0] \level_1_sums[12][6] ;
wire   [5:0] \level_1_sums[12][7] ;
wire   [5:0] \level_1_sums[12][8] ;
wire   [5:0] \level_1_sums[12][9] ;
wire   [5:0] \level_1_sums[12][10] ;
wire   [5:0] \level_1_sums[12][11] ;
wire   [5:0] \level_1_sums[12][12] ;
wire   [5:0] \level_1_sums[12][13] ;
wire   [5:0] \level_1_sums[12][14] ;
wire   [5:0] \level_1_sums[12][15] ;
wire   [5:0] \level_1_sums[12][16] ;
wire   [5:0] \level_1_sums[12][17] ;
wire   [5:0] \level_1_sums[12][18] ;
wire   [5:0] \level_1_sums[12][19] ;
wire   [5:0] \level_1_sums[12][20] ;
wire   [5:0] \level_1_sums[12][21] ;
wire   [5:0] \level_1_sums[12][22] ;
wire   [5:0] \level_1_sums[12][23] ;
wire   [5:0] \level_1_sums[12][24] ;
wire   [5:0] \level_1_sums[12][25] ;
wire   [5:0] \level_1_sums[12][26] ;
wire   [5:0] \level_1_sums[12][27] ;
wire   [5:0] \level_1_sums[12][28] ;
wire   [5:0] \level_1_sums[12][29] ;
wire   [5:0] \level_1_sums[12][30] ;
wire   [5:0] \level_1_sums[12][31] ;
wire   [5:0] \level_1_sums[12][32] ;
wire   [5:0] \level_1_sums[12][33] ;
wire   [5:0] \level_1_sums[12][34] ;
wire   [5:0] \level_1_sums[12][35] ;
wire   [5:0] \level_1_sums[12][36] ;
wire   [5:0] \level_1_sums[12][37] ;
wire   [5:0] \level_1_sums[12][38] ;
wire   [5:0] \level_1_sums[12][39] ;
wire   [5:0] \level_1_sums[12][40] ;
wire   [5:0] \level_1_sums[12][41] ;
wire   [5:0] \level_1_sums[12][42] ;
wire   [5:0] \level_1_sums[12][43] ;
wire   [5:0] \level_1_sums[12][44] ;
wire   [5:0] \level_1_sums[12][45] ;
wire   [5:0] \level_1_sums[12][46] ;
wire   [5:0] \level_1_sums[12][47] ;
wire   [5:0] \level_1_sums[12][48] ;
wire   [5:0] \level_1_sums[12][49] ;
wire   [5:0] \level_1_sums[12][50] ;
wire   [5:0] \level_1_sums[12][51] ;
wire   [5:0] \level_1_sums[12][52] ;
wire   [5:0] \level_1_sums[12][53] ;
wire   [5:0] \level_1_sums[12][54] ;
wire   [5:0] \level_1_sums[12][55] ;
wire   [5:0] \level_1_sums[12][56] ;
wire   [5:0] \level_1_sums[12][57] ;
wire   [5:0] \level_1_sums[12][58] ;
wire   [5:0] \level_1_sums[12][59] ;
wire   [5:0] \level_1_sums[12][60] ;
wire   [5:0] \level_1_sums[12][61] ;
wire   [5:0] \level_1_sums[12][62] ;
wire   [5:0] \level_1_sums[12][63] ;
wire   [5:0] \level_1_sums[12][64] ;
wire   [5:0] \level_1_sums[12][65] ;
wire   [5:0] \level_1_sums[12][66] ;
wire   [5:0] \level_1_sums[12][67] ;
wire   [5:0] \level_1_sums[12][68] ;
wire   [5:0] \level_1_sums[12][69] ;
wire   [5:0] \level_1_sums[12][70] ;
wire   [5:0] \level_1_sums[12][71] ;
wire   [5:0] \level_1_sums[12][72] ;
wire   [5:0] \level_1_sums[12][73] ;
wire   [5:0] \level_1_sums[12][74] ;
wire   [5:0] \level_1_sums[12][75] ;
wire   [5:0] \level_1_sums[12][76] ;
wire   [5:0] \level_1_sums[12][77] ;
wire   [5:0] \level_1_sums[12][78] ;
wire   [5:0] \level_1_sums[12][79] ;
wire   [5:0] \level_1_sums[12][80] ;
wire   [5:0] \level_1_sums[12][81] ;
wire   [5:0] \level_1_sums[12][82] ;
wire   [5:0] \level_1_sums[12][83] ;
wire   [5:0] \level_1_sums[12][84] ;
wire   [5:0] \level_1_sums[12][85] ;
wire   [5:0] \level_1_sums[12][86] ;
wire   [5:0] \level_1_sums[12][87] ;
wire   [5:0] \level_1_sums[12][88] ;
wire   [5:0] \level_1_sums[12][89] ;
wire   [5:0] \level_1_sums[12][90] ;
wire   [5:0] \level_1_sums[12][91] ;
wire   [5:0] \level_1_sums[12][92] ;
wire   [5:0] \level_1_sums[12][93] ;
wire   [5:0] \level_1_sums[12][94] ;
wire   [5:0] \level_1_sums[12][95] ;
wire   [5:0] \level_1_sums[12][96] ;
wire   [5:0] \level_1_sums[12][97] ;
wire   [5:0] \level_1_sums[12][98] ;
wire   [5:0] \level_1_sums[12][99] ;
wire   [5:0] \level_1_sums[12][100] ;
wire   [5:0] \level_1_sums[12][101] ;
wire   [5:0] \level_1_sums[12][102] ;
wire   [5:0] \level_1_sums[12][103] ;
wire   [5:0] \level_1_sums[12][104] ;
wire   [5:0] \level_1_sums[12][105] ;
wire   [5:0] \level_1_sums[12][106] ;
wire   [5:0] \level_1_sums[12][107] ;
wire   [5:0] \level_1_sums[12][108] ;
wire   [5:0] \level_1_sums[12][109] ;
wire   [5:0] \level_1_sums[12][110] ;
wire   [5:0] \level_1_sums[12][111] ;
wire   [5:0] \level_1_sums[12][112] ;
wire   [5:0] \level_1_sums[12][113] ;
wire   [5:0] \level_1_sums[12][114] ;
wire   [5:0] \level_1_sums[12][115] ;
wire   [5:0] \level_1_sums[12][116] ;
wire   [5:0] \level_1_sums[12][117] ;
wire   [5:0] \level_1_sums[12][118] ;
wire   [5:0] \level_1_sums[12][119] ;
wire   [5:0] \level_1_sums[12][120] ;
wire   [5:0] \level_1_sums[12][121] ;
wire   [5:0] \level_1_sums[12][122] ;
wire   [5:0] \level_1_sums[12][123] ;
wire   [5:0] \level_1_sums[12][124] ;
wire   [5:0] \level_1_sums[12][125] ;
wire   [5:0] \level_1_sums[12][126] ;
wire   [5:0] \level_1_sums[12][127] ;
wire   [5:0] \level_1_sums[13][0] ;
wire   [5:0] \level_1_sums[13][1] ;
wire   [5:0] \level_1_sums[13][2] ;
wire   [5:0] \level_1_sums[13][3] ;
wire   [5:0] \level_1_sums[13][4] ;
wire   [5:0] \level_1_sums[13][5] ;
wire   [5:0] \level_1_sums[13][6] ;
wire   [5:0] \level_1_sums[13][7] ;
wire   [5:0] \level_1_sums[13][8] ;
wire   [5:0] \level_1_sums[13][9] ;
wire   [5:0] \level_1_sums[13][10] ;
wire   [5:0] \level_1_sums[13][11] ;
wire   [5:0] \level_1_sums[13][12] ;
wire   [5:0] \level_1_sums[13][13] ;
wire   [5:0] \level_1_sums[13][14] ;
wire   [5:0] \level_1_sums[13][15] ;
wire   [5:0] \level_1_sums[13][16] ;
wire   [5:0] \level_1_sums[13][17] ;
wire   [5:0] \level_1_sums[13][18] ;
wire   [5:0] \level_1_sums[13][19] ;
wire   [5:0] \level_1_sums[13][20] ;
wire   [5:0] \level_1_sums[13][21] ;
wire   [5:0] \level_1_sums[13][22] ;
wire   [5:0] \level_1_sums[13][23] ;
wire   [5:0] \level_1_sums[13][24] ;
wire   [5:0] \level_1_sums[13][25] ;
wire   [5:0] \level_1_sums[13][26] ;
wire   [5:0] \level_1_sums[13][27] ;
wire   [5:0] \level_1_sums[13][28] ;
wire   [5:0] \level_1_sums[13][29] ;
wire   [5:0] \level_1_sums[13][30] ;
wire   [5:0] \level_1_sums[13][31] ;
wire   [5:0] \level_1_sums[13][32] ;
wire   [5:0] \level_1_sums[13][33] ;
wire   [5:0] \level_1_sums[13][34] ;
wire   [5:0] \level_1_sums[13][35] ;
wire   [5:0] \level_1_sums[13][36] ;
wire   [5:0] \level_1_sums[13][37] ;
wire   [5:0] \level_1_sums[13][38] ;
wire   [5:0] \level_1_sums[13][39] ;
wire   [5:0] \level_1_sums[13][40] ;
wire   [5:0] \level_1_sums[13][41] ;
wire   [5:0] \level_1_sums[13][42] ;
wire   [5:0] \level_1_sums[13][43] ;
wire   [5:0] \level_1_sums[13][44] ;
wire   [5:0] \level_1_sums[13][45] ;
wire   [5:0] \level_1_sums[13][46] ;
wire   [5:0] \level_1_sums[13][47] ;
wire   [5:0] \level_1_sums[13][48] ;
wire   [5:0] \level_1_sums[13][49] ;
wire   [5:0] \level_1_sums[13][50] ;
wire   [5:0] \level_1_sums[13][51] ;
wire   [5:0] \level_1_sums[13][52] ;
wire   [5:0] \level_1_sums[13][53] ;
wire   [5:0] \level_1_sums[13][54] ;
wire   [5:0] \level_1_sums[13][55] ;
wire   [5:0] \level_1_sums[13][56] ;
wire   [5:0] \level_1_sums[13][57] ;
wire   [5:0] \level_1_sums[13][58] ;
wire   [5:0] \level_1_sums[13][59] ;
wire   [5:0] \level_1_sums[13][60] ;
wire   [5:0] \level_1_sums[13][61] ;
wire   [5:0] \level_1_sums[13][62] ;
wire   [5:0] \level_1_sums[13][63] ;
wire   [5:0] \level_1_sums[13][64] ;
wire   [5:0] \level_1_sums[13][65] ;
wire   [5:0] \level_1_sums[13][66] ;
wire   [5:0] \level_1_sums[13][67] ;
wire   [5:0] \level_1_sums[13][68] ;
wire   [5:0] \level_1_sums[13][69] ;
wire   [5:0] \level_1_sums[13][70] ;
wire   [5:0] \level_1_sums[13][71] ;
wire   [5:0] \level_1_sums[13][72] ;
wire   [5:0] \level_1_sums[13][73] ;
wire   [5:0] \level_1_sums[13][74] ;
wire   [5:0] \level_1_sums[13][75] ;
wire   [5:0] \level_1_sums[13][76] ;
wire   [5:0] \level_1_sums[13][77] ;
wire   [5:0] \level_1_sums[13][78] ;
wire   [5:0] \level_1_sums[13][79] ;
wire   [5:0] \level_1_sums[13][80] ;
wire   [5:0] \level_1_sums[13][81] ;
wire   [5:0] \level_1_sums[13][82] ;
wire   [5:0] \level_1_sums[13][83] ;
wire   [5:0] \level_1_sums[13][84] ;
wire   [5:0] \level_1_sums[13][85] ;
wire   [5:0] \level_1_sums[13][86] ;
wire   [5:0] \level_1_sums[13][87] ;
wire   [5:0] \level_1_sums[13][88] ;
wire   [5:0] \level_1_sums[13][89] ;
wire   [5:0] \level_1_sums[13][90] ;
wire   [5:0] \level_1_sums[13][91] ;
wire   [5:0] \level_1_sums[13][92] ;
wire   [5:0] \level_1_sums[13][93] ;
wire   [5:0] \level_1_sums[13][94] ;
wire   [5:0] \level_1_sums[13][95] ;
wire   [5:0] \level_1_sums[13][96] ;
wire   [5:0] \level_1_sums[13][97] ;
wire   [5:0] \level_1_sums[13][98] ;
wire   [5:0] \level_1_sums[13][99] ;
wire   [5:0] \level_1_sums[13][100] ;
wire   [5:0] \level_1_sums[13][101] ;
wire   [5:0] \level_1_sums[13][102] ;
wire   [5:0] \level_1_sums[13][103] ;
wire   [5:0] \level_1_sums[13][104] ;
wire   [5:0] \level_1_sums[13][105] ;
wire   [5:0] \level_1_sums[13][106] ;
wire   [5:0] \level_1_sums[13][107] ;
wire   [5:0] \level_1_sums[13][108] ;
wire   [5:0] \level_1_sums[13][109] ;
wire   [5:0] \level_1_sums[13][110] ;
wire   [5:0] \level_1_sums[13][111] ;
wire   [5:0] \level_1_sums[13][112] ;
wire   [5:0] \level_1_sums[13][113] ;
wire   [5:0] \level_1_sums[13][114] ;
wire   [5:0] \level_1_sums[13][115] ;
wire   [5:0] \level_1_sums[13][116] ;
wire   [5:0] \level_1_sums[13][117] ;
wire   [5:0] \level_1_sums[13][118] ;
wire   [5:0] \level_1_sums[13][119] ;
wire   [5:0] \level_1_sums[13][120] ;
wire   [5:0] \level_1_sums[13][121] ;
wire   [5:0] \level_1_sums[13][122] ;
wire   [5:0] \level_1_sums[13][123] ;
wire   [5:0] \level_1_sums[13][124] ;
wire   [5:0] \level_1_sums[13][125] ;
wire   [5:0] \level_1_sums[13][126] ;
wire   [5:0] \level_1_sums[13][127] ;
wire   [5:0] \level_1_sums[14][0] ;
wire   [5:0] \level_1_sums[14][1] ;
wire   [5:0] \level_1_sums[14][2] ;
wire   [5:0] \level_1_sums[14][3] ;
wire   [5:0] \level_1_sums[14][4] ;
wire   [5:0] \level_1_sums[14][5] ;
wire   [5:0] \level_1_sums[14][6] ;
wire   [5:0] \level_1_sums[14][7] ;
wire   [5:0] \level_1_sums[14][8] ;
wire   [5:0] \level_1_sums[14][9] ;
wire   [5:0] \level_1_sums[14][10] ;
wire   [5:0] \level_1_sums[14][11] ;
wire   [5:0] \level_1_sums[14][12] ;
wire   [5:0] \level_1_sums[14][13] ;
wire   [5:0] \level_1_sums[14][14] ;
wire   [5:0] \level_1_sums[14][15] ;
wire   [5:0] \level_1_sums[14][16] ;
wire   [5:0] \level_1_sums[14][17] ;
wire   [5:0] \level_1_sums[14][18] ;
wire   [5:0] \level_1_sums[14][19] ;
wire   [5:0] \level_1_sums[14][20] ;
wire   [5:0] \level_1_sums[14][21] ;
wire   [5:0] \level_1_sums[14][22] ;
wire   [5:0] \level_1_sums[14][23] ;
wire   [5:0] \level_1_sums[14][24] ;
wire   [5:0] \level_1_sums[14][25] ;
wire   [5:0] \level_1_sums[14][26] ;
wire   [5:0] \level_1_sums[14][27] ;
wire   [5:0] \level_1_sums[14][28] ;
wire   [5:0] \level_1_sums[14][29] ;
wire   [5:0] \level_1_sums[14][30] ;
wire   [5:0] \level_1_sums[14][31] ;
wire   [5:0] \level_1_sums[14][32] ;
wire   [5:0] \level_1_sums[14][33] ;
wire   [5:0] \level_1_sums[14][34] ;
wire   [5:0] \level_1_sums[14][35] ;
wire   [5:0] \level_1_sums[14][36] ;
wire   [5:0] \level_1_sums[14][37] ;
wire   [5:0] \level_1_sums[14][38] ;
wire   [5:0] \level_1_sums[14][39] ;
wire   [5:0] \level_1_sums[14][40] ;
wire   [5:0] \level_1_sums[14][41] ;
wire   [5:0] \level_1_sums[14][42] ;
wire   [5:0] \level_1_sums[14][43] ;
wire   [5:0] \level_1_sums[14][44] ;
wire   [5:0] \level_1_sums[14][45] ;
wire   [5:0] \level_1_sums[14][46] ;
wire   [5:0] \level_1_sums[14][47] ;
wire   [5:0] \level_1_sums[14][48] ;
wire   [5:0] \level_1_sums[14][49] ;
wire   [5:0] \level_1_sums[14][50] ;
wire   [5:0] \level_1_sums[14][51] ;
wire   [5:0] \level_1_sums[14][52] ;
wire   [5:0] \level_1_sums[14][53] ;
wire   [5:0] \level_1_sums[14][54] ;
wire   [5:0] \level_1_sums[14][55] ;
wire   [5:0] \level_1_sums[14][56] ;
wire   [5:0] \level_1_sums[14][57] ;
wire   [5:0] \level_1_sums[14][58] ;
wire   [5:0] \level_1_sums[14][59] ;
wire   [5:0] \level_1_sums[14][60] ;
wire   [5:0] \level_1_sums[14][61] ;
wire   [5:0] \level_1_sums[14][62] ;
wire   [5:0] \level_1_sums[14][63] ;
wire   [5:0] \level_1_sums[14][64] ;
wire   [5:0] \level_1_sums[14][65] ;
wire   [5:0] \level_1_sums[14][66] ;
wire   [5:0] \level_1_sums[14][67] ;
wire   [5:0] \level_1_sums[14][68] ;
wire   [5:0] \level_1_sums[14][69] ;
wire   [5:0] \level_1_sums[14][70] ;
wire   [5:0] \level_1_sums[14][71] ;
wire   [5:0] \level_1_sums[14][72] ;
wire   [5:0] \level_1_sums[14][73] ;
wire   [5:0] \level_1_sums[14][74] ;
wire   [5:0] \level_1_sums[14][75] ;
wire   [5:0] \level_1_sums[14][76] ;
wire   [5:0] \level_1_sums[14][77] ;
wire   [5:0] \level_1_sums[14][78] ;
wire   [5:0] \level_1_sums[14][79] ;
wire   [5:0] \level_1_sums[14][80] ;
wire   [5:0] \level_1_sums[14][81] ;
wire   [5:0] \level_1_sums[14][82] ;
wire   [5:0] \level_1_sums[14][83] ;
wire   [5:0] \level_1_sums[14][84] ;
wire   [5:0] \level_1_sums[14][85] ;
wire   [5:0] \level_1_sums[14][86] ;
wire   [5:0] \level_1_sums[14][87] ;
wire   [5:0] \level_1_sums[14][88] ;
wire   [5:0] \level_1_sums[14][89] ;
wire   [5:0] \level_1_sums[14][90] ;
wire   [5:0] \level_1_sums[14][91] ;
wire   [5:0] \level_1_sums[14][92] ;
wire   [5:0] \level_1_sums[14][93] ;
wire   [5:0] \level_1_sums[14][94] ;
wire   [5:0] \level_1_sums[14][95] ;
wire   [5:0] \level_1_sums[14][96] ;
wire   [5:0] \level_1_sums[14][97] ;
wire   [5:0] \level_1_sums[14][98] ;
wire   [5:0] \level_1_sums[14][99] ;
wire   [5:0] \level_1_sums[14][100] ;
wire   [5:0] \level_1_sums[14][101] ;
wire   [5:0] \level_1_sums[14][102] ;
wire   [5:0] \level_1_sums[14][103] ;
wire   [5:0] \level_1_sums[14][104] ;
wire   [5:0] \level_1_sums[14][105] ;
wire   [5:0] \level_1_sums[14][106] ;
wire   [5:0] \level_1_sums[14][107] ;
wire   [5:0] \level_1_sums[14][108] ;
wire   [5:0] \level_1_sums[14][109] ;
wire   [5:0] \level_1_sums[14][110] ;
wire   [5:0] \level_1_sums[14][111] ;
wire   [5:0] \level_1_sums[14][112] ;
wire   [5:0] \level_1_sums[14][113] ;
wire   [5:0] \level_1_sums[14][114] ;
wire   [5:0] \level_1_sums[14][115] ;
wire   [5:0] \level_1_sums[14][116] ;
wire   [5:0] \level_1_sums[14][117] ;
wire   [5:0] \level_1_sums[14][118] ;
wire   [5:0] \level_1_sums[14][119] ;
wire   [5:0] \level_1_sums[14][120] ;
wire   [5:0] \level_1_sums[14][121] ;
wire   [5:0] \level_1_sums[14][122] ;
wire   [5:0] \level_1_sums[14][123] ;
wire   [5:0] \level_1_sums[14][124] ;
wire   [5:0] \level_1_sums[14][125] ;
wire   [5:0] \level_1_sums[14][126] ;
wire   [5:0] \level_1_sums[14][127] ;
wire   [5:0] \level_1_sums[15][0] ;
wire   [5:0] \level_1_sums[15][1] ;
wire   [5:0] \level_1_sums[15][2] ;
wire   [5:0] \level_1_sums[15][3] ;
wire   [5:0] \level_1_sums[15][4] ;
wire   [5:0] \level_1_sums[15][5] ;
wire   [5:0] \level_1_sums[15][6] ;
wire   [5:0] \level_1_sums[15][7] ;
wire   [5:0] \level_1_sums[15][8] ;
wire   [5:0] \level_1_sums[15][9] ;
wire   [5:0] \level_1_sums[15][10] ;
wire   [5:0] \level_1_sums[15][11] ;
wire   [5:0] \level_1_sums[15][12] ;
wire   [5:0] \level_1_sums[15][13] ;
wire   [5:0] \level_1_sums[15][14] ;
wire   [5:0] \level_1_sums[15][15] ;
wire   [5:0] \level_1_sums[15][16] ;
wire   [5:0] \level_1_sums[15][17] ;
wire   [5:0] \level_1_sums[15][18] ;
wire   [5:0] \level_1_sums[15][19] ;
wire   [5:0] \level_1_sums[15][20] ;
wire   [5:0] \level_1_sums[15][21] ;
wire   [5:0] \level_1_sums[15][22] ;
wire   [5:0] \level_1_sums[15][23] ;
wire   [5:0] \level_1_sums[15][24] ;
wire   [5:0] \level_1_sums[15][25] ;
wire   [5:0] \level_1_sums[15][26] ;
wire   [5:0] \level_1_sums[15][27] ;
wire   [5:0] \level_1_sums[15][28] ;
wire   [5:0] \level_1_sums[15][29] ;
wire   [5:0] \level_1_sums[15][30] ;
wire   [5:0] \level_1_sums[15][31] ;
wire   [5:0] \level_1_sums[15][32] ;
wire   [5:0] \level_1_sums[15][33] ;
wire   [5:0] \level_1_sums[15][34] ;
wire   [5:0] \level_1_sums[15][35] ;
wire   [5:0] \level_1_sums[15][36] ;
wire   [5:0] \level_1_sums[15][37] ;
wire   [5:0] \level_1_sums[15][38] ;
wire   [5:0] \level_1_sums[15][39] ;
wire   [5:0] \level_1_sums[15][40] ;
wire   [5:0] \level_1_sums[15][41] ;
wire   [5:0] \level_1_sums[15][42] ;
wire   [5:0] \level_1_sums[15][43] ;
wire   [5:0] \level_1_sums[15][44] ;
wire   [5:0] \level_1_sums[15][45] ;
wire   [5:0] \level_1_sums[15][46] ;
wire   [5:0] \level_1_sums[15][47] ;
wire   [5:0] \level_1_sums[15][48] ;
wire   [5:0] \level_1_sums[15][49] ;
wire   [5:0] \level_1_sums[15][50] ;
wire   [5:0] \level_1_sums[15][51] ;
wire   [5:0] \level_1_sums[15][52] ;
wire   [5:0] \level_1_sums[15][53] ;
wire   [5:0] \level_1_sums[15][54] ;
wire   [5:0] \level_1_sums[15][55] ;
wire   [5:0] \level_1_sums[15][56] ;
wire   [5:0] \level_1_sums[15][57] ;
wire   [5:0] \level_1_sums[15][58] ;
wire   [5:0] \level_1_sums[15][59] ;
wire   [5:0] \level_1_sums[15][60] ;
wire   [5:0] \level_1_sums[15][61] ;
wire   [5:0] \level_1_sums[15][62] ;
wire   [5:0] \level_1_sums[15][63] ;
wire   [5:0] \level_1_sums[15][64] ;
wire   [5:0] \level_1_sums[15][65] ;
wire   [5:0] \level_1_sums[15][66] ;
wire   [5:0] \level_1_sums[15][67] ;
wire   [5:0] \level_1_sums[15][68] ;
wire   [5:0] \level_1_sums[15][69] ;
wire   [5:0] \level_1_sums[15][70] ;
wire   [5:0] \level_1_sums[15][71] ;
wire   [5:0] \level_1_sums[15][72] ;
wire   [5:0] \level_1_sums[15][73] ;
wire   [5:0] \level_1_sums[15][74] ;
wire   [5:0] \level_1_sums[15][75] ;
wire   [5:0] \level_1_sums[15][76] ;
wire   [5:0] \level_1_sums[15][77] ;
wire   [5:0] \level_1_sums[15][78] ;
wire   [5:0] \level_1_sums[15][79] ;
wire   [5:0] \level_1_sums[15][80] ;
wire   [5:0] \level_1_sums[15][81] ;
wire   [5:0] \level_1_sums[15][82] ;
wire   [5:0] \level_1_sums[15][83] ;
wire   [5:0] \level_1_sums[15][84] ;
wire   [5:0] \level_1_sums[15][85] ;
wire   [5:0] \level_1_sums[15][86] ;
wire   [5:0] \level_1_sums[15][87] ;
wire   [5:0] \level_1_sums[15][88] ;
wire   [5:0] \level_1_sums[15][89] ;
wire   [5:0] \level_1_sums[15][90] ;
wire   [5:0] \level_1_sums[15][91] ;
wire   [5:0] \level_1_sums[15][92] ;
wire   [5:0] \level_1_sums[15][93] ;
wire   [5:0] \level_1_sums[15][94] ;
wire   [5:0] \level_1_sums[15][95] ;
wire   [5:0] \level_1_sums[15][96] ;
wire   [5:0] \level_1_sums[15][97] ;
wire   [5:0] \level_1_sums[15][98] ;
wire   [5:0] \level_1_sums[15][99] ;
wire   [5:0] \level_1_sums[15][100] ;
wire   [5:0] \level_1_sums[15][101] ;
wire   [5:0] \level_1_sums[15][102] ;
wire   [5:0] \level_1_sums[15][103] ;
wire   [5:0] \level_1_sums[15][104] ;
wire   [5:0] \level_1_sums[15][105] ;
wire   [5:0] \level_1_sums[15][106] ;
wire   [5:0] \level_1_sums[15][107] ;
wire   [5:0] \level_1_sums[15][108] ;
wire   [5:0] \level_1_sums[15][109] ;
wire   [5:0] \level_1_sums[15][110] ;
wire   [5:0] \level_1_sums[15][111] ;
wire   [5:0] \level_1_sums[15][112] ;
wire   [5:0] \level_1_sums[15][113] ;
wire   [5:0] \level_1_sums[15][114] ;
wire   [5:0] \level_1_sums[15][115] ;
wire   [5:0] \level_1_sums[15][116] ;
wire   [5:0] \level_1_sums[15][117] ;
wire   [5:0] \level_1_sums[15][118] ;
wire   [5:0] \level_1_sums[15][119] ;
wire   [5:0] \level_1_sums[15][120] ;
wire   [5:0] \level_1_sums[15][121] ;
wire   [5:0] \level_1_sums[15][122] ;
wire   [5:0] \level_1_sums[15][123] ;
wire   [5:0] \level_1_sums[15][124] ;
wire   [5:0] \level_1_sums[15][125] ;
wire   [5:0] \level_1_sums[15][126] ;
wire   [5:0] \level_1_sums[15][127] ;
wire   [5:0] \level_1_sums[16][0] ;
wire   [5:0] \level_1_sums[16][1] ;
wire   [5:0] \level_1_sums[16][2] ;
wire   [5:0] \level_1_sums[16][3] ;
wire   [5:0] \level_1_sums[16][4] ;
wire   [5:0] \level_1_sums[16][5] ;
wire   [5:0] \level_1_sums[16][6] ;
wire   [5:0] \level_1_sums[16][7] ;
wire   [5:0] \level_1_sums[16][8] ;
wire   [5:0] \level_1_sums[16][9] ;
wire   [5:0] \level_1_sums[16][10] ;
wire   [5:0] \level_1_sums[16][11] ;
wire   [5:0] \level_1_sums[16][12] ;
wire   [5:0] \level_1_sums[16][13] ;
wire   [5:0] \level_1_sums[16][14] ;
wire   [5:0] \level_1_sums[16][15] ;
wire   [5:0] \level_1_sums[16][16] ;
wire   [5:0] \level_1_sums[16][17] ;
wire   [5:0] \level_1_sums[16][18] ;
wire   [5:0] \level_1_sums[16][19] ;
wire   [5:0] \level_1_sums[16][20] ;
wire   [5:0] \level_1_sums[16][21] ;
wire   [5:0] \level_1_sums[16][22] ;
wire   [5:0] \level_1_sums[16][23] ;
wire   [5:0] \level_1_sums[16][24] ;
wire   [5:0] \level_1_sums[16][25] ;
wire   [5:0] \level_1_sums[16][26] ;
wire   [5:0] \level_1_sums[16][27] ;
wire   [5:0] \level_1_sums[16][28] ;
wire   [5:0] \level_1_sums[16][29] ;
wire   [5:0] \level_1_sums[16][30] ;
wire   [5:0] \level_1_sums[16][31] ;
wire   [5:0] \level_1_sums[16][32] ;
wire   [5:0] \level_1_sums[16][33] ;
wire   [5:0] \level_1_sums[16][34] ;
wire   [5:0] \level_1_sums[16][35] ;
wire   [5:0] \level_1_sums[16][36] ;
wire   [5:0] \level_1_sums[16][37] ;
wire   [5:0] \level_1_sums[16][38] ;
wire   [5:0] \level_1_sums[16][39] ;
wire   [5:0] \level_1_sums[16][40] ;
wire   [5:0] \level_1_sums[16][41] ;
wire   [5:0] \level_1_sums[16][42] ;
wire   [5:0] \level_1_sums[16][43] ;
wire   [5:0] \level_1_sums[16][44] ;
wire   [5:0] \level_1_sums[16][45] ;
wire   [5:0] \level_1_sums[16][46] ;
wire   [5:0] \level_1_sums[16][47] ;
wire   [5:0] \level_1_sums[16][48] ;
wire   [5:0] \level_1_sums[16][49] ;
wire   [5:0] \level_1_sums[16][50] ;
wire   [5:0] \level_1_sums[16][51] ;
wire   [5:0] \level_1_sums[16][52] ;
wire   [5:0] \level_1_sums[16][53] ;
wire   [5:0] \level_1_sums[16][54] ;
wire   [5:0] \level_1_sums[16][55] ;
wire   [5:0] \level_1_sums[16][56] ;
wire   [5:0] \level_1_sums[16][57] ;
wire   [5:0] \level_1_sums[16][58] ;
wire   [5:0] \level_1_sums[16][59] ;
wire   [5:0] \level_1_sums[16][60] ;
wire   [5:0] \level_1_sums[16][61] ;
wire   [5:0] \level_1_sums[16][62] ;
wire   [5:0] \level_1_sums[16][63] ;
wire   [5:0] \level_1_sums[16][64] ;
wire   [5:0] \level_1_sums[16][65] ;
wire   [5:0] \level_1_sums[16][66] ;
wire   [5:0] \level_1_sums[16][67] ;
wire   [5:0] \level_1_sums[16][68] ;
wire   [5:0] \level_1_sums[16][69] ;
wire   [5:0] \level_1_sums[16][70] ;
wire   [5:0] \level_1_sums[16][71] ;
wire   [5:0] \level_1_sums[16][72] ;
wire   [5:0] \level_1_sums[16][73] ;
wire   [5:0] \level_1_sums[16][74] ;
wire   [5:0] \level_1_sums[16][75] ;
wire   [5:0] \level_1_sums[16][76] ;
wire   [5:0] \level_1_sums[16][77] ;
wire   [5:0] \level_1_sums[16][78] ;
wire   [5:0] \level_1_sums[16][79] ;
wire   [5:0] \level_1_sums[16][80] ;
wire   [5:0] \level_1_sums[16][81] ;
wire   [5:0] \level_1_sums[16][82] ;
wire   [5:0] \level_1_sums[16][83] ;
wire   [5:0] \level_1_sums[16][84] ;
wire   [5:0] \level_1_sums[16][85] ;
wire   [5:0] \level_1_sums[16][86] ;
wire   [5:0] \level_1_sums[16][87] ;
wire   [5:0] \level_1_sums[16][88] ;
wire   [5:0] \level_1_sums[16][89] ;
wire   [5:0] \level_1_sums[16][90] ;
wire   [5:0] \level_1_sums[16][91] ;
wire   [5:0] \level_1_sums[16][92] ;
wire   [5:0] \level_1_sums[16][93] ;
wire   [5:0] \level_1_sums[16][94] ;
wire   [5:0] \level_1_sums[16][95] ;
wire   [5:0] \level_1_sums[16][96] ;
wire   [5:0] \level_1_sums[16][97] ;
wire   [5:0] \level_1_sums[16][98] ;
wire   [5:0] \level_1_sums[16][99] ;
wire   [5:0] \level_1_sums[16][100] ;
wire   [5:0] \level_1_sums[16][101] ;
wire   [5:0] \level_1_sums[16][102] ;
wire   [5:0] \level_1_sums[16][103] ;
wire   [5:0] \level_1_sums[16][104] ;
wire   [5:0] \level_1_sums[16][105] ;
wire   [5:0] \level_1_sums[16][106] ;
wire   [5:0] \level_1_sums[16][107] ;
wire   [5:0] \level_1_sums[16][108] ;
wire   [5:0] \level_1_sums[16][109] ;
wire   [5:0] \level_1_sums[16][110] ;
wire   [5:0] \level_1_sums[16][111] ;
wire   [5:0] \level_1_sums[16][112] ;
wire   [5:0] \level_1_sums[16][113] ;
wire   [5:0] \level_1_sums[16][114] ;
wire   [5:0] \level_1_sums[16][115] ;
wire   [5:0] \level_1_sums[16][116] ;
wire   [5:0] \level_1_sums[16][117] ;
wire   [5:0] \level_1_sums[16][118] ;
wire   [5:0] \level_1_sums[16][119] ;
wire   [5:0] \level_1_sums[16][120] ;
wire   [5:0] \level_1_sums[16][121] ;
wire   [5:0] \level_1_sums[16][122] ;
wire   [5:0] \level_1_sums[16][123] ;
wire   [5:0] \level_1_sums[16][124] ;
wire   [5:0] \level_1_sums[16][125] ;
wire   [5:0] \level_1_sums[16][126] ;
wire   [5:0] \level_1_sums[16][127] ;
wire   [5:0] \level_1_sums[17][0] ;
wire   [5:0] \level_1_sums[17][1] ;
wire   [5:0] \level_1_sums[17][2] ;
wire   [5:0] \level_1_sums[17][3] ;
wire   [5:0] \level_1_sums[17][4] ;
wire   [5:0] \level_1_sums[17][5] ;
wire   [5:0] \level_1_sums[17][6] ;
wire   [5:0] \level_1_sums[17][7] ;
wire   [5:0] \level_1_sums[17][8] ;
wire   [5:0] \level_1_sums[17][9] ;
wire   [5:0] \level_1_sums[17][10] ;
wire   [5:0] \level_1_sums[17][11] ;
wire   [5:0] \level_1_sums[17][12] ;
wire   [5:0] \level_1_sums[17][13] ;
wire   [5:0] \level_1_sums[17][14] ;
wire   [5:0] \level_1_sums[17][15] ;
wire   [5:0] \level_1_sums[17][16] ;
wire   [5:0] \level_1_sums[17][17] ;
wire   [5:0] \level_1_sums[17][18] ;
wire   [5:0] \level_1_sums[17][19] ;
wire   [5:0] \level_1_sums[17][20] ;
wire   [5:0] \level_1_sums[17][21] ;
wire   [5:0] \level_1_sums[17][22] ;
wire   [5:0] \level_1_sums[17][23] ;
wire   [5:0] \level_1_sums[17][24] ;
wire   [5:0] \level_1_sums[17][25] ;
wire   [5:0] \level_1_sums[17][26] ;
wire   [5:0] \level_1_sums[17][27] ;
wire   [5:0] \level_1_sums[17][28] ;
wire   [5:0] \level_1_sums[17][29] ;
wire   [5:0] \level_1_sums[17][30] ;
wire   [5:0] \level_1_sums[17][31] ;
wire   [5:0] \level_1_sums[17][32] ;
wire   [5:0] \level_1_sums[17][33] ;
wire   [5:0] \level_1_sums[17][34] ;
wire   [5:0] \level_1_sums[17][35] ;
wire   [5:0] \level_1_sums[17][36] ;
wire   [5:0] \level_1_sums[17][37] ;
wire   [5:0] \level_1_sums[17][38] ;
wire   [5:0] \level_1_sums[17][39] ;
wire   [5:0] \level_1_sums[17][40] ;
wire   [5:0] \level_1_sums[17][41] ;
wire   [5:0] \level_1_sums[17][42] ;
wire   [5:0] \level_1_sums[17][43] ;
wire   [5:0] \level_1_sums[17][44] ;
wire   [5:0] \level_1_sums[17][45] ;
wire   [5:0] \level_1_sums[17][46] ;
wire   [5:0] \level_1_sums[17][47] ;
wire   [5:0] \level_1_sums[17][48] ;
wire   [5:0] \level_1_sums[17][49] ;
wire   [5:0] \level_1_sums[17][50] ;
wire   [5:0] \level_1_sums[17][51] ;
wire   [5:0] \level_1_sums[17][52] ;
wire   [5:0] \level_1_sums[17][53] ;
wire   [5:0] \level_1_sums[17][54] ;
wire   [5:0] \level_1_sums[17][55] ;
wire   [5:0] \level_1_sums[17][56] ;
wire   [5:0] \level_1_sums[17][57] ;
wire   [5:0] \level_1_sums[17][58] ;
wire   [5:0] \level_1_sums[17][59] ;
wire   [5:0] \level_1_sums[17][60] ;
wire   [5:0] \level_1_sums[17][61] ;
wire   [5:0] \level_1_sums[17][62] ;
wire   [5:0] \level_1_sums[17][63] ;
wire   [5:0] \level_1_sums[17][64] ;
wire   [5:0] \level_1_sums[17][65] ;
wire   [5:0] \level_1_sums[17][66] ;
wire   [5:0] \level_1_sums[17][67] ;
wire   [5:0] \level_1_sums[17][68] ;
wire   [5:0] \level_1_sums[17][69] ;
wire   [5:0] \level_1_sums[17][70] ;
wire   [5:0] \level_1_sums[17][71] ;
wire   [5:0] \level_1_sums[17][72] ;
wire   [5:0] \level_1_sums[17][73] ;
wire   [5:0] \level_1_sums[17][74] ;
wire   [5:0] \level_1_sums[17][75] ;
wire   [5:0] \level_1_sums[17][76] ;
wire   [5:0] \level_1_sums[17][77] ;
wire   [5:0] \level_1_sums[17][78] ;
wire   [5:0] \level_1_sums[17][79] ;
wire   [5:0] \level_1_sums[17][80] ;
wire   [5:0] \level_1_sums[17][81] ;
wire   [5:0] \level_1_sums[17][82] ;
wire   [5:0] \level_1_sums[17][83] ;
wire   [5:0] \level_1_sums[17][84] ;
wire   [5:0] \level_1_sums[17][85] ;
wire   [5:0] \level_1_sums[17][86] ;
wire   [5:0] \level_1_sums[17][87] ;
wire   [5:0] \level_1_sums[17][88] ;
wire   [5:0] \level_1_sums[17][89] ;
wire   [5:0] \level_1_sums[17][90] ;
wire   [5:0] \level_1_sums[17][91] ;
wire   [5:0] \level_1_sums[17][92] ;
wire   [5:0] \level_1_sums[17][93] ;
wire   [5:0] \level_1_sums[17][94] ;
wire   [5:0] \level_1_sums[17][95] ;
wire   [5:0] \level_1_sums[17][96] ;
wire   [5:0] \level_1_sums[17][97] ;
wire   [5:0] \level_1_sums[17][98] ;
wire   [5:0] \level_1_sums[17][99] ;
wire   [5:0] \level_1_sums[17][100] ;
wire   [5:0] \level_1_sums[17][101] ;
wire   [5:0] \level_1_sums[17][102] ;
wire   [5:0] \level_1_sums[17][103] ;
wire   [5:0] \level_1_sums[17][104] ;
wire   [5:0] \level_1_sums[17][105] ;
wire   [5:0] \level_1_sums[17][106] ;
wire   [5:0] \level_1_sums[17][107] ;
wire   [5:0] \level_1_sums[17][108] ;
wire   [5:0] \level_1_sums[17][109] ;
wire   [5:0] \level_1_sums[17][110] ;
wire   [5:0] \level_1_sums[17][111] ;
wire   [5:0] \level_1_sums[17][112] ;
wire   [5:0] \level_1_sums[17][113] ;
wire   [5:0] \level_1_sums[17][114] ;
wire   [5:0] \level_1_sums[17][115] ;
wire   [5:0] \level_1_sums[17][116] ;
wire   [5:0] \level_1_sums[17][117] ;
wire   [5:0] \level_1_sums[17][118] ;
wire   [5:0] \level_1_sums[17][119] ;
wire   [5:0] \level_1_sums[17][120] ;
wire   [5:0] \level_1_sums[17][121] ;
wire   [5:0] \level_1_sums[17][122] ;
wire   [5:0] \level_1_sums[17][123] ;
wire   [5:0] \level_1_sums[17][124] ;
wire   [5:0] \level_1_sums[17][125] ;
wire   [5:0] \level_1_sums[17][126] ;
wire   [5:0] \level_1_sums[17][127] ;
wire   [5:0] \level_1_sums[18][0] ;
wire   [5:0] \level_1_sums[18][1] ;
wire   [5:0] \level_1_sums[18][2] ;
wire   [5:0] \level_1_sums[18][3] ;
wire   [5:0] \level_1_sums[18][4] ;
wire   [5:0] \level_1_sums[18][5] ;
wire   [5:0] \level_1_sums[18][6] ;
wire   [5:0] \level_1_sums[18][7] ;
wire   [5:0] \level_1_sums[18][8] ;
wire   [5:0] \level_1_sums[18][9] ;
wire   [5:0] \level_1_sums[18][10] ;
wire   [5:0] \level_1_sums[18][11] ;
wire   [5:0] \level_1_sums[18][12] ;
wire   [5:0] \level_1_sums[18][13] ;
wire   [5:0] \level_1_sums[18][14] ;
wire   [5:0] \level_1_sums[18][15] ;
wire   [5:0] \level_1_sums[18][16] ;
wire   [5:0] \level_1_sums[18][17] ;
wire   [5:0] \level_1_sums[18][18] ;
wire   [5:0] \level_1_sums[18][19] ;
wire   [5:0] \level_1_sums[18][20] ;
wire   [5:0] \level_1_sums[18][21] ;
wire   [5:0] \level_1_sums[18][22] ;
wire   [5:0] \level_1_sums[18][23] ;
wire   [5:0] \level_1_sums[18][24] ;
wire   [5:0] \level_1_sums[18][25] ;
wire   [5:0] \level_1_sums[18][26] ;
wire   [5:0] \level_1_sums[18][27] ;
wire   [5:0] \level_1_sums[18][28] ;
wire   [5:0] \level_1_sums[18][29] ;
wire   [5:0] \level_1_sums[18][30] ;
wire   [5:0] \level_1_sums[18][31] ;
wire   [5:0] \level_1_sums[18][32] ;
wire   [5:0] \level_1_sums[18][33] ;
wire   [5:0] \level_1_sums[18][34] ;
wire   [5:0] \level_1_sums[18][35] ;
wire   [5:0] \level_1_sums[18][36] ;
wire   [5:0] \level_1_sums[18][37] ;
wire   [5:0] \level_1_sums[18][38] ;
wire   [5:0] \level_1_sums[18][39] ;
wire   [5:0] \level_1_sums[18][40] ;
wire   [5:0] \level_1_sums[18][41] ;
wire   [5:0] \level_1_sums[18][42] ;
wire   [5:0] \level_1_sums[18][43] ;
wire   [5:0] \level_1_sums[18][44] ;
wire   [5:0] \level_1_sums[18][45] ;
wire   [5:0] \level_1_sums[18][46] ;
wire   [5:0] \level_1_sums[18][47] ;
wire   [5:0] \level_1_sums[18][48] ;
wire   [5:0] \level_1_sums[18][49] ;
wire   [5:0] \level_1_sums[18][50] ;
wire   [5:0] \level_1_sums[18][51] ;
wire   [5:0] \level_1_sums[18][52] ;
wire   [5:0] \level_1_sums[18][53] ;
wire   [5:0] \level_1_sums[18][54] ;
wire   [5:0] \level_1_sums[18][55] ;
wire   [5:0] \level_1_sums[18][56] ;
wire   [5:0] \level_1_sums[18][57] ;
wire   [5:0] \level_1_sums[18][58] ;
wire   [5:0] \level_1_sums[18][59] ;
wire   [5:0] \level_1_sums[18][60] ;
wire   [5:0] \level_1_sums[18][61] ;
wire   [5:0] \level_1_sums[18][62] ;
wire   [5:0] \level_1_sums[18][63] ;
wire   [5:0] \level_1_sums[18][64] ;
wire   [5:0] \level_1_sums[18][65] ;
wire   [5:0] \level_1_sums[18][66] ;
wire   [5:0] \level_1_sums[18][67] ;
wire   [5:0] \level_1_sums[18][68] ;
wire   [5:0] \level_1_sums[18][69] ;
wire   [5:0] \level_1_sums[18][70] ;
wire   [5:0] \level_1_sums[18][71] ;
wire   [5:0] \level_1_sums[18][72] ;
wire   [5:0] \level_1_sums[18][73] ;
wire   [5:0] \level_1_sums[18][74] ;
wire   [5:0] \level_1_sums[18][75] ;
wire   [5:0] \level_1_sums[18][76] ;
wire   [5:0] \level_1_sums[18][77] ;
wire   [5:0] \level_1_sums[18][78] ;
wire   [5:0] \level_1_sums[18][79] ;
wire   [5:0] \level_1_sums[18][80] ;
wire   [5:0] \level_1_sums[18][81] ;
wire   [5:0] \level_1_sums[18][82] ;
wire   [5:0] \level_1_sums[18][83] ;
wire   [5:0] \level_1_sums[18][84] ;
wire   [5:0] \level_1_sums[18][85] ;
wire   [5:0] \level_1_sums[18][86] ;
wire   [5:0] \level_1_sums[18][87] ;
wire   [5:0] \level_1_sums[18][88] ;
wire   [5:0] \level_1_sums[18][89] ;
wire   [5:0] \level_1_sums[18][90] ;
wire   [5:0] \level_1_sums[18][91] ;
wire   [5:0] \level_1_sums[18][92] ;
wire   [5:0] \level_1_sums[18][93] ;
wire   [5:0] \level_1_sums[18][94] ;
wire   [5:0] \level_1_sums[18][95] ;
wire   [5:0] \level_1_sums[18][96] ;
wire   [5:0] \level_1_sums[18][97] ;
wire   [5:0] \level_1_sums[18][98] ;
wire   [5:0] \level_1_sums[18][99] ;
wire   [5:0] \level_1_sums[18][100] ;
wire   [5:0] \level_1_sums[18][101] ;
wire   [5:0] \level_1_sums[18][102] ;
wire   [5:0] \level_1_sums[18][103] ;
wire   [5:0] \level_1_sums[18][104] ;
wire   [5:0] \level_1_sums[18][105] ;
wire   [5:0] \level_1_sums[18][106] ;
wire   [5:0] \level_1_sums[18][107] ;
wire   [5:0] \level_1_sums[18][108] ;
wire   [5:0] \level_1_sums[18][109] ;
wire   [5:0] \level_1_sums[18][110] ;
wire   [5:0] \level_1_sums[18][111] ;
wire   [5:0] \level_1_sums[18][112] ;
wire   [5:0] \level_1_sums[18][113] ;
wire   [5:0] \level_1_sums[18][114] ;
wire   [5:0] \level_1_sums[18][115] ;
wire   [5:0] \level_1_sums[18][116] ;
wire   [5:0] \level_1_sums[18][117] ;
wire   [5:0] \level_1_sums[18][118] ;
wire   [5:0] \level_1_sums[18][119] ;
wire   [5:0] \level_1_sums[18][120] ;
wire   [5:0] \level_1_sums[18][121] ;
wire   [5:0] \level_1_sums[18][122] ;
wire   [5:0] \level_1_sums[18][123] ;
wire   [5:0] \level_1_sums[18][124] ;
wire   [5:0] \level_1_sums[18][125] ;
wire   [5:0] \level_1_sums[18][126] ;
wire   [5:0] \level_1_sums[18][127] ;
wire   [5:0] \level_1_sums[19][0] ;
wire   [5:0] \level_1_sums[19][1] ;
wire   [5:0] \level_1_sums[19][2] ;
wire   [5:0] \level_1_sums[19][3] ;
wire   [5:0] \level_1_sums[19][4] ;
wire   [5:0] \level_1_sums[19][5] ;
wire   [5:0] \level_1_sums[19][6] ;
wire   [5:0] \level_1_sums[19][7] ;
wire   [5:0] \level_1_sums[19][8] ;
wire   [5:0] \level_1_sums[19][9] ;
wire   [5:0] \level_1_sums[19][10] ;
wire   [5:0] \level_1_sums[19][11] ;
wire   [5:0] \level_1_sums[19][12] ;
wire   [5:0] \level_1_sums[19][13] ;
wire   [5:0] \level_1_sums[19][14] ;
wire   [5:0] \level_1_sums[19][15] ;
wire   [5:0] \level_1_sums[19][16] ;
wire   [5:0] \level_1_sums[19][17] ;
wire   [5:0] \level_1_sums[19][18] ;
wire   [5:0] \level_1_sums[19][19] ;
wire   [5:0] \level_1_sums[19][20] ;
wire   [5:0] \level_1_sums[19][21] ;
wire   [5:0] \level_1_sums[19][22] ;
wire   [5:0] \level_1_sums[19][23] ;
wire   [5:0] \level_1_sums[19][24] ;
wire   [5:0] \level_1_sums[19][25] ;
wire   [5:0] \level_1_sums[19][26] ;
wire   [5:0] \level_1_sums[19][27] ;
wire   [5:0] \level_1_sums[19][28] ;
wire   [5:0] \level_1_sums[19][29] ;
wire   [5:0] \level_1_sums[19][30] ;
wire   [5:0] \level_1_sums[19][31] ;
wire   [5:0] \level_1_sums[19][32] ;
wire   [5:0] \level_1_sums[19][33] ;
wire   [5:0] \level_1_sums[19][34] ;
wire   [5:0] \level_1_sums[19][35] ;
wire   [5:0] \level_1_sums[19][36] ;
wire   [5:0] \level_1_sums[19][37] ;
wire   [5:0] \level_1_sums[19][38] ;
wire   [5:0] \level_1_sums[19][39] ;
wire   [5:0] \level_1_sums[19][40] ;
wire   [5:0] \level_1_sums[19][41] ;
wire   [5:0] \level_1_sums[19][42] ;
wire   [5:0] \level_1_sums[19][43] ;
wire   [5:0] \level_1_sums[19][44] ;
wire   [5:0] \level_1_sums[19][45] ;
wire   [5:0] \level_1_sums[19][46] ;
wire   [5:0] \level_1_sums[19][47] ;
wire   [5:0] \level_1_sums[19][48] ;
wire   [5:0] \level_1_sums[19][49] ;
wire   [5:0] \level_1_sums[19][50] ;
wire   [5:0] \level_1_sums[19][51] ;
wire   [5:0] \level_1_sums[19][52] ;
wire   [5:0] \level_1_sums[19][53] ;
wire   [5:0] \level_1_sums[19][54] ;
wire   [5:0] \level_1_sums[19][55] ;
wire   [5:0] \level_1_sums[19][56] ;
wire   [5:0] \level_1_sums[19][57] ;
wire   [5:0] \level_1_sums[19][58] ;
wire   [5:0] \level_1_sums[19][59] ;
wire   [5:0] \level_1_sums[19][60] ;
wire   [5:0] \level_1_sums[19][61] ;
wire   [5:0] \level_1_sums[19][62] ;
wire   [5:0] \level_1_sums[19][63] ;
wire   [5:0] \level_1_sums[19][64] ;
wire   [5:0] \level_1_sums[19][65] ;
wire   [5:0] \level_1_sums[19][66] ;
wire   [5:0] \level_1_sums[19][67] ;
wire   [5:0] \level_1_sums[19][68] ;
wire   [5:0] \level_1_sums[19][69] ;
wire   [5:0] \level_1_sums[19][70] ;
wire   [5:0] \level_1_sums[19][71] ;
wire   [5:0] \level_1_sums[19][72] ;
wire   [5:0] \level_1_sums[19][73] ;
wire   [5:0] \level_1_sums[19][74] ;
wire   [5:0] \level_1_sums[19][75] ;
wire   [5:0] \level_1_sums[19][76] ;
wire   [5:0] \level_1_sums[19][77] ;
wire   [5:0] \level_1_sums[19][78] ;
wire   [5:0] \level_1_sums[19][79] ;
wire   [5:0] \level_1_sums[19][80] ;
wire   [5:0] \level_1_sums[19][81] ;
wire   [5:0] \level_1_sums[19][82] ;
wire   [5:0] \level_1_sums[19][83] ;
wire   [5:0] \level_1_sums[19][84] ;
wire   [5:0] \level_1_sums[19][85] ;
wire   [5:0] \level_1_sums[19][86] ;
wire   [5:0] \level_1_sums[19][87] ;
wire   [5:0] \level_1_sums[19][88] ;
wire   [5:0] \level_1_sums[19][89] ;
wire   [5:0] \level_1_sums[19][90] ;
wire   [5:0] \level_1_sums[19][91] ;
wire   [5:0] \level_1_sums[19][92] ;
wire   [5:0] \level_1_sums[19][93] ;
wire   [5:0] \level_1_sums[19][94] ;
wire   [5:0] \level_1_sums[19][95] ;
wire   [5:0] \level_1_sums[19][96] ;
wire   [5:0] \level_1_sums[19][97] ;
wire   [5:0] \level_1_sums[19][98] ;
wire   [5:0] \level_1_sums[19][99] ;
wire   [5:0] \level_1_sums[19][100] ;
wire   [5:0] \level_1_sums[19][101] ;
wire   [5:0] \level_1_sums[19][102] ;
wire   [5:0] \level_1_sums[19][103] ;
wire   [5:0] \level_1_sums[19][104] ;
wire   [5:0] \level_1_sums[19][105] ;
wire   [5:0] \level_1_sums[19][106] ;
wire   [5:0] \level_1_sums[19][107] ;
wire   [5:0] \level_1_sums[19][108] ;
wire   [5:0] \level_1_sums[19][109] ;
wire   [5:0] \level_1_sums[19][110] ;
wire   [5:0] \level_1_sums[19][111] ;
wire   [5:0] \level_1_sums[19][112] ;
wire   [5:0] \level_1_sums[19][113] ;
wire   [5:0] \level_1_sums[19][114] ;
wire   [5:0] \level_1_sums[19][115] ;
wire   [5:0] \level_1_sums[19][116] ;
wire   [5:0] \level_1_sums[19][117] ;
wire   [5:0] \level_1_sums[19][118] ;
wire   [5:0] \level_1_sums[19][119] ;
wire   [5:0] \level_1_sums[19][120] ;
wire   [5:0] \level_1_sums[19][121] ;
wire   [5:0] \level_1_sums[19][122] ;
wire   [5:0] \level_1_sums[19][123] ;
wire   [5:0] \level_1_sums[19][124] ;
wire   [5:0] \level_1_sums[19][125] ;
wire   [5:0] \level_1_sums[19][126] ;
wire   [5:0] \level_1_sums[19][127] ;
wire   [9:0] \biases_l1_ext[0] ;
wire   [9:0] \biases_l1_ext[1] ;
wire   [9:0] \biases_l1_ext[2] ;
wire   [9:0] \biases_l1_ext[3] ;
wire   [9:0] \biases_l1_ext[4] ;
wire   [9:0] \biases_l1_ext[5] ;
wire   [9:0] \biases_l1_ext[6] ;
wire   [9:0] \biases_l1_ext[7] ;
wire   [9:0] \biases_l1_ext[8] ;
wire   [9:0] \biases_l1_ext[9] ;
wire   [9:0] \biases_l1_ext[10] ;
wire   [9:0] \biases_l1_ext[11] ;
wire   [9:0] \biases_l1_ext[12] ;
wire   [9:0] \biases_l1_ext[13] ;
wire   [9:0] \biases_l1_ext[14] ;
wire   [9:0] \biases_l1_ext[15] ;
wire   [9:0] \biases_l1_ext[16] ;
wire   [9:0] \biases_l1_ext[17] ;
wire   [9:0] \biases_l1_ext[18] ;
wire   [9:0] \biases_l1_ext[19] ;
wire   [6:0] \biases_l1[0] ;
wire   [6:0] \biases_l1[1] ;
wire   [6:0] \biases_l1[2] ;
wire   [6:0] \biases_l1[3] ;
wire   [6:0] \biases_l1[4] ;
wire   [6:0] \biases_l1[5] ;
wire   [6:0] \biases_l1[6] ;
wire   [6:0] \biases_l1[7] ;
wire   [6:0] \biases_l1[8] ;
wire   [6:0] \biases_l1[9] ;
wire   [6:0] \biases_l1[10] ;
wire   [6:0] \biases_l1[11] ;
wire   [6:0] \biases_l1[12] ;
wire   [6:0] \biases_l1[13] ;
wire   [6:0] \biases_l1[14] ;
wire   [6:0] \biases_l1[15] ;
wire   [6:0] \biases_l1[16] ;
wire   [6:0] \biases_l1[17] ;
wire   [6:0] \biases_l1[18] ;
wire   [6:0] \biases_l1[19] ;
wire   [4:0] \A[0][0] ;
wire   [4:0] \A[0][1] ;
wire   [4:0] \A[0][2] ;
wire   [4:0] \A[0][3] ;
wire   [4:0] \A[0][4] ;
wire   [4:0] \A[0][5] ;
wire   [4:0] \A[0][6] ;
wire   [4:0] \A[0][7] ;
wire   [4:0] \A[0][8] ;
wire   [4:0] \A[0][9] ;
wire   [4:0] \A[0][10] ;
wire   [4:0] \A[0][11] ;
wire   [4:0] \A[0][12] ;
wire   [4:0] \A[0][13] ;
wire   [4:0] \A[0][14] ;
wire   [4:0] \A[0][15] ;
wire   [4:0] \A[0][16] ;
wire   [4:0] \A[0][17] ;
wire   [4:0] \A[0][18] ;
wire   [4:0] \A[0][19] ;
wire   [4:0] \A[0][20] ;
wire   [4:0] \A[0][21] ;
wire   [4:0] \A[0][22] ;
wire   [4:0] \A[0][23] ;
wire   [4:0] \A[0][24] ;
wire   [4:0] \A[0][25] ;
wire   [4:0] \A[0][26] ;
wire   [4:0] \A[0][27] ;
wire   [4:0] \A[0][28] ;
wire   [4:0] \A[0][29] ;
wire   [4:0] \A[0][30] ;
wire   [4:0] \A[0][31] ;
wire   [4:0] \A[0][32] ;
wire   [4:0] \A[0][33] ;
wire   [4:0] \A[0][34] ;
wire   [4:0] \A[0][35] ;
wire   [4:0] \A[0][36] ;
wire   [4:0] \A[0][37] ;
wire   [4:0] \A[0][38] ;
wire   [4:0] \A[0][39] ;
wire   [4:0] \A[0][40] ;
wire   [4:0] \A[0][41] ;
wire   [4:0] \A[0][42] ;
wire   [4:0] \A[0][43] ;
wire   [4:0] \A[0][44] ;
wire   [4:0] \A[0][45] ;
wire   [4:0] \A[0][46] ;
wire   [4:0] \A[0][47] ;
wire   [4:0] \A[0][48] ;
wire   [4:0] \A[0][49] ;
wire   [4:0] \A[0][50] ;
wire   [4:0] \A[0][51] ;
wire   [4:0] \A[0][52] ;
wire   [4:0] \A[0][53] ;
wire   [4:0] \A[0][54] ;
wire   [4:0] \A[0][55] ;
wire   [4:0] \A[0][56] ;
wire   [4:0] \A[0][57] ;
wire   [4:0] \A[0][58] ;
wire   [4:0] \A[0][59] ;
wire   [4:0] \A[0][60] ;
wire   [4:0] \A[0][61] ;
wire   [4:0] \A[0][62] ;
wire   [4:0] \A[0][63] ;
wire   [4:0] \A[0][64] ;
wire   [4:0] \A[0][65] ;
wire   [4:0] \A[0][66] ;
wire   [4:0] \A[0][67] ;
wire   [4:0] \A[0][68] ;
wire   [4:0] \A[0][69] ;
wire   [4:0] \A[0][70] ;
wire   [4:0] \A[0][71] ;
wire   [4:0] \A[0][72] ;
wire   [4:0] \A[0][73] ;
wire   [4:0] \A[0][74] ;
wire   [4:0] \A[0][75] ;
wire   [4:0] \A[0][76] ;
wire   [4:0] \A[0][77] ;
wire   [4:0] \A[0][78] ;
wire   [4:0] \A[0][79] ;
wire   [4:0] \A[0][80] ;
wire   [4:0] \A[0][81] ;
wire   [4:0] \A[0][82] ;
wire   [4:0] \A[0][83] ;
wire   [4:0] \A[0][84] ;
wire   [4:0] \A[0][85] ;
wire   [4:0] \A[0][86] ;
wire   [4:0] \A[0][87] ;
wire   [4:0] \A[0][88] ;
wire   [4:0] \A[0][89] ;
wire   [4:0] \A[0][90] ;
wire   [4:0] \A[0][91] ;
wire   [4:0] \A[0][92] ;
wire   [4:0] \A[0][93] ;
wire   [4:0] \A[0][94] ;
wire   [4:0] \A[0][95] ;
wire   [4:0] \A[0][96] ;
wire   [4:0] \A[0][97] ;
wire   [4:0] \A[0][98] ;
wire   [4:0] \A[0][99] ;
wire   [4:0] \A[0][100] ;
wire   [4:0] \A[0][101] ;
wire   [4:0] \A[0][102] ;
wire   [4:0] \A[0][103] ;
wire   [4:0] \A[0][104] ;
wire   [4:0] \A[0][105] ;
wire   [4:0] \A[0][106] ;
wire   [4:0] \A[0][107] ;
wire   [4:0] \A[0][108] ;
wire   [4:0] \A[0][109] ;
wire   [4:0] \A[0][110] ;
wire   [4:0] \A[0][111] ;
wire   [4:0] \A[0][112] ;
wire   [4:0] \A[0][113] ;
wire   [4:0] \A[0][114] ;
wire   [4:0] \A[0][115] ;
wire   [4:0] \A[0][116] ;
wire   [4:0] \A[0][117] ;
wire   [4:0] \A[0][118] ;
wire   [4:0] \A[0][119] ;
wire   [4:0] \A[0][120] ;
wire   [4:0] \A[0][121] ;
wire   [4:0] \A[0][122] ;
wire   [4:0] \A[0][123] ;
wire   [4:0] \A[0][124] ;
wire   [4:0] \A[0][125] ;
wire   [4:0] \A[0][126] ;
wire   [4:0] \A[0][127] ;
wire   [4:0] \A[0][128] ;
wire   [4:0] \A[0][129] ;
wire   [4:0] \A[0][130] ;
wire   [4:0] \A[0][131] ;
wire   [4:0] \A[0][132] ;
wire   [4:0] \A[0][133] ;
wire   [4:0] \A[0][134] ;
wire   [4:0] \A[0][135] ;
wire   [4:0] \A[0][136] ;
wire   [4:0] \A[0][137] ;
wire   [4:0] \A[0][138] ;
wire   [4:0] \A[0][139] ;
wire   [4:0] \A[0][140] ;
wire   [4:0] \A[0][141] ;
wire   [4:0] \A[0][142] ;
wire   [4:0] \A[0][143] ;
wire   [4:0] \A[0][144] ;
wire   [4:0] \A[0][145] ;
wire   [4:0] \A[0][146] ;
wire   [4:0] \A[0][147] ;
wire   [4:0] \A[0][148] ;
wire   [4:0] \A[0][149] ;
wire   [4:0] \A[0][150] ;
wire   [4:0] \A[0][151] ;
wire   [4:0] \A[0][152] ;
wire   [4:0] \A[0][153] ;
wire   [4:0] \A[0][154] ;
wire   [4:0] \A[0][155] ;
wire   [4:0] \A[0][156] ;
wire   [4:0] \A[0][157] ;
wire   [4:0] \A[0][158] ;
wire   [4:0] \A[0][159] ;
wire   [4:0] \A[0][160] ;
wire   [4:0] \A[0][161] ;
wire   [4:0] \A[0][162] ;
wire   [4:0] \A[0][163] ;
wire   [4:0] \A[0][164] ;
wire   [4:0] \A[0][165] ;
wire   [4:0] \A[0][166] ;
wire   [4:0] \A[0][167] ;
wire   [4:0] \A[0][168] ;
wire   [4:0] \A[0][169] ;
wire   [4:0] \A[0][170] ;
wire   [4:0] \A[0][171] ;
wire   [4:0] \A[0][172] ;
wire   [4:0] \A[0][173] ;
wire   [4:0] \A[0][174] ;
wire   [4:0] \A[0][175] ;
wire   [4:0] \A[0][176] ;
wire   [4:0] \A[0][177] ;
wire   [4:0] \A[0][178] ;
wire   [4:0] \A[0][179] ;
wire   [4:0] \A[0][180] ;
wire   [4:0] \A[0][181] ;
wire   [4:0] \A[0][182] ;
wire   [4:0] \A[0][183] ;
wire   [4:0] \A[0][184] ;
wire   [4:0] \A[0][185] ;
wire   [4:0] \A[0][186] ;
wire   [4:0] \A[0][187] ;
wire   [4:0] \A[0][188] ;
wire   [4:0] \A[0][189] ;
wire   [4:0] \A[0][190] ;
wire   [4:0] \A[0][191] ;
wire   [4:0] \A[0][192] ;
wire   [4:0] \A[0][193] ;
wire   [4:0] \A[0][194] ;
wire   [4:0] \A[0][195] ;
wire   [4:0] \A[0][196] ;
wire   [4:0] \A[0][197] ;
wire   [4:0] \A[0][198] ;
wire   [4:0] \A[0][199] ;
wire   [4:0] \A[0][200] ;
wire   [4:0] \A[0][201] ;
wire   [4:0] \A[0][202] ;
wire   [4:0] \A[0][203] ;
wire   [4:0] \A[0][204] ;
wire   [4:0] \A[0][205] ;
wire   [4:0] \A[0][206] ;
wire   [4:0] \A[0][207] ;
wire   [4:0] \A[0][208] ;
wire   [4:0] \A[0][209] ;
wire   [4:0] \A[0][210] ;
wire   [4:0] \A[0][211] ;
wire   [4:0] \A[0][212] ;
wire   [4:0] \A[0][213] ;
wire   [4:0] \A[0][214] ;
wire   [4:0] \A[0][215] ;
wire   [4:0] \A[0][216] ;
wire   [4:0] \A[0][217] ;
wire   [4:0] \A[0][218] ;
wire   [4:0] \A[0][219] ;
wire   [4:0] \A[0][220] ;
wire   [4:0] \A[0][221] ;
wire   [4:0] \A[0][222] ;
wire   [4:0] \A[0][223] ;
wire   [4:0] \A[0][224] ;
wire   [4:0] \A[0][225] ;
wire   [4:0] \A[0][226] ;
wire   [4:0] \A[0][227] ;
wire   [4:0] \A[0][228] ;
wire   [4:0] \A[0][229] ;
wire   [4:0] \A[0][230] ;
wire   [4:0] \A[0][231] ;
wire   [4:0] \A[0][232] ;
wire   [4:0] \A[0][233] ;
wire   [4:0] \A[0][234] ;
wire   [4:0] \A[0][235] ;
wire   [4:0] \A[0][236] ;
wire   [4:0] \A[0][237] ;
wire   [4:0] \A[0][238] ;
wire   [4:0] \A[0][239] ;
wire   [4:0] \A[0][240] ;
wire   [4:0] \A[0][241] ;
wire   [4:0] \A[0][242] ;
wire   [4:0] \A[0][243] ;
wire   [4:0] \A[0][244] ;
wire   [4:0] \A[0][245] ;
wire   [4:0] \A[0][246] ;
wire   [4:0] \A[0][247] ;
wire   [4:0] \A[0][248] ;
wire   [4:0] \A[0][249] ;
wire   [4:0] \A[0][250] ;
wire   [4:0] \A[0][251] ;
wire   [4:0] \A[0][252] ;
wire   [4:0] \A[0][253] ;
wire   [4:0] \A[0][254] ;
wire   [4:0] \A[0][255] ;
wire   [4:0] \A[1][0] ;
wire   [4:0] \A[1][1] ;
wire   [4:0] \A[1][2] ;
wire   [4:0] \A[1][3] ;
wire   [4:0] \A[1][4] ;
wire   [4:0] \A[1][5] ;
wire   [4:0] \A[1][6] ;
wire   [4:0] \A[1][7] ;
wire   [4:0] \A[1][8] ;
wire   [4:0] \A[1][9] ;
wire   [4:0] \A[1][10] ;
wire   [4:0] \A[1][11] ;
wire   [4:0] \A[1][12] ;
wire   [4:0] \A[1][13] ;
wire   [4:0] \A[1][14] ;
wire   [4:0] \A[1][15] ;
wire   [4:0] \A[1][16] ;
wire   [4:0] \A[1][17] ;
wire   [4:0] \A[1][18] ;
wire   [4:0] \A[1][19] ;
wire   [4:0] \A[1][20] ;
wire   [4:0] \A[1][21] ;
wire   [4:0] \A[1][22] ;
wire   [4:0] \A[1][23] ;
wire   [4:0] \A[1][24] ;
wire   [4:0] \A[1][25] ;
wire   [4:0] \A[1][26] ;
wire   [4:0] \A[1][27] ;
wire   [4:0] \A[1][28] ;
wire   [4:0] \A[1][29] ;
wire   [4:0] \A[1][30] ;
wire   [4:0] \A[1][31] ;
wire   [4:0] \A[1][32] ;
wire   [4:0] \A[1][33] ;
wire   [4:0] \A[1][34] ;
wire   [4:0] \A[1][35] ;
wire   [4:0] \A[1][36] ;
wire   [4:0] \A[1][37] ;
wire   [4:0] \A[1][38] ;
wire   [4:0] \A[1][39] ;
wire   [4:0] \A[1][40] ;
wire   [4:0] \A[1][41] ;
wire   [4:0] \A[1][42] ;
wire   [4:0] \A[1][43] ;
wire   [4:0] \A[1][44] ;
wire   [4:0] \A[1][45] ;
wire   [4:0] \A[1][46] ;
wire   [4:0] \A[1][47] ;
wire   [4:0] \A[1][48] ;
wire   [4:0] \A[1][49] ;
wire   [4:0] \A[1][50] ;
wire   [4:0] \A[1][51] ;
wire   [4:0] \A[1][52] ;
wire   [4:0] \A[1][53] ;
wire   [4:0] \A[1][54] ;
wire   [4:0] \A[1][55] ;
wire   [4:0] \A[1][56] ;
wire   [4:0] \A[1][57] ;
wire   [4:0] \A[1][58] ;
wire   [4:0] \A[1][59] ;
wire   [4:0] \A[1][60] ;
wire   [4:0] \A[1][61] ;
wire   [4:0] \A[1][62] ;
wire   [4:0] \A[1][63] ;
wire   [4:0] \A[1][64] ;
wire   [4:0] \A[1][65] ;
wire   [4:0] \A[1][66] ;
wire   [4:0] \A[1][67] ;
wire   [4:0] \A[1][68] ;
wire   [4:0] \A[1][69] ;
wire   [4:0] \A[1][70] ;
wire   [4:0] \A[1][71] ;
wire   [4:0] \A[1][72] ;
wire   [4:0] \A[1][73] ;
wire   [4:0] \A[1][74] ;
wire   [4:0] \A[1][75] ;
wire   [4:0] \A[1][76] ;
wire   [4:0] \A[1][77] ;
wire   [4:0] \A[1][78] ;
wire   [4:0] \A[1][79] ;
wire   [4:0] \A[1][80] ;
wire   [4:0] \A[1][81] ;
wire   [4:0] \A[1][82] ;
wire   [4:0] \A[1][83] ;
wire   [4:0] \A[1][84] ;
wire   [4:0] \A[1][85] ;
wire   [4:0] \A[1][86] ;
wire   [4:0] \A[1][87] ;
wire   [4:0] \A[1][88] ;
wire   [4:0] \A[1][89] ;
wire   [4:0] \A[1][90] ;
wire   [4:0] \A[1][91] ;
wire   [4:0] \A[1][92] ;
wire   [4:0] \A[1][93] ;
wire   [4:0] \A[1][94] ;
wire   [4:0] \A[1][95] ;
wire   [4:0] \A[1][96] ;
wire   [4:0] \A[1][97] ;
wire   [4:0] \A[1][98] ;
wire   [4:0] \A[1][99] ;
wire   [4:0] \A[1][100] ;
wire   [4:0] \A[1][101] ;
wire   [4:0] \A[1][102] ;
wire   [4:0] \A[1][103] ;
wire   [4:0] \A[1][104] ;
wire   [4:0] \A[1][105] ;
wire   [4:0] \A[1][106] ;
wire   [4:0] \A[1][107] ;
wire   [4:0] \A[1][108] ;
wire   [4:0] \A[1][109] ;
wire   [4:0] \A[1][110] ;
wire   [4:0] \A[1][111] ;
wire   [4:0] \A[1][112] ;
wire   [4:0] \A[1][113] ;
wire   [4:0] \A[1][114] ;
wire   [4:0] \A[1][115] ;
wire   [4:0] \A[1][116] ;
wire   [4:0] \A[1][117] ;
wire   [4:0] \A[1][118] ;
wire   [4:0] \A[1][119] ;
wire   [4:0] \A[1][120] ;
wire   [4:0] \A[1][121] ;
wire   [4:0] \A[1][122] ;
wire   [4:0] \A[1][123] ;
wire   [4:0] \A[1][124] ;
wire   [4:0] \A[1][125] ;
wire   [4:0] \A[1][126] ;
wire   [4:0] \A[1][127] ;
wire   [4:0] \A[1][128] ;
wire   [4:0] \A[1][129] ;
wire   [4:0] \A[1][130] ;
wire   [4:0] \A[1][131] ;
wire   [4:0] \A[1][132] ;
wire   [4:0] \A[1][133] ;
wire   [4:0] \A[1][134] ;
wire   [4:0] \A[1][135] ;
wire   [4:0] \A[1][136] ;
wire   [4:0] \A[1][137] ;
wire   [4:0] \A[1][138] ;
wire   [4:0] \A[1][139] ;
wire   [4:0] \A[1][140] ;
wire   [4:0] \A[1][141] ;
wire   [4:0] \A[1][142] ;
wire   [4:0] \A[1][143] ;
wire   [4:0] \A[1][144] ;
wire   [4:0] \A[1][145] ;
wire   [4:0] \A[1][146] ;
wire   [4:0] \A[1][147] ;
wire   [4:0] \A[1][148] ;
wire   [4:0] \A[1][149] ;
wire   [4:0] \A[1][150] ;
wire   [4:0] \A[1][151] ;
wire   [4:0] \A[1][152] ;
wire   [4:0] \A[1][153] ;
wire   [4:0] \A[1][154] ;
wire   [4:0] \A[1][155] ;
wire   [4:0] \A[1][156] ;
wire   [4:0] \A[1][157] ;
wire   [4:0] \A[1][158] ;
wire   [4:0] \A[1][159] ;
wire   [4:0] \A[1][160] ;
wire   [4:0] \A[1][161] ;
wire   [4:0] \A[1][162] ;
wire   [4:0] \A[1][163] ;
wire   [4:0] \A[1][164] ;
wire   [4:0] \A[1][165] ;
wire   [4:0] \A[1][166] ;
wire   [4:0] \A[1][167] ;
wire   [4:0] \A[1][168] ;
wire   [4:0] \A[1][169] ;
wire   [4:0] \A[1][170] ;
wire   [4:0] \A[1][171] ;
wire   [4:0] \A[1][172] ;
wire   [4:0] \A[1][173] ;
wire   [4:0] \A[1][174] ;
wire   [4:0] \A[1][175] ;
wire   [4:0] \A[1][176] ;
wire   [4:0] \A[1][177] ;
wire   [4:0] \A[1][178] ;
wire   [4:0] \A[1][179] ;
wire   [4:0] \A[1][180] ;
wire   [4:0] \A[1][181] ;
wire   [4:0] \A[1][182] ;
wire   [4:0] \A[1][183] ;
wire   [4:0] \A[1][184] ;
wire   [4:0] \A[1][185] ;
wire   [4:0] \A[1][186] ;
wire   [4:0] \A[1][187] ;
wire   [4:0] \A[1][188] ;
wire   [4:0] \A[1][189] ;
wire   [4:0] \A[1][190] ;
wire   [4:0] \A[1][191] ;
wire   [4:0] \A[1][192] ;
wire   [4:0] \A[1][193] ;
wire   [4:0] \A[1][194] ;
wire   [4:0] \A[1][195] ;
wire   [4:0] \A[1][196] ;
wire   [4:0] \A[1][197] ;
wire   [4:0] \A[1][198] ;
wire   [4:0] \A[1][199] ;
wire   [4:0] \A[1][200] ;
wire   [4:0] \A[1][201] ;
wire   [4:0] \A[1][202] ;
wire   [4:0] \A[1][203] ;
wire   [4:0] \A[1][204] ;
wire   [4:0] \A[1][205] ;
wire   [4:0] \A[1][206] ;
wire   [4:0] \A[1][207] ;
wire   [4:0] \A[1][208] ;
wire   [4:0] \A[1][209] ;
wire   [4:0] \A[1][210] ;
wire   [4:0] \A[1][211] ;
wire   [4:0] \A[1][212] ;
wire   [4:0] \A[1][213] ;
wire   [4:0] \A[1][214] ;
wire   [4:0] \A[1][215] ;
wire   [4:0] \A[1][216] ;
wire   [4:0] \A[1][217] ;
wire   [4:0] \A[1][218] ;
wire   [4:0] \A[1][219] ;
wire   [4:0] \A[1][220] ;
wire   [4:0] \A[1][221] ;
wire   [4:0] \A[1][222] ;
wire   [4:0] \A[1][223] ;
wire   [4:0] \A[1][224] ;
wire   [4:0] \A[1][225] ;
wire   [4:0] \A[1][226] ;
wire   [4:0] \A[1][227] ;
wire   [4:0] \A[1][228] ;
wire   [4:0] \A[1][229] ;
wire   [4:0] \A[1][230] ;
wire   [4:0] \A[1][231] ;
wire   [4:0] \A[1][232] ;
wire   [4:0] \A[1][233] ;
wire   [4:0] \A[1][234] ;
wire   [4:0] \A[1][235] ;
wire   [4:0] \A[1][236] ;
wire   [4:0] \A[1][237] ;
wire   [4:0] \A[1][238] ;
wire   [4:0] \A[1][239] ;
wire   [4:0] \A[1][240] ;
wire   [4:0] \A[1][241] ;
wire   [4:0] \A[1][242] ;
wire   [4:0] \A[1][243] ;
wire   [4:0] \A[1][244] ;
wire   [4:0] \A[1][245] ;
wire   [4:0] \A[1][246] ;
wire   [4:0] \A[1][247] ;
wire   [4:0] \A[1][248] ;
wire   [4:0] \A[1][249] ;
wire   [4:0] \A[1][250] ;
wire   [4:0] \A[1][251] ;
wire   [4:0] \A[1][252] ;
wire   [4:0] \A[1][253] ;
wire   [4:0] \A[1][254] ;
wire   [4:0] \A[1][255] ;
wire   [4:0] \A[2][0] ;
wire   [4:0] \A[2][1] ;
wire   [4:0] \A[2][2] ;
wire   [4:0] \A[2][3] ;
wire   [4:0] \A[2][4] ;
wire   [4:0] \A[2][5] ;
wire   [4:0] \A[2][6] ;
wire   [4:0] \A[2][7] ;
wire   [4:0] \A[2][8] ;
wire   [4:0] \A[2][9] ;
wire   [4:0] \A[2][10] ;
wire   [4:0] \A[2][11] ;
wire   [4:0] \A[2][12] ;
wire   [4:0] \A[2][13] ;
wire   [4:0] \A[2][14] ;
wire   [4:0] \A[2][15] ;
wire   [4:0] \A[2][16] ;
wire   [4:0] \A[2][17] ;
wire   [4:0] \A[2][18] ;
wire   [4:0] \A[2][19] ;
wire   [4:0] \A[2][20] ;
wire   [4:0] \A[2][21] ;
wire   [4:0] \A[2][22] ;
wire   [4:0] \A[2][23] ;
wire   [4:0] \A[2][24] ;
wire   [4:0] \A[2][25] ;
wire   [4:0] \A[2][26] ;
wire   [4:0] \A[2][27] ;
wire   [4:0] \A[2][28] ;
wire   [4:0] \A[2][29] ;
wire   [4:0] \A[2][30] ;
wire   [4:0] \A[2][31] ;
wire   [4:0] \A[2][32] ;
wire   [4:0] \A[2][33] ;
wire   [4:0] \A[2][34] ;
wire   [4:0] \A[2][35] ;
wire   [4:0] \A[2][36] ;
wire   [4:0] \A[2][37] ;
wire   [4:0] \A[2][38] ;
wire   [4:0] \A[2][39] ;
wire   [4:0] \A[2][40] ;
wire   [4:0] \A[2][41] ;
wire   [4:0] \A[2][42] ;
wire   [4:0] \A[2][43] ;
wire   [4:0] \A[2][44] ;
wire   [4:0] \A[2][45] ;
wire   [4:0] \A[2][46] ;
wire   [4:0] \A[2][47] ;
wire   [4:0] \A[2][48] ;
wire   [4:0] \A[2][49] ;
wire   [4:0] \A[2][50] ;
wire   [4:0] \A[2][51] ;
wire   [4:0] \A[2][52] ;
wire   [4:0] \A[2][53] ;
wire   [4:0] \A[2][54] ;
wire   [4:0] \A[2][55] ;
wire   [4:0] \A[2][56] ;
wire   [4:0] \A[2][57] ;
wire   [4:0] \A[2][58] ;
wire   [4:0] \A[2][59] ;
wire   [4:0] \A[2][60] ;
wire   [4:0] \A[2][61] ;
wire   [4:0] \A[2][62] ;
wire   [4:0] \A[2][63] ;
wire   [4:0] \A[2][64] ;
wire   [4:0] \A[2][65] ;
wire   [4:0] \A[2][66] ;
wire   [4:0] \A[2][67] ;
wire   [4:0] \A[2][68] ;
wire   [4:0] \A[2][69] ;
wire   [4:0] \A[2][70] ;
wire   [4:0] \A[2][71] ;
wire   [4:0] \A[2][72] ;
wire   [4:0] \A[2][73] ;
wire   [4:0] \A[2][74] ;
wire   [4:0] \A[2][75] ;
wire   [4:0] \A[2][76] ;
wire   [4:0] \A[2][77] ;
wire   [4:0] \A[2][78] ;
wire   [4:0] \A[2][79] ;
wire   [4:0] \A[2][80] ;
wire   [4:0] \A[2][81] ;
wire   [4:0] \A[2][82] ;
wire   [4:0] \A[2][83] ;
wire   [4:0] \A[2][84] ;
wire   [4:0] \A[2][85] ;
wire   [4:0] \A[2][86] ;
wire   [4:0] \A[2][87] ;
wire   [4:0] \A[2][88] ;
wire   [4:0] \A[2][89] ;
wire   [4:0] \A[2][90] ;
wire   [4:0] \A[2][91] ;
wire   [4:0] \A[2][92] ;
wire   [4:0] \A[2][93] ;
wire   [4:0] \A[2][94] ;
wire   [4:0] \A[2][95] ;
wire   [4:0] \A[2][96] ;
wire   [4:0] \A[2][97] ;
wire   [4:0] \A[2][98] ;
wire   [4:0] \A[2][99] ;
wire   [4:0] \A[2][100] ;
wire   [4:0] \A[2][101] ;
wire   [4:0] \A[2][102] ;
wire   [4:0] \A[2][103] ;
wire   [4:0] \A[2][104] ;
wire   [4:0] \A[2][105] ;
wire   [4:0] \A[2][106] ;
wire   [4:0] \A[2][107] ;
wire   [4:0] \A[2][108] ;
wire   [4:0] \A[2][109] ;
wire   [4:0] \A[2][110] ;
wire   [4:0] \A[2][111] ;
wire   [4:0] \A[2][112] ;
wire   [4:0] \A[2][113] ;
wire   [4:0] \A[2][114] ;
wire   [4:0] \A[2][115] ;
wire   [4:0] \A[2][116] ;
wire   [4:0] \A[2][117] ;
wire   [4:0] \A[2][118] ;
wire   [4:0] \A[2][119] ;
wire   [4:0] \A[2][120] ;
wire   [4:0] \A[2][121] ;
wire   [4:0] \A[2][122] ;
wire   [4:0] \A[2][123] ;
wire   [4:0] \A[2][124] ;
wire   [4:0] \A[2][125] ;
wire   [4:0] \A[2][126] ;
wire   [4:0] \A[2][127] ;
wire   [4:0] \A[2][128] ;
wire   [4:0] \A[2][129] ;
wire   [4:0] \A[2][130] ;
wire   [4:0] \A[2][131] ;
wire   [4:0] \A[2][132] ;
wire   [4:0] \A[2][133] ;
wire   [4:0] \A[2][134] ;
wire   [4:0] \A[2][135] ;
wire   [4:0] \A[2][136] ;
wire   [4:0] \A[2][137] ;
wire   [4:0] \A[2][138] ;
wire   [4:0] \A[2][139] ;
wire   [4:0] \A[2][140] ;
wire   [4:0] \A[2][141] ;
wire   [4:0] \A[2][142] ;
wire   [4:0] \A[2][143] ;
wire   [4:0] \A[2][144] ;
wire   [4:0] \A[2][145] ;
wire   [4:0] \A[2][146] ;
wire   [4:0] \A[2][147] ;
wire   [4:0] \A[2][148] ;
wire   [4:0] \A[2][149] ;
wire   [4:0] \A[2][150] ;
wire   [4:0] \A[2][151] ;
wire   [4:0] \A[2][152] ;
wire   [4:0] \A[2][153] ;
wire   [4:0] \A[2][154] ;
wire   [4:0] \A[2][155] ;
wire   [4:0] \A[2][156] ;
wire   [4:0] \A[2][157] ;
wire   [4:0] \A[2][158] ;
wire   [4:0] \A[2][159] ;
wire   [4:0] \A[2][160] ;
wire   [4:0] \A[2][161] ;
wire   [4:0] \A[2][162] ;
wire   [4:0] \A[2][163] ;
wire   [4:0] \A[2][164] ;
wire   [4:0] \A[2][165] ;
wire   [4:0] \A[2][166] ;
wire   [4:0] \A[2][167] ;
wire   [4:0] \A[2][168] ;
wire   [4:0] \A[2][169] ;
wire   [4:0] \A[2][170] ;
wire   [4:0] \A[2][171] ;
wire   [4:0] \A[2][172] ;
wire   [4:0] \A[2][173] ;
wire   [4:0] \A[2][174] ;
wire   [4:0] \A[2][175] ;
wire   [4:0] \A[2][176] ;
wire   [4:0] \A[2][177] ;
wire   [4:0] \A[2][178] ;
wire   [4:0] \A[2][179] ;
wire   [4:0] \A[2][180] ;
wire   [4:0] \A[2][181] ;
wire   [4:0] \A[2][182] ;
wire   [4:0] \A[2][183] ;
wire   [4:0] \A[2][184] ;
wire   [4:0] \A[2][185] ;
wire   [4:0] \A[2][186] ;
wire   [4:0] \A[2][187] ;
wire   [4:0] \A[2][188] ;
wire   [4:0] \A[2][189] ;
wire   [4:0] \A[2][190] ;
wire   [4:0] \A[2][191] ;
wire   [4:0] \A[2][192] ;
wire   [4:0] \A[2][193] ;
wire   [4:0] \A[2][194] ;
wire   [4:0] \A[2][195] ;
wire   [4:0] \A[2][196] ;
wire   [4:0] \A[2][197] ;
wire   [4:0] \A[2][198] ;
wire   [4:0] \A[2][199] ;
wire   [4:0] \A[2][200] ;
wire   [4:0] \A[2][201] ;
wire   [4:0] \A[2][202] ;
wire   [4:0] \A[2][203] ;
wire   [4:0] \A[2][204] ;
wire   [4:0] \A[2][205] ;
wire   [4:0] \A[2][206] ;
wire   [4:0] \A[2][207] ;
wire   [4:0] \A[2][208] ;
wire   [4:0] \A[2][209] ;
wire   [4:0] \A[2][210] ;
wire   [4:0] \A[2][211] ;
wire   [4:0] \A[2][212] ;
wire   [4:0] \A[2][213] ;
wire   [4:0] \A[2][214] ;
wire   [4:0] \A[2][215] ;
wire   [4:0] \A[2][216] ;
wire   [4:0] \A[2][217] ;
wire   [4:0] \A[2][218] ;
wire   [4:0] \A[2][219] ;
wire   [4:0] \A[2][220] ;
wire   [4:0] \A[2][221] ;
wire   [4:0] \A[2][222] ;
wire   [4:0] \A[2][223] ;
wire   [4:0] \A[2][224] ;
wire   [4:0] \A[2][225] ;
wire   [4:0] \A[2][226] ;
wire   [4:0] \A[2][227] ;
wire   [4:0] \A[2][228] ;
wire   [4:0] \A[2][229] ;
wire   [4:0] \A[2][230] ;
wire   [4:0] \A[2][231] ;
wire   [4:0] \A[2][232] ;
wire   [4:0] \A[2][233] ;
wire   [4:0] \A[2][234] ;
wire   [4:0] \A[2][235] ;
wire   [4:0] \A[2][236] ;
wire   [4:0] \A[2][237] ;
wire   [4:0] \A[2][238] ;
wire   [4:0] \A[2][239] ;
wire   [4:0] \A[2][240] ;
wire   [4:0] \A[2][241] ;
wire   [4:0] \A[2][242] ;
wire   [4:0] \A[2][243] ;
wire   [4:0] \A[2][244] ;
wire   [4:0] \A[2][245] ;
wire   [4:0] \A[2][246] ;
wire   [4:0] \A[2][247] ;
wire   [4:0] \A[2][248] ;
wire   [4:0] \A[2][249] ;
wire   [4:0] \A[2][250] ;
wire   [4:0] \A[2][251] ;
wire   [4:0] \A[2][252] ;
wire   [4:0] \A[2][253] ;
wire   [4:0] \A[2][254] ;
wire   [4:0] \A[2][255] ;
wire   [4:0] \A[3][0] ;
wire   [4:0] \A[3][1] ;
wire   [4:0] \A[3][2] ;
wire   [4:0] \A[3][3] ;
wire   [4:0] \A[3][4] ;
wire   [4:0] \A[3][5] ;
wire   [4:0] \A[3][6] ;
wire   [4:0] \A[3][7] ;
wire   [4:0] \A[3][8] ;
wire   [4:0] \A[3][9] ;
wire   [4:0] \A[3][10] ;
wire   [4:0] \A[3][11] ;
wire   [4:0] \A[3][12] ;
wire   [4:0] \A[3][13] ;
wire   [4:0] \A[3][14] ;
wire   [4:0] \A[3][15] ;
wire   [4:0] \A[3][16] ;
wire   [4:0] \A[3][17] ;
wire   [4:0] \A[3][18] ;
wire   [4:0] \A[3][19] ;
wire   [4:0] \A[3][20] ;
wire   [4:0] \A[3][21] ;
wire   [4:0] \A[3][22] ;
wire   [4:0] \A[3][23] ;
wire   [4:0] \A[3][24] ;
wire   [4:0] \A[3][25] ;
wire   [4:0] \A[3][26] ;
wire   [4:0] \A[3][27] ;
wire   [4:0] \A[3][28] ;
wire   [4:0] \A[3][29] ;
wire   [4:0] \A[3][30] ;
wire   [4:0] \A[3][31] ;
wire   [4:0] \A[3][32] ;
wire   [4:0] \A[3][33] ;
wire   [4:0] \A[3][34] ;
wire   [4:0] \A[3][35] ;
wire   [4:0] \A[3][36] ;
wire   [4:0] \A[3][37] ;
wire   [4:0] \A[3][38] ;
wire   [4:0] \A[3][39] ;
wire   [4:0] \A[3][40] ;
wire   [4:0] \A[3][41] ;
wire   [4:0] \A[3][42] ;
wire   [4:0] \A[3][43] ;
wire   [4:0] \A[3][44] ;
wire   [4:0] \A[3][45] ;
wire   [4:0] \A[3][46] ;
wire   [4:0] \A[3][47] ;
wire   [4:0] \A[3][48] ;
wire   [4:0] \A[3][49] ;
wire   [4:0] \A[3][50] ;
wire   [4:0] \A[3][51] ;
wire   [4:0] \A[3][52] ;
wire   [4:0] \A[3][53] ;
wire   [4:0] \A[3][54] ;
wire   [4:0] \A[3][55] ;
wire   [4:0] \A[3][56] ;
wire   [4:0] \A[3][57] ;
wire   [4:0] \A[3][58] ;
wire   [4:0] \A[3][59] ;
wire   [4:0] \A[3][60] ;
wire   [4:0] \A[3][61] ;
wire   [4:0] \A[3][62] ;
wire   [4:0] \A[3][63] ;
wire   [4:0] \A[3][64] ;
wire   [4:0] \A[3][65] ;
wire   [4:0] \A[3][66] ;
wire   [4:0] \A[3][67] ;
wire   [4:0] \A[3][68] ;
wire   [4:0] \A[3][69] ;
wire   [4:0] \A[3][70] ;
wire   [4:0] \A[3][71] ;
wire   [4:0] \A[3][72] ;
wire   [4:0] \A[3][73] ;
wire   [4:0] \A[3][74] ;
wire   [4:0] \A[3][75] ;
wire   [4:0] \A[3][76] ;
wire   [4:0] \A[3][77] ;
wire   [4:0] \A[3][78] ;
wire   [4:0] \A[3][79] ;
wire   [4:0] \A[3][80] ;
wire   [4:0] \A[3][81] ;
wire   [4:0] \A[3][82] ;
wire   [4:0] \A[3][83] ;
wire   [4:0] \A[3][84] ;
wire   [4:0] \A[3][85] ;
wire   [4:0] \A[3][86] ;
wire   [4:0] \A[3][87] ;
wire   [4:0] \A[3][88] ;
wire   [4:0] \A[3][89] ;
wire   [4:0] \A[3][90] ;
wire   [4:0] \A[3][91] ;
wire   [4:0] \A[3][92] ;
wire   [4:0] \A[3][93] ;
wire   [4:0] \A[3][94] ;
wire   [4:0] \A[3][95] ;
wire   [4:0] \A[3][96] ;
wire   [4:0] \A[3][97] ;
wire   [4:0] \A[3][98] ;
wire   [4:0] \A[3][99] ;
wire   [4:0] \A[3][100] ;
wire   [4:0] \A[3][101] ;
wire   [4:0] \A[3][102] ;
wire   [4:0] \A[3][103] ;
wire   [4:0] \A[3][104] ;
wire   [4:0] \A[3][105] ;
wire   [4:0] \A[3][106] ;
wire   [4:0] \A[3][107] ;
wire   [4:0] \A[3][108] ;
wire   [4:0] \A[3][109] ;
wire   [4:0] \A[3][110] ;
wire   [4:0] \A[3][111] ;
wire   [4:0] \A[3][112] ;
wire   [4:0] \A[3][113] ;
wire   [4:0] \A[3][114] ;
wire   [4:0] \A[3][115] ;
wire   [4:0] \A[3][116] ;
wire   [4:0] \A[3][117] ;
wire   [4:0] \A[3][118] ;
wire   [4:0] \A[3][119] ;
wire   [4:0] \A[3][120] ;
wire   [4:0] \A[3][121] ;
wire   [4:0] \A[3][122] ;
wire   [4:0] \A[3][123] ;
wire   [4:0] \A[3][124] ;
wire   [4:0] \A[3][125] ;
wire   [4:0] \A[3][126] ;
wire   [4:0] \A[3][127] ;
wire   [4:0] \A[3][128] ;
wire   [4:0] \A[3][129] ;
wire   [4:0] \A[3][130] ;
wire   [4:0] \A[3][131] ;
wire   [4:0] \A[3][132] ;
wire   [4:0] \A[3][133] ;
wire   [4:0] \A[3][134] ;
wire   [4:0] \A[3][135] ;
wire   [4:0] \A[3][136] ;
wire   [4:0] \A[3][137] ;
wire   [4:0] \A[3][138] ;
wire   [4:0] \A[3][139] ;
wire   [4:0] \A[3][140] ;
wire   [4:0] \A[3][141] ;
wire   [4:0] \A[3][142] ;
wire   [4:0] \A[3][143] ;
wire   [4:0] \A[3][144] ;
wire   [4:0] \A[3][145] ;
wire   [4:0] \A[3][146] ;
wire   [4:0] \A[3][147] ;
wire   [4:0] \A[3][148] ;
wire   [4:0] \A[3][149] ;
wire   [4:0] \A[3][150] ;
wire   [4:0] \A[3][151] ;
wire   [4:0] \A[3][152] ;
wire   [4:0] \A[3][153] ;
wire   [4:0] \A[3][154] ;
wire   [4:0] \A[3][155] ;
wire   [4:0] \A[3][156] ;
wire   [4:0] \A[3][157] ;
wire   [4:0] \A[3][158] ;
wire   [4:0] \A[3][159] ;
wire   [4:0] \A[3][160] ;
wire   [4:0] \A[3][161] ;
wire   [4:0] \A[3][162] ;
wire   [4:0] \A[3][163] ;
wire   [4:0] \A[3][164] ;
wire   [4:0] \A[3][165] ;
wire   [4:0] \A[3][166] ;
wire   [4:0] \A[3][167] ;
wire   [4:0] \A[3][168] ;
wire   [4:0] \A[3][169] ;
wire   [4:0] \A[3][170] ;
wire   [4:0] \A[3][171] ;
wire   [4:0] \A[3][172] ;
wire   [4:0] \A[3][173] ;
wire   [4:0] \A[3][174] ;
wire   [4:0] \A[3][175] ;
wire   [4:0] \A[3][176] ;
wire   [4:0] \A[3][177] ;
wire   [4:0] \A[3][178] ;
wire   [4:0] \A[3][179] ;
wire   [4:0] \A[3][180] ;
wire   [4:0] \A[3][181] ;
wire   [4:0] \A[3][182] ;
wire   [4:0] \A[3][183] ;
wire   [4:0] \A[3][184] ;
wire   [4:0] \A[3][185] ;
wire   [4:0] \A[3][186] ;
wire   [4:0] \A[3][187] ;
wire   [4:0] \A[3][188] ;
wire   [4:0] \A[3][189] ;
wire   [4:0] \A[3][190] ;
wire   [4:0] \A[3][191] ;
wire   [4:0] \A[3][192] ;
wire   [4:0] \A[3][193] ;
wire   [4:0] \A[3][194] ;
wire   [4:0] \A[3][195] ;
wire   [4:0] \A[3][196] ;
wire   [4:0] \A[3][197] ;
wire   [4:0] \A[3][198] ;
wire   [4:0] \A[3][199] ;
wire   [4:0] \A[3][200] ;
wire   [4:0] \A[3][201] ;
wire   [4:0] \A[3][202] ;
wire   [4:0] \A[3][203] ;
wire   [4:0] \A[3][204] ;
wire   [4:0] \A[3][205] ;
wire   [4:0] \A[3][206] ;
wire   [4:0] \A[3][207] ;
wire   [4:0] \A[3][208] ;
wire   [4:0] \A[3][209] ;
wire   [4:0] \A[3][210] ;
wire   [4:0] \A[3][211] ;
wire   [4:0] \A[3][212] ;
wire   [4:0] \A[3][213] ;
wire   [4:0] \A[3][214] ;
wire   [4:0] \A[3][215] ;
wire   [4:0] \A[3][216] ;
wire   [4:0] \A[3][217] ;
wire   [4:0] \A[3][218] ;
wire   [4:0] \A[3][219] ;
wire   [4:0] \A[3][220] ;
wire   [4:0] \A[3][221] ;
wire   [4:0] \A[3][222] ;
wire   [4:0] \A[3][223] ;
wire   [4:0] \A[3][224] ;
wire   [4:0] \A[3][225] ;
wire   [4:0] \A[3][226] ;
wire   [4:0] \A[3][227] ;
wire   [4:0] \A[3][228] ;
wire   [4:0] \A[3][229] ;
wire   [4:0] \A[3][230] ;
wire   [4:0] \A[3][231] ;
wire   [4:0] \A[3][232] ;
wire   [4:0] \A[3][233] ;
wire   [4:0] \A[3][234] ;
wire   [4:0] \A[3][235] ;
wire   [4:0] \A[3][236] ;
wire   [4:0] \A[3][237] ;
wire   [4:0] \A[3][238] ;
wire   [4:0] \A[3][239] ;
wire   [4:0] \A[3][240] ;
wire   [4:0] \A[3][241] ;
wire   [4:0] \A[3][242] ;
wire   [4:0] \A[3][243] ;
wire   [4:0] \A[3][244] ;
wire   [4:0] \A[3][245] ;
wire   [4:0] \A[3][246] ;
wire   [4:0] \A[3][247] ;
wire   [4:0] \A[3][248] ;
wire   [4:0] \A[3][249] ;
wire   [4:0] \A[3][250] ;
wire   [4:0] \A[3][251] ;
wire   [4:0] \A[3][252] ;
wire   [4:0] \A[3][253] ;
wire   [4:0] \A[3][254] ;
wire   [4:0] \A[3][255] ;
wire   [4:0] \A[4][0] ;
wire   [4:0] \A[4][1] ;
wire   [4:0] \A[4][2] ;
wire   [4:0] \A[4][3] ;
wire   [4:0] \A[4][4] ;
wire   [4:0] \A[4][5] ;
wire   [4:0] \A[4][6] ;
wire   [4:0] \A[4][7] ;
wire   [4:0] \A[4][8] ;
wire   [4:0] \A[4][9] ;
wire   [4:0] \A[4][10] ;
wire   [4:0] \A[4][11] ;
wire   [4:0] \A[4][12] ;
wire   [4:0] \A[4][13] ;
wire   [4:0] \A[4][14] ;
wire   [4:0] \A[4][15] ;
wire   [4:0] \A[4][16] ;
wire   [4:0] \A[4][17] ;
wire   [4:0] \A[4][18] ;
wire   [4:0] \A[4][19] ;
wire   [4:0] \A[4][20] ;
wire   [4:0] \A[4][21] ;
wire   [4:0] \A[4][22] ;
wire   [4:0] \A[4][23] ;
wire   [4:0] \A[4][24] ;
wire   [4:0] \A[4][25] ;
wire   [4:0] \A[4][26] ;
wire   [4:0] \A[4][27] ;
wire   [4:0] \A[4][28] ;
wire   [4:0] \A[4][29] ;
wire   [4:0] \A[4][30] ;
wire   [4:0] \A[4][31] ;
wire   [4:0] \A[4][32] ;
wire   [4:0] \A[4][33] ;
wire   [4:0] \A[4][34] ;
wire   [4:0] \A[4][35] ;
wire   [4:0] \A[4][36] ;
wire   [4:0] \A[4][37] ;
wire   [4:0] \A[4][38] ;
wire   [4:0] \A[4][39] ;
wire   [4:0] \A[4][40] ;
wire   [4:0] \A[4][41] ;
wire   [4:0] \A[4][42] ;
wire   [4:0] \A[4][43] ;
wire   [4:0] \A[4][44] ;
wire   [4:0] \A[4][45] ;
wire   [4:0] \A[4][46] ;
wire   [4:0] \A[4][47] ;
wire   [4:0] \A[4][48] ;
wire   [4:0] \A[4][49] ;
wire   [4:0] \A[4][50] ;
wire   [4:0] \A[4][51] ;
wire   [4:0] \A[4][52] ;
wire   [4:0] \A[4][53] ;
wire   [4:0] \A[4][54] ;
wire   [4:0] \A[4][55] ;
wire   [4:0] \A[4][56] ;
wire   [4:0] \A[4][57] ;
wire   [4:0] \A[4][58] ;
wire   [4:0] \A[4][59] ;
wire   [4:0] \A[4][60] ;
wire   [4:0] \A[4][61] ;
wire   [4:0] \A[4][62] ;
wire   [4:0] \A[4][63] ;
wire   [4:0] \A[4][64] ;
wire   [4:0] \A[4][65] ;
wire   [4:0] \A[4][66] ;
wire   [4:0] \A[4][67] ;
wire   [4:0] \A[4][68] ;
wire   [4:0] \A[4][69] ;
wire   [4:0] \A[4][70] ;
wire   [4:0] \A[4][71] ;
wire   [4:0] \A[4][72] ;
wire   [4:0] \A[4][73] ;
wire   [4:0] \A[4][74] ;
wire   [4:0] \A[4][75] ;
wire   [4:0] \A[4][76] ;
wire   [4:0] \A[4][77] ;
wire   [4:0] \A[4][78] ;
wire   [4:0] \A[4][79] ;
wire   [4:0] \A[4][80] ;
wire   [4:0] \A[4][81] ;
wire   [4:0] \A[4][82] ;
wire   [4:0] \A[4][83] ;
wire   [4:0] \A[4][84] ;
wire   [4:0] \A[4][85] ;
wire   [4:0] \A[4][86] ;
wire   [4:0] \A[4][87] ;
wire   [4:0] \A[4][88] ;
wire   [4:0] \A[4][89] ;
wire   [4:0] \A[4][90] ;
wire   [4:0] \A[4][91] ;
wire   [4:0] \A[4][92] ;
wire   [4:0] \A[4][93] ;
wire   [4:0] \A[4][94] ;
wire   [4:0] \A[4][95] ;
wire   [4:0] \A[4][96] ;
wire   [4:0] \A[4][97] ;
wire   [4:0] \A[4][98] ;
wire   [4:0] \A[4][99] ;
wire   [4:0] \A[4][100] ;
wire   [4:0] \A[4][101] ;
wire   [4:0] \A[4][102] ;
wire   [4:0] \A[4][103] ;
wire   [4:0] \A[4][104] ;
wire   [4:0] \A[4][105] ;
wire   [4:0] \A[4][106] ;
wire   [4:0] \A[4][107] ;
wire   [4:0] \A[4][108] ;
wire   [4:0] \A[4][109] ;
wire   [4:0] \A[4][110] ;
wire   [4:0] \A[4][111] ;
wire   [4:0] \A[4][112] ;
wire   [4:0] \A[4][113] ;
wire   [4:0] \A[4][114] ;
wire   [4:0] \A[4][115] ;
wire   [4:0] \A[4][116] ;
wire   [4:0] \A[4][117] ;
wire   [4:0] \A[4][118] ;
wire   [4:0] \A[4][119] ;
wire   [4:0] \A[4][120] ;
wire   [4:0] \A[4][121] ;
wire   [4:0] \A[4][122] ;
wire   [4:0] \A[4][123] ;
wire   [4:0] \A[4][124] ;
wire   [4:0] \A[4][125] ;
wire   [4:0] \A[4][126] ;
wire   [4:0] \A[4][127] ;
wire   [4:0] \A[4][128] ;
wire   [4:0] \A[4][129] ;
wire   [4:0] \A[4][130] ;
wire   [4:0] \A[4][131] ;
wire   [4:0] \A[4][132] ;
wire   [4:0] \A[4][133] ;
wire   [4:0] \A[4][134] ;
wire   [4:0] \A[4][135] ;
wire   [4:0] \A[4][136] ;
wire   [4:0] \A[4][137] ;
wire   [4:0] \A[4][138] ;
wire   [4:0] \A[4][139] ;
wire   [4:0] \A[4][140] ;
wire   [4:0] \A[4][141] ;
wire   [4:0] \A[4][142] ;
wire   [4:0] \A[4][143] ;
wire   [4:0] \A[4][144] ;
wire   [4:0] \A[4][145] ;
wire   [4:0] \A[4][146] ;
wire   [4:0] \A[4][147] ;
wire   [4:0] \A[4][148] ;
wire   [4:0] \A[4][149] ;
wire   [4:0] \A[4][150] ;
wire   [4:0] \A[4][151] ;
wire   [4:0] \A[4][152] ;
wire   [4:0] \A[4][153] ;
wire   [4:0] \A[4][154] ;
wire   [4:0] \A[4][155] ;
wire   [4:0] \A[4][156] ;
wire   [4:0] \A[4][157] ;
wire   [4:0] \A[4][158] ;
wire   [4:0] \A[4][159] ;
wire   [4:0] \A[4][160] ;
wire   [4:0] \A[4][161] ;
wire   [4:0] \A[4][162] ;
wire   [4:0] \A[4][163] ;
wire   [4:0] \A[4][164] ;
wire   [4:0] \A[4][165] ;
wire   [4:0] \A[4][166] ;
wire   [4:0] \A[4][167] ;
wire   [4:0] \A[4][168] ;
wire   [4:0] \A[4][169] ;
wire   [4:0] \A[4][170] ;
wire   [4:0] \A[4][171] ;
wire   [4:0] \A[4][172] ;
wire   [4:0] \A[4][173] ;
wire   [4:0] \A[4][174] ;
wire   [4:0] \A[4][175] ;
wire   [4:0] \A[4][176] ;
wire   [4:0] \A[4][177] ;
wire   [4:0] \A[4][178] ;
wire   [4:0] \A[4][179] ;
wire   [4:0] \A[4][180] ;
wire   [4:0] \A[4][181] ;
wire   [4:0] \A[4][182] ;
wire   [4:0] \A[4][183] ;
wire   [4:0] \A[4][184] ;
wire   [4:0] \A[4][185] ;
wire   [4:0] \A[4][186] ;
wire   [4:0] \A[4][187] ;
wire   [4:0] \A[4][188] ;
wire   [4:0] \A[4][189] ;
wire   [4:0] \A[4][190] ;
wire   [4:0] \A[4][191] ;
wire   [4:0] \A[4][192] ;
wire   [4:0] \A[4][193] ;
wire   [4:0] \A[4][194] ;
wire   [4:0] \A[4][195] ;
wire   [4:0] \A[4][196] ;
wire   [4:0] \A[4][197] ;
wire   [4:0] \A[4][198] ;
wire   [4:0] \A[4][199] ;
wire   [4:0] \A[4][200] ;
wire   [4:0] \A[4][201] ;
wire   [4:0] \A[4][202] ;
wire   [4:0] \A[4][203] ;
wire   [4:0] \A[4][204] ;
wire   [4:0] \A[4][205] ;
wire   [4:0] \A[4][206] ;
wire   [4:0] \A[4][207] ;
wire   [4:0] \A[4][208] ;
wire   [4:0] \A[4][209] ;
wire   [4:0] \A[4][210] ;
wire   [4:0] \A[4][211] ;
wire   [4:0] \A[4][212] ;
wire   [4:0] \A[4][213] ;
wire   [4:0] \A[4][214] ;
wire   [4:0] \A[4][215] ;
wire   [4:0] \A[4][216] ;
wire   [4:0] \A[4][217] ;
wire   [4:0] \A[4][218] ;
wire   [4:0] \A[4][219] ;
wire   [4:0] \A[4][220] ;
wire   [4:0] \A[4][221] ;
wire   [4:0] \A[4][222] ;
wire   [4:0] \A[4][223] ;
wire   [4:0] \A[4][224] ;
wire   [4:0] \A[4][225] ;
wire   [4:0] \A[4][226] ;
wire   [4:0] \A[4][227] ;
wire   [4:0] \A[4][228] ;
wire   [4:0] \A[4][229] ;
wire   [4:0] \A[4][230] ;
wire   [4:0] \A[4][231] ;
wire   [4:0] \A[4][232] ;
wire   [4:0] \A[4][233] ;
wire   [4:0] \A[4][234] ;
wire   [4:0] \A[4][235] ;
wire   [4:0] \A[4][236] ;
wire   [4:0] \A[4][237] ;
wire   [4:0] \A[4][238] ;
wire   [4:0] \A[4][239] ;
wire   [4:0] \A[4][240] ;
wire   [4:0] \A[4][241] ;
wire   [4:0] \A[4][242] ;
wire   [4:0] \A[4][243] ;
wire   [4:0] \A[4][244] ;
wire   [4:0] \A[4][245] ;
wire   [4:0] \A[4][246] ;
wire   [4:0] \A[4][247] ;
wire   [4:0] \A[4][248] ;
wire   [4:0] \A[4][249] ;
wire   [4:0] \A[4][250] ;
wire   [4:0] \A[4][251] ;
wire   [4:0] \A[4][252] ;
wire   [4:0] \A[4][253] ;
wire   [4:0] \A[4][254] ;
wire   [4:0] \A[4][255] ;
wire   [4:0] \A[5][0] ;
wire   [4:0] \A[5][1] ;
wire   [4:0] \A[5][2] ;
wire   [4:0] \A[5][3] ;
wire   [4:0] \A[5][4] ;
wire   [4:0] \A[5][5] ;
wire   [4:0] \A[5][6] ;
wire   [4:0] \A[5][7] ;
wire   [4:0] \A[5][8] ;
wire   [4:0] \A[5][9] ;
wire   [4:0] \A[5][10] ;
wire   [4:0] \A[5][11] ;
wire   [4:0] \A[5][12] ;
wire   [4:0] \A[5][13] ;
wire   [4:0] \A[5][14] ;
wire   [4:0] \A[5][15] ;
wire   [4:0] \A[5][16] ;
wire   [4:0] \A[5][17] ;
wire   [4:0] \A[5][18] ;
wire   [4:0] \A[5][19] ;
wire   [4:0] \A[5][20] ;
wire   [4:0] \A[5][21] ;
wire   [4:0] \A[5][22] ;
wire   [4:0] \A[5][23] ;
wire   [4:0] \A[5][24] ;
wire   [4:0] \A[5][25] ;
wire   [4:0] \A[5][26] ;
wire   [4:0] \A[5][27] ;
wire   [4:0] \A[5][28] ;
wire   [4:0] \A[5][29] ;
wire   [4:0] \A[5][30] ;
wire   [4:0] \A[5][31] ;
wire   [4:0] \A[5][32] ;
wire   [4:0] \A[5][33] ;
wire   [4:0] \A[5][34] ;
wire   [4:0] \A[5][35] ;
wire   [4:0] \A[5][36] ;
wire   [4:0] \A[5][37] ;
wire   [4:0] \A[5][38] ;
wire   [4:0] \A[5][39] ;
wire   [4:0] \A[5][40] ;
wire   [4:0] \A[5][41] ;
wire   [4:0] \A[5][42] ;
wire   [4:0] \A[5][43] ;
wire   [4:0] \A[5][44] ;
wire   [4:0] \A[5][45] ;
wire   [4:0] \A[5][46] ;
wire   [4:0] \A[5][47] ;
wire   [4:0] \A[5][48] ;
wire   [4:0] \A[5][49] ;
wire   [4:0] \A[5][50] ;
wire   [4:0] \A[5][51] ;
wire   [4:0] \A[5][52] ;
wire   [4:0] \A[5][53] ;
wire   [4:0] \A[5][54] ;
wire   [4:0] \A[5][55] ;
wire   [4:0] \A[5][56] ;
wire   [4:0] \A[5][57] ;
wire   [4:0] \A[5][58] ;
wire   [4:0] \A[5][59] ;
wire   [4:0] \A[5][60] ;
wire   [4:0] \A[5][61] ;
wire   [4:0] \A[5][62] ;
wire   [4:0] \A[5][63] ;
wire   [4:0] \A[5][64] ;
wire   [4:0] \A[5][65] ;
wire   [4:0] \A[5][66] ;
wire   [4:0] \A[5][67] ;
wire   [4:0] \A[5][68] ;
wire   [4:0] \A[5][69] ;
wire   [4:0] \A[5][70] ;
wire   [4:0] \A[5][71] ;
wire   [4:0] \A[5][72] ;
wire   [4:0] \A[5][73] ;
wire   [4:0] \A[5][74] ;
wire   [4:0] \A[5][75] ;
wire   [4:0] \A[5][76] ;
wire   [4:0] \A[5][77] ;
wire   [4:0] \A[5][78] ;
wire   [4:0] \A[5][79] ;
wire   [4:0] \A[5][80] ;
wire   [4:0] \A[5][81] ;
wire   [4:0] \A[5][82] ;
wire   [4:0] \A[5][83] ;
wire   [4:0] \A[5][84] ;
wire   [4:0] \A[5][85] ;
wire   [4:0] \A[5][86] ;
wire   [4:0] \A[5][87] ;
wire   [4:0] \A[5][88] ;
wire   [4:0] \A[5][89] ;
wire   [4:0] \A[5][90] ;
wire   [4:0] \A[5][91] ;
wire   [4:0] \A[5][92] ;
wire   [4:0] \A[5][93] ;
wire   [4:0] \A[5][94] ;
wire   [4:0] \A[5][95] ;
wire   [4:0] \A[5][96] ;
wire   [4:0] \A[5][97] ;
wire   [4:0] \A[5][98] ;
wire   [4:0] \A[5][99] ;
wire   [4:0] \A[5][100] ;
wire   [4:0] \A[5][101] ;
wire   [4:0] \A[5][102] ;
wire   [4:0] \A[5][103] ;
wire   [4:0] \A[5][104] ;
wire   [4:0] \A[5][105] ;
wire   [4:0] \A[5][106] ;
wire   [4:0] \A[5][107] ;
wire   [4:0] \A[5][108] ;
wire   [4:0] \A[5][109] ;
wire   [4:0] \A[5][110] ;
wire   [4:0] \A[5][111] ;
wire   [4:0] \A[5][112] ;
wire   [4:0] \A[5][113] ;
wire   [4:0] \A[5][114] ;
wire   [4:0] \A[5][115] ;
wire   [4:0] \A[5][116] ;
wire   [4:0] \A[5][117] ;
wire   [4:0] \A[5][118] ;
wire   [4:0] \A[5][119] ;
wire   [4:0] \A[5][120] ;
wire   [4:0] \A[5][121] ;
wire   [4:0] \A[5][122] ;
wire   [4:0] \A[5][123] ;
wire   [4:0] \A[5][124] ;
wire   [4:0] \A[5][125] ;
wire   [4:0] \A[5][126] ;
wire   [4:0] \A[5][127] ;
wire   [4:0] \A[5][128] ;
wire   [4:0] \A[5][129] ;
wire   [4:0] \A[5][130] ;
wire   [4:0] \A[5][131] ;
wire   [4:0] \A[5][132] ;
wire   [4:0] \A[5][133] ;
wire   [4:0] \A[5][134] ;
wire   [4:0] \A[5][135] ;
wire   [4:0] \A[5][136] ;
wire   [4:0] \A[5][137] ;
wire   [4:0] \A[5][138] ;
wire   [4:0] \A[5][139] ;
wire   [4:0] \A[5][140] ;
wire   [4:0] \A[5][141] ;
wire   [4:0] \A[5][142] ;
wire   [4:0] \A[5][143] ;
wire   [4:0] \A[5][144] ;
wire   [4:0] \A[5][145] ;
wire   [4:0] \A[5][146] ;
wire   [4:0] \A[5][147] ;
wire   [4:0] \A[5][148] ;
wire   [4:0] \A[5][149] ;
wire   [4:0] \A[5][150] ;
wire   [4:0] \A[5][151] ;
wire   [4:0] \A[5][152] ;
wire   [4:0] \A[5][153] ;
wire   [4:0] \A[5][154] ;
wire   [4:0] \A[5][155] ;
wire   [4:0] \A[5][156] ;
wire   [4:0] \A[5][157] ;
wire   [4:0] \A[5][158] ;
wire   [4:0] \A[5][159] ;
wire   [4:0] \A[5][160] ;
wire   [4:0] \A[5][161] ;
wire   [4:0] \A[5][162] ;
wire   [4:0] \A[5][163] ;
wire   [4:0] \A[5][164] ;
wire   [4:0] \A[5][165] ;
wire   [4:0] \A[5][166] ;
wire   [4:0] \A[5][167] ;
wire   [4:0] \A[5][168] ;
wire   [4:0] \A[5][169] ;
wire   [4:0] \A[5][170] ;
wire   [4:0] \A[5][171] ;
wire   [4:0] \A[5][172] ;
wire   [4:0] \A[5][173] ;
wire   [4:0] \A[5][174] ;
wire   [4:0] \A[5][175] ;
wire   [4:0] \A[5][176] ;
wire   [4:0] \A[5][177] ;
wire   [4:0] \A[5][178] ;
wire   [4:0] \A[5][179] ;
wire   [4:0] \A[5][180] ;
wire   [4:0] \A[5][181] ;
wire   [4:0] \A[5][182] ;
wire   [4:0] \A[5][183] ;
wire   [4:0] \A[5][184] ;
wire   [4:0] \A[5][185] ;
wire   [4:0] \A[5][186] ;
wire   [4:0] \A[5][187] ;
wire   [4:0] \A[5][188] ;
wire   [4:0] \A[5][189] ;
wire   [4:0] \A[5][190] ;
wire   [4:0] \A[5][191] ;
wire   [4:0] \A[5][192] ;
wire   [4:0] \A[5][193] ;
wire   [4:0] \A[5][194] ;
wire   [4:0] \A[5][195] ;
wire   [4:0] \A[5][196] ;
wire   [4:0] \A[5][197] ;
wire   [4:0] \A[5][198] ;
wire   [4:0] \A[5][199] ;
wire   [4:0] \A[5][200] ;
wire   [4:0] \A[5][201] ;
wire   [4:0] \A[5][202] ;
wire   [4:0] \A[5][203] ;
wire   [4:0] \A[5][204] ;
wire   [4:0] \A[5][205] ;
wire   [4:0] \A[5][206] ;
wire   [4:0] \A[5][207] ;
wire   [4:0] \A[5][208] ;
wire   [4:0] \A[5][209] ;
wire   [4:0] \A[5][210] ;
wire   [4:0] \A[5][211] ;
wire   [4:0] \A[5][212] ;
wire   [4:0] \A[5][213] ;
wire   [4:0] \A[5][214] ;
wire   [4:0] \A[5][215] ;
wire   [4:0] \A[5][216] ;
wire   [4:0] \A[5][217] ;
wire   [4:0] \A[5][218] ;
wire   [4:0] \A[5][219] ;
wire   [4:0] \A[5][220] ;
wire   [4:0] \A[5][221] ;
wire   [4:0] \A[5][222] ;
wire   [4:0] \A[5][223] ;
wire   [4:0] \A[5][224] ;
wire   [4:0] \A[5][225] ;
wire   [4:0] \A[5][226] ;
wire   [4:0] \A[5][227] ;
wire   [4:0] \A[5][228] ;
wire   [4:0] \A[5][229] ;
wire   [4:0] \A[5][230] ;
wire   [4:0] \A[5][231] ;
wire   [4:0] \A[5][232] ;
wire   [4:0] \A[5][233] ;
wire   [4:0] \A[5][234] ;
wire   [4:0] \A[5][235] ;
wire   [4:0] \A[5][236] ;
wire   [4:0] \A[5][237] ;
wire   [4:0] \A[5][238] ;
wire   [4:0] \A[5][239] ;
wire   [4:0] \A[5][240] ;
wire   [4:0] \A[5][241] ;
wire   [4:0] \A[5][242] ;
wire   [4:0] \A[5][243] ;
wire   [4:0] \A[5][244] ;
wire   [4:0] \A[5][245] ;
wire   [4:0] \A[5][246] ;
wire   [4:0] \A[5][247] ;
wire   [4:0] \A[5][248] ;
wire   [4:0] \A[5][249] ;
wire   [4:0] \A[5][250] ;
wire   [4:0] \A[5][251] ;
wire   [4:0] \A[5][252] ;
wire   [4:0] \A[5][253] ;
wire   [4:0] \A[5][254] ;
wire   [4:0] \A[5][255] ;
wire   [4:0] \A[6][0] ;
wire   [4:0] \A[6][1] ;
wire   [4:0] \A[6][2] ;
wire   [4:0] \A[6][3] ;
wire   [4:0] \A[6][4] ;
wire   [4:0] \A[6][5] ;
wire   [4:0] \A[6][6] ;
wire   [4:0] \A[6][7] ;
wire   [4:0] \A[6][8] ;
wire   [4:0] \A[6][9] ;
wire   [4:0] \A[6][10] ;
wire   [4:0] \A[6][11] ;
wire   [4:0] \A[6][12] ;
wire   [4:0] \A[6][13] ;
wire   [4:0] \A[6][14] ;
wire   [4:0] \A[6][15] ;
wire   [4:0] \A[6][16] ;
wire   [4:0] \A[6][17] ;
wire   [4:0] \A[6][18] ;
wire   [4:0] \A[6][19] ;
wire   [4:0] \A[6][20] ;
wire   [4:0] \A[6][21] ;
wire   [4:0] \A[6][22] ;
wire   [4:0] \A[6][23] ;
wire   [4:0] \A[6][24] ;
wire   [4:0] \A[6][25] ;
wire   [4:0] \A[6][26] ;
wire   [4:0] \A[6][27] ;
wire   [4:0] \A[6][28] ;
wire   [4:0] \A[6][29] ;
wire   [4:0] \A[6][30] ;
wire   [4:0] \A[6][31] ;
wire   [4:0] \A[6][32] ;
wire   [4:0] \A[6][33] ;
wire   [4:0] \A[6][34] ;
wire   [4:0] \A[6][35] ;
wire   [4:0] \A[6][36] ;
wire   [4:0] \A[6][37] ;
wire   [4:0] \A[6][38] ;
wire   [4:0] \A[6][39] ;
wire   [4:0] \A[6][40] ;
wire   [4:0] \A[6][41] ;
wire   [4:0] \A[6][42] ;
wire   [4:0] \A[6][43] ;
wire   [4:0] \A[6][44] ;
wire   [4:0] \A[6][45] ;
wire   [4:0] \A[6][46] ;
wire   [4:0] \A[6][47] ;
wire   [4:0] \A[6][48] ;
wire   [4:0] \A[6][49] ;
wire   [4:0] \A[6][50] ;
wire   [4:0] \A[6][51] ;
wire   [4:0] \A[6][52] ;
wire   [4:0] \A[6][53] ;
wire   [4:0] \A[6][54] ;
wire   [4:0] \A[6][55] ;
wire   [4:0] \A[6][56] ;
wire   [4:0] \A[6][57] ;
wire   [4:0] \A[6][58] ;
wire   [4:0] \A[6][59] ;
wire   [4:0] \A[6][60] ;
wire   [4:0] \A[6][61] ;
wire   [4:0] \A[6][62] ;
wire   [4:0] \A[6][63] ;
wire   [4:0] \A[6][64] ;
wire   [4:0] \A[6][65] ;
wire   [4:0] \A[6][66] ;
wire   [4:0] \A[6][67] ;
wire   [4:0] \A[6][68] ;
wire   [4:0] \A[6][69] ;
wire   [4:0] \A[6][70] ;
wire   [4:0] \A[6][71] ;
wire   [4:0] \A[6][72] ;
wire   [4:0] \A[6][73] ;
wire   [4:0] \A[6][74] ;
wire   [4:0] \A[6][75] ;
wire   [4:0] \A[6][76] ;
wire   [4:0] \A[6][77] ;
wire   [4:0] \A[6][78] ;
wire   [4:0] \A[6][79] ;
wire   [4:0] \A[6][80] ;
wire   [4:0] \A[6][81] ;
wire   [4:0] \A[6][82] ;
wire   [4:0] \A[6][83] ;
wire   [4:0] \A[6][84] ;
wire   [4:0] \A[6][85] ;
wire   [4:0] \A[6][86] ;
wire   [4:0] \A[6][87] ;
wire   [4:0] \A[6][88] ;
wire   [4:0] \A[6][89] ;
wire   [4:0] \A[6][90] ;
wire   [4:0] \A[6][91] ;
wire   [4:0] \A[6][92] ;
wire   [4:0] \A[6][93] ;
wire   [4:0] \A[6][94] ;
wire   [4:0] \A[6][95] ;
wire   [4:0] \A[6][96] ;
wire   [4:0] \A[6][97] ;
wire   [4:0] \A[6][98] ;
wire   [4:0] \A[6][99] ;
wire   [4:0] \A[6][100] ;
wire   [4:0] \A[6][101] ;
wire   [4:0] \A[6][102] ;
wire   [4:0] \A[6][103] ;
wire   [4:0] \A[6][104] ;
wire   [4:0] \A[6][105] ;
wire   [4:0] \A[6][106] ;
wire   [4:0] \A[6][107] ;
wire   [4:0] \A[6][108] ;
wire   [4:0] \A[6][109] ;
wire   [4:0] \A[6][110] ;
wire   [4:0] \A[6][111] ;
wire   [4:0] \A[6][112] ;
wire   [4:0] \A[6][113] ;
wire   [4:0] \A[6][114] ;
wire   [4:0] \A[6][115] ;
wire   [4:0] \A[6][116] ;
wire   [4:0] \A[6][117] ;
wire   [4:0] \A[6][118] ;
wire   [4:0] \A[6][119] ;
wire   [4:0] \A[6][120] ;
wire   [4:0] \A[6][121] ;
wire   [4:0] \A[6][122] ;
wire   [4:0] \A[6][123] ;
wire   [4:0] \A[6][124] ;
wire   [4:0] \A[6][125] ;
wire   [4:0] \A[6][126] ;
wire   [4:0] \A[6][127] ;
wire   [4:0] \A[6][128] ;
wire   [4:0] \A[6][129] ;
wire   [4:0] \A[6][130] ;
wire   [4:0] \A[6][131] ;
wire   [4:0] \A[6][132] ;
wire   [4:0] \A[6][133] ;
wire   [4:0] \A[6][134] ;
wire   [4:0] \A[6][135] ;
wire   [4:0] \A[6][136] ;
wire   [4:0] \A[6][137] ;
wire   [4:0] \A[6][138] ;
wire   [4:0] \A[6][139] ;
wire   [4:0] \A[6][140] ;
wire   [4:0] \A[6][141] ;
wire   [4:0] \A[6][142] ;
wire   [4:0] \A[6][143] ;
wire   [4:0] \A[6][144] ;
wire   [4:0] \A[6][145] ;
wire   [4:0] \A[6][146] ;
wire   [4:0] \A[6][147] ;
wire   [4:0] \A[6][148] ;
wire   [4:0] \A[6][149] ;
wire   [4:0] \A[6][150] ;
wire   [4:0] \A[6][151] ;
wire   [4:0] \A[6][152] ;
wire   [4:0] \A[6][153] ;
wire   [4:0] \A[6][154] ;
wire   [4:0] \A[6][155] ;
wire   [4:0] \A[6][156] ;
wire   [4:0] \A[6][157] ;
wire   [4:0] \A[6][158] ;
wire   [4:0] \A[6][159] ;
wire   [4:0] \A[6][160] ;
wire   [4:0] \A[6][161] ;
wire   [4:0] \A[6][162] ;
wire   [4:0] \A[6][163] ;
wire   [4:0] \A[6][164] ;
wire   [4:0] \A[6][165] ;
wire   [4:0] \A[6][166] ;
wire   [4:0] \A[6][167] ;
wire   [4:0] \A[6][168] ;
wire   [4:0] \A[6][169] ;
wire   [4:0] \A[6][170] ;
wire   [4:0] \A[6][171] ;
wire   [4:0] \A[6][172] ;
wire   [4:0] \A[6][173] ;
wire   [4:0] \A[6][174] ;
wire   [4:0] \A[6][175] ;
wire   [4:0] \A[6][176] ;
wire   [4:0] \A[6][177] ;
wire   [4:0] \A[6][178] ;
wire   [4:0] \A[6][179] ;
wire   [4:0] \A[6][180] ;
wire   [4:0] \A[6][181] ;
wire   [4:0] \A[6][182] ;
wire   [4:0] \A[6][183] ;
wire   [4:0] \A[6][184] ;
wire   [4:0] \A[6][185] ;
wire   [4:0] \A[6][186] ;
wire   [4:0] \A[6][187] ;
wire   [4:0] \A[6][188] ;
wire   [4:0] \A[6][189] ;
wire   [4:0] \A[6][190] ;
wire   [4:0] \A[6][191] ;
wire   [4:0] \A[6][192] ;
wire   [4:0] \A[6][193] ;
wire   [4:0] \A[6][194] ;
wire   [4:0] \A[6][195] ;
wire   [4:0] \A[6][196] ;
wire   [4:0] \A[6][197] ;
wire   [4:0] \A[6][198] ;
wire   [4:0] \A[6][199] ;
wire   [4:0] \A[6][200] ;
wire   [4:0] \A[6][201] ;
wire   [4:0] \A[6][202] ;
wire   [4:0] \A[6][203] ;
wire   [4:0] \A[6][204] ;
wire   [4:0] \A[6][205] ;
wire   [4:0] \A[6][206] ;
wire   [4:0] \A[6][207] ;
wire   [4:0] \A[6][208] ;
wire   [4:0] \A[6][209] ;
wire   [4:0] \A[6][210] ;
wire   [4:0] \A[6][211] ;
wire   [4:0] \A[6][212] ;
wire   [4:0] \A[6][213] ;
wire   [4:0] \A[6][214] ;
wire   [4:0] \A[6][215] ;
wire   [4:0] \A[6][216] ;
wire   [4:0] \A[6][217] ;
wire   [4:0] \A[6][218] ;
wire   [4:0] \A[6][219] ;
wire   [4:0] \A[6][220] ;
wire   [4:0] \A[6][221] ;
wire   [4:0] \A[6][222] ;
wire   [4:0] \A[6][223] ;
wire   [4:0] \A[6][224] ;
wire   [4:0] \A[6][225] ;
wire   [4:0] \A[6][226] ;
wire   [4:0] \A[6][227] ;
wire   [4:0] \A[6][228] ;
wire   [4:0] \A[6][229] ;
wire   [4:0] \A[6][230] ;
wire   [4:0] \A[6][231] ;
wire   [4:0] \A[6][232] ;
wire   [4:0] \A[6][233] ;
wire   [4:0] \A[6][234] ;
wire   [4:0] \A[6][235] ;
wire   [4:0] \A[6][236] ;
wire   [4:0] \A[6][237] ;
wire   [4:0] \A[6][238] ;
wire   [4:0] \A[6][239] ;
wire   [4:0] \A[6][240] ;
wire   [4:0] \A[6][241] ;
wire   [4:0] \A[6][242] ;
wire   [4:0] \A[6][243] ;
wire   [4:0] \A[6][244] ;
wire   [4:0] \A[6][245] ;
wire   [4:0] \A[6][246] ;
wire   [4:0] \A[6][247] ;
wire   [4:0] \A[6][248] ;
wire   [4:0] \A[6][249] ;
wire   [4:0] \A[6][250] ;
wire   [4:0] \A[6][251] ;
wire   [4:0] \A[6][252] ;
wire   [4:0] \A[6][253] ;
wire   [4:0] \A[6][254] ;
wire   [4:0] \A[6][255] ;
wire   [4:0] \A[7][0] ;
wire   [4:0] \A[7][1] ;
wire   [4:0] \A[7][2] ;
wire   [4:0] \A[7][3] ;
wire   [4:0] \A[7][4] ;
wire   [4:0] \A[7][5] ;
wire   [4:0] \A[7][6] ;
wire   [4:0] \A[7][7] ;
wire   [4:0] \A[7][8] ;
wire   [4:0] \A[7][9] ;
wire   [4:0] \A[7][10] ;
wire   [4:0] \A[7][11] ;
wire   [4:0] \A[7][12] ;
wire   [4:0] \A[7][13] ;
wire   [4:0] \A[7][14] ;
wire   [4:0] \A[7][15] ;
wire   [4:0] \A[7][16] ;
wire   [4:0] \A[7][17] ;
wire   [4:0] \A[7][18] ;
wire   [4:0] \A[7][19] ;
wire   [4:0] \A[7][20] ;
wire   [4:0] \A[7][21] ;
wire   [4:0] \A[7][22] ;
wire   [4:0] \A[7][23] ;
wire   [4:0] \A[7][24] ;
wire   [4:0] \A[7][25] ;
wire   [4:0] \A[7][26] ;
wire   [4:0] \A[7][27] ;
wire   [4:0] \A[7][28] ;
wire   [4:0] \A[7][29] ;
wire   [4:0] \A[7][30] ;
wire   [4:0] \A[7][31] ;
wire   [4:0] \A[7][32] ;
wire   [4:0] \A[7][33] ;
wire   [4:0] \A[7][34] ;
wire   [4:0] \A[7][35] ;
wire   [4:0] \A[7][36] ;
wire   [4:0] \A[7][37] ;
wire   [4:0] \A[7][38] ;
wire   [4:0] \A[7][39] ;
wire   [4:0] \A[7][40] ;
wire   [4:0] \A[7][41] ;
wire   [4:0] \A[7][42] ;
wire   [4:0] \A[7][43] ;
wire   [4:0] \A[7][44] ;
wire   [4:0] \A[7][45] ;
wire   [4:0] \A[7][46] ;
wire   [4:0] \A[7][47] ;
wire   [4:0] \A[7][48] ;
wire   [4:0] \A[7][49] ;
wire   [4:0] \A[7][50] ;
wire   [4:0] \A[7][51] ;
wire   [4:0] \A[7][52] ;
wire   [4:0] \A[7][53] ;
wire   [4:0] \A[7][54] ;
wire   [4:0] \A[7][55] ;
wire   [4:0] \A[7][56] ;
wire   [4:0] \A[7][57] ;
wire   [4:0] \A[7][58] ;
wire   [4:0] \A[7][59] ;
wire   [4:0] \A[7][60] ;
wire   [4:0] \A[7][61] ;
wire   [4:0] \A[7][62] ;
wire   [4:0] \A[7][63] ;
wire   [4:0] \A[7][64] ;
wire   [4:0] \A[7][65] ;
wire   [4:0] \A[7][66] ;
wire   [4:0] \A[7][67] ;
wire   [4:0] \A[7][68] ;
wire   [4:0] \A[7][69] ;
wire   [4:0] \A[7][70] ;
wire   [4:0] \A[7][71] ;
wire   [4:0] \A[7][72] ;
wire   [4:0] \A[7][73] ;
wire   [4:0] \A[7][74] ;
wire   [4:0] \A[7][75] ;
wire   [4:0] \A[7][76] ;
wire   [4:0] \A[7][77] ;
wire   [4:0] \A[7][78] ;
wire   [4:0] \A[7][79] ;
wire   [4:0] \A[7][80] ;
wire   [4:0] \A[7][81] ;
wire   [4:0] \A[7][82] ;
wire   [4:0] \A[7][83] ;
wire   [4:0] \A[7][84] ;
wire   [4:0] \A[7][85] ;
wire   [4:0] \A[7][86] ;
wire   [4:0] \A[7][87] ;
wire   [4:0] \A[7][88] ;
wire   [4:0] \A[7][89] ;
wire   [4:0] \A[7][90] ;
wire   [4:0] \A[7][91] ;
wire   [4:0] \A[7][92] ;
wire   [4:0] \A[7][93] ;
wire   [4:0] \A[7][94] ;
wire   [4:0] \A[7][95] ;
wire   [4:0] \A[7][96] ;
wire   [4:0] \A[7][97] ;
wire   [4:0] \A[7][98] ;
wire   [4:0] \A[7][99] ;
wire   [4:0] \A[7][100] ;
wire   [4:0] \A[7][101] ;
wire   [4:0] \A[7][102] ;
wire   [4:0] \A[7][103] ;
wire   [4:0] \A[7][104] ;
wire   [4:0] \A[7][105] ;
wire   [4:0] \A[7][106] ;
wire   [4:0] \A[7][107] ;
wire   [4:0] \A[7][108] ;
wire   [4:0] \A[7][109] ;
wire   [4:0] \A[7][110] ;
wire   [4:0] \A[7][111] ;
wire   [4:0] \A[7][112] ;
wire   [4:0] \A[7][113] ;
wire   [4:0] \A[7][114] ;
wire   [4:0] \A[7][115] ;
wire   [4:0] \A[7][116] ;
wire   [4:0] \A[7][117] ;
wire   [4:0] \A[7][118] ;
wire   [4:0] \A[7][119] ;
wire   [4:0] \A[7][120] ;
wire   [4:0] \A[7][121] ;
wire   [4:0] \A[7][122] ;
wire   [4:0] \A[7][123] ;
wire   [4:0] \A[7][124] ;
wire   [4:0] \A[7][125] ;
wire   [4:0] \A[7][126] ;
wire   [4:0] \A[7][127] ;
wire   [4:0] \A[7][128] ;
wire   [4:0] \A[7][129] ;
wire   [4:0] \A[7][130] ;
wire   [4:0] \A[7][131] ;
wire   [4:0] \A[7][132] ;
wire   [4:0] \A[7][133] ;
wire   [4:0] \A[7][134] ;
wire   [4:0] \A[7][135] ;
wire   [4:0] \A[7][136] ;
wire   [4:0] \A[7][137] ;
wire   [4:0] \A[7][138] ;
wire   [4:0] \A[7][139] ;
wire   [4:0] \A[7][140] ;
wire   [4:0] \A[7][141] ;
wire   [4:0] \A[7][142] ;
wire   [4:0] \A[7][143] ;
wire   [4:0] \A[7][144] ;
wire   [4:0] \A[7][145] ;
wire   [4:0] \A[7][146] ;
wire   [4:0] \A[7][147] ;
wire   [4:0] \A[7][148] ;
wire   [4:0] \A[7][149] ;
wire   [4:0] \A[7][150] ;
wire   [4:0] \A[7][151] ;
wire   [4:0] \A[7][152] ;
wire   [4:0] \A[7][153] ;
wire   [4:0] \A[7][154] ;
wire   [4:0] \A[7][155] ;
wire   [4:0] \A[7][156] ;
wire   [4:0] \A[7][157] ;
wire   [4:0] \A[7][158] ;
wire   [4:0] \A[7][159] ;
wire   [4:0] \A[7][160] ;
wire   [4:0] \A[7][161] ;
wire   [4:0] \A[7][162] ;
wire   [4:0] \A[7][163] ;
wire   [4:0] \A[7][164] ;
wire   [4:0] \A[7][165] ;
wire   [4:0] \A[7][166] ;
wire   [4:0] \A[7][167] ;
wire   [4:0] \A[7][168] ;
wire   [4:0] \A[7][169] ;
wire   [4:0] \A[7][170] ;
wire   [4:0] \A[7][171] ;
wire   [4:0] \A[7][172] ;
wire   [4:0] \A[7][173] ;
wire   [4:0] \A[7][174] ;
wire   [4:0] \A[7][175] ;
wire   [4:0] \A[7][176] ;
wire   [4:0] \A[7][177] ;
wire   [4:0] \A[7][178] ;
wire   [4:0] \A[7][179] ;
wire   [4:0] \A[7][180] ;
wire   [4:0] \A[7][181] ;
wire   [4:0] \A[7][182] ;
wire   [4:0] \A[7][183] ;
wire   [4:0] \A[7][184] ;
wire   [4:0] \A[7][185] ;
wire   [4:0] \A[7][186] ;
wire   [4:0] \A[7][187] ;
wire   [4:0] \A[7][188] ;
wire   [4:0] \A[7][189] ;
wire   [4:0] \A[7][190] ;
wire   [4:0] \A[7][191] ;
wire   [4:0] \A[7][192] ;
wire   [4:0] \A[7][193] ;
wire   [4:0] \A[7][194] ;
wire   [4:0] \A[7][195] ;
wire   [4:0] \A[7][196] ;
wire   [4:0] \A[7][197] ;
wire   [4:0] \A[7][198] ;
wire   [4:0] \A[7][199] ;
wire   [4:0] \A[7][200] ;
wire   [4:0] \A[7][201] ;
wire   [4:0] \A[7][202] ;
wire   [4:0] \A[7][203] ;
wire   [4:0] \A[7][204] ;
wire   [4:0] \A[7][205] ;
wire   [4:0] \A[7][206] ;
wire   [4:0] \A[7][207] ;
wire   [4:0] \A[7][208] ;
wire   [4:0] \A[7][209] ;
wire   [4:0] \A[7][210] ;
wire   [4:0] \A[7][211] ;
wire   [4:0] \A[7][212] ;
wire   [4:0] \A[7][213] ;
wire   [4:0] \A[7][214] ;
wire   [4:0] \A[7][215] ;
wire   [4:0] \A[7][216] ;
wire   [4:0] \A[7][217] ;
wire   [4:0] \A[7][218] ;
wire   [4:0] \A[7][219] ;
wire   [4:0] \A[7][220] ;
wire   [4:0] \A[7][221] ;
wire   [4:0] \A[7][222] ;
wire   [4:0] \A[7][223] ;
wire   [4:0] \A[7][224] ;
wire   [4:0] \A[7][225] ;
wire   [4:0] \A[7][226] ;
wire   [4:0] \A[7][227] ;
wire   [4:0] \A[7][228] ;
wire   [4:0] \A[7][229] ;
wire   [4:0] \A[7][230] ;
wire   [4:0] \A[7][231] ;
wire   [4:0] \A[7][232] ;
wire   [4:0] \A[7][233] ;
wire   [4:0] \A[7][234] ;
wire   [4:0] \A[7][235] ;
wire   [4:0] \A[7][236] ;
wire   [4:0] \A[7][237] ;
wire   [4:0] \A[7][238] ;
wire   [4:0] \A[7][239] ;
wire   [4:0] \A[7][240] ;
wire   [4:0] \A[7][241] ;
wire   [4:0] \A[7][242] ;
wire   [4:0] \A[7][243] ;
wire   [4:0] \A[7][244] ;
wire   [4:0] \A[7][245] ;
wire   [4:0] \A[7][246] ;
wire   [4:0] \A[7][247] ;
wire   [4:0] \A[7][248] ;
wire   [4:0] \A[7][249] ;
wire   [4:0] \A[7][250] ;
wire   [4:0] \A[7][251] ;
wire   [4:0] \A[7][252] ;
wire   [4:0] \A[7][253] ;
wire   [4:0] \A[7][254] ;
wire   [4:0] \A[7][255] ;
wire   [4:0] \A[8][0] ;
wire   [4:0] \A[8][1] ;
wire   [4:0] \A[8][2] ;
wire   [4:0] \A[8][3] ;
wire   [4:0] \A[8][4] ;
wire   [4:0] \A[8][5] ;
wire   [4:0] \A[8][6] ;
wire   [4:0] \A[8][7] ;
wire   [4:0] \A[8][8] ;
wire   [4:0] \A[8][9] ;
wire   [4:0] \A[8][10] ;
wire   [4:0] \A[8][11] ;
wire   [4:0] \A[8][12] ;
wire   [4:0] \A[8][13] ;
wire   [4:0] \A[8][14] ;
wire   [4:0] \A[8][15] ;
wire   [4:0] \A[8][16] ;
wire   [4:0] \A[8][17] ;
wire   [4:0] \A[8][18] ;
wire   [4:0] \A[8][19] ;
wire   [4:0] \A[8][20] ;
wire   [4:0] \A[8][21] ;
wire   [4:0] \A[8][22] ;
wire   [4:0] \A[8][23] ;
wire   [4:0] \A[8][24] ;
wire   [4:0] \A[8][25] ;
wire   [4:0] \A[8][26] ;
wire   [4:0] \A[8][27] ;
wire   [4:0] \A[8][28] ;
wire   [4:0] \A[8][29] ;
wire   [4:0] \A[8][30] ;
wire   [4:0] \A[8][31] ;
wire   [4:0] \A[8][32] ;
wire   [4:0] \A[8][33] ;
wire   [4:0] \A[8][34] ;
wire   [4:0] \A[8][35] ;
wire   [4:0] \A[8][36] ;
wire   [4:0] \A[8][37] ;
wire   [4:0] \A[8][38] ;
wire   [4:0] \A[8][39] ;
wire   [4:0] \A[8][40] ;
wire   [4:0] \A[8][41] ;
wire   [4:0] \A[8][42] ;
wire   [4:0] \A[8][43] ;
wire   [4:0] \A[8][44] ;
wire   [4:0] \A[8][45] ;
wire   [4:0] \A[8][46] ;
wire   [4:0] \A[8][47] ;
wire   [4:0] \A[8][48] ;
wire   [4:0] \A[8][49] ;
wire   [4:0] \A[8][50] ;
wire   [4:0] \A[8][51] ;
wire   [4:0] \A[8][52] ;
wire   [4:0] \A[8][53] ;
wire   [4:0] \A[8][54] ;
wire   [4:0] \A[8][55] ;
wire   [4:0] \A[8][56] ;
wire   [4:0] \A[8][57] ;
wire   [4:0] \A[8][58] ;
wire   [4:0] \A[8][59] ;
wire   [4:0] \A[8][60] ;
wire   [4:0] \A[8][61] ;
wire   [4:0] \A[8][62] ;
wire   [4:0] \A[8][63] ;
wire   [4:0] \A[8][64] ;
wire   [4:0] \A[8][65] ;
wire   [4:0] \A[8][66] ;
wire   [4:0] \A[8][67] ;
wire   [4:0] \A[8][68] ;
wire   [4:0] \A[8][69] ;
wire   [4:0] \A[8][70] ;
wire   [4:0] \A[8][71] ;
wire   [4:0] \A[8][72] ;
wire   [4:0] \A[8][73] ;
wire   [4:0] \A[8][74] ;
wire   [4:0] \A[8][75] ;
wire   [4:0] \A[8][76] ;
wire   [4:0] \A[8][77] ;
wire   [4:0] \A[8][78] ;
wire   [4:0] \A[8][79] ;
wire   [4:0] \A[8][80] ;
wire   [4:0] \A[8][81] ;
wire   [4:0] \A[8][82] ;
wire   [4:0] \A[8][83] ;
wire   [4:0] \A[8][84] ;
wire   [4:0] \A[8][85] ;
wire   [4:0] \A[8][86] ;
wire   [4:0] \A[8][87] ;
wire   [4:0] \A[8][88] ;
wire   [4:0] \A[8][89] ;
wire   [4:0] \A[8][90] ;
wire   [4:0] \A[8][91] ;
wire   [4:0] \A[8][92] ;
wire   [4:0] \A[8][93] ;
wire   [4:0] \A[8][94] ;
wire   [4:0] \A[8][95] ;
wire   [4:0] \A[8][96] ;
wire   [4:0] \A[8][97] ;
wire   [4:0] \A[8][98] ;
wire   [4:0] \A[8][99] ;
wire   [4:0] \A[8][100] ;
wire   [4:0] \A[8][101] ;
wire   [4:0] \A[8][102] ;
wire   [4:0] \A[8][103] ;
wire   [4:0] \A[8][104] ;
wire   [4:0] \A[8][105] ;
wire   [4:0] \A[8][106] ;
wire   [4:0] \A[8][107] ;
wire   [4:0] \A[8][108] ;
wire   [4:0] \A[8][109] ;
wire   [4:0] \A[8][110] ;
wire   [4:0] \A[8][111] ;
wire   [4:0] \A[8][112] ;
wire   [4:0] \A[8][113] ;
wire   [4:0] \A[8][114] ;
wire   [4:0] \A[8][115] ;
wire   [4:0] \A[8][116] ;
wire   [4:0] \A[8][117] ;
wire   [4:0] \A[8][118] ;
wire   [4:0] \A[8][119] ;
wire   [4:0] \A[8][120] ;
wire   [4:0] \A[8][121] ;
wire   [4:0] \A[8][122] ;
wire   [4:0] \A[8][123] ;
wire   [4:0] \A[8][124] ;
wire   [4:0] \A[8][125] ;
wire   [4:0] \A[8][126] ;
wire   [4:0] \A[8][127] ;
wire   [4:0] \A[8][128] ;
wire   [4:0] \A[8][129] ;
wire   [4:0] \A[8][130] ;
wire   [4:0] \A[8][131] ;
wire   [4:0] \A[8][132] ;
wire   [4:0] \A[8][133] ;
wire   [4:0] \A[8][134] ;
wire   [4:0] \A[8][135] ;
wire   [4:0] \A[8][136] ;
wire   [4:0] \A[8][137] ;
wire   [4:0] \A[8][138] ;
wire   [4:0] \A[8][139] ;
wire   [4:0] \A[8][140] ;
wire   [4:0] \A[8][141] ;
wire   [4:0] \A[8][142] ;
wire   [4:0] \A[8][143] ;
wire   [4:0] \A[8][144] ;
wire   [4:0] \A[8][145] ;
wire   [4:0] \A[8][146] ;
wire   [4:0] \A[8][147] ;
wire   [4:0] \A[8][148] ;
wire   [4:0] \A[8][149] ;
wire   [4:0] \A[8][150] ;
wire   [4:0] \A[8][151] ;
wire   [4:0] \A[8][152] ;
wire   [4:0] \A[8][153] ;
wire   [4:0] \A[8][154] ;
wire   [4:0] \A[8][155] ;
wire   [4:0] \A[8][156] ;
wire   [4:0] \A[8][157] ;
wire   [4:0] \A[8][158] ;
wire   [4:0] \A[8][159] ;
wire   [4:0] \A[8][160] ;
wire   [4:0] \A[8][161] ;
wire   [4:0] \A[8][162] ;
wire   [4:0] \A[8][163] ;
wire   [4:0] \A[8][164] ;
wire   [4:0] \A[8][165] ;
wire   [4:0] \A[8][166] ;
wire   [4:0] \A[8][167] ;
wire   [4:0] \A[8][168] ;
wire   [4:0] \A[8][169] ;
wire   [4:0] \A[8][170] ;
wire   [4:0] \A[8][171] ;
wire   [4:0] \A[8][172] ;
wire   [4:0] \A[8][173] ;
wire   [4:0] \A[8][174] ;
wire   [4:0] \A[8][175] ;
wire   [4:0] \A[8][176] ;
wire   [4:0] \A[8][177] ;
wire   [4:0] \A[8][178] ;
wire   [4:0] \A[8][179] ;
wire   [4:0] \A[8][180] ;
wire   [4:0] \A[8][181] ;
wire   [4:0] \A[8][182] ;
wire   [4:0] \A[8][183] ;
wire   [4:0] \A[8][184] ;
wire   [4:0] \A[8][185] ;
wire   [4:0] \A[8][186] ;
wire   [4:0] \A[8][187] ;
wire   [4:0] \A[8][188] ;
wire   [4:0] \A[8][189] ;
wire   [4:0] \A[8][190] ;
wire   [4:0] \A[8][191] ;
wire   [4:0] \A[8][192] ;
wire   [4:0] \A[8][193] ;
wire   [4:0] \A[8][194] ;
wire   [4:0] \A[8][195] ;
wire   [4:0] \A[8][196] ;
wire   [4:0] \A[8][197] ;
wire   [4:0] \A[8][198] ;
wire   [4:0] \A[8][199] ;
wire   [4:0] \A[8][200] ;
wire   [4:0] \A[8][201] ;
wire   [4:0] \A[8][202] ;
wire   [4:0] \A[8][203] ;
wire   [4:0] \A[8][204] ;
wire   [4:0] \A[8][205] ;
wire   [4:0] \A[8][206] ;
wire   [4:0] \A[8][207] ;
wire   [4:0] \A[8][208] ;
wire   [4:0] \A[8][209] ;
wire   [4:0] \A[8][210] ;
wire   [4:0] \A[8][211] ;
wire   [4:0] \A[8][212] ;
wire   [4:0] \A[8][213] ;
wire   [4:0] \A[8][214] ;
wire   [4:0] \A[8][215] ;
wire   [4:0] \A[8][216] ;
wire   [4:0] \A[8][217] ;
wire   [4:0] \A[8][218] ;
wire   [4:0] \A[8][219] ;
wire   [4:0] \A[8][220] ;
wire   [4:0] \A[8][221] ;
wire   [4:0] \A[8][222] ;
wire   [4:0] \A[8][223] ;
wire   [4:0] \A[8][224] ;
wire   [4:0] \A[8][225] ;
wire   [4:0] \A[8][226] ;
wire   [4:0] \A[8][227] ;
wire   [4:0] \A[8][228] ;
wire   [4:0] \A[8][229] ;
wire   [4:0] \A[8][230] ;
wire   [4:0] \A[8][231] ;
wire   [4:0] \A[8][232] ;
wire   [4:0] \A[8][233] ;
wire   [4:0] \A[8][234] ;
wire   [4:0] \A[8][235] ;
wire   [4:0] \A[8][236] ;
wire   [4:0] \A[8][237] ;
wire   [4:0] \A[8][238] ;
wire   [4:0] \A[8][239] ;
wire   [4:0] \A[8][240] ;
wire   [4:0] \A[8][241] ;
wire   [4:0] \A[8][242] ;
wire   [4:0] \A[8][243] ;
wire   [4:0] \A[8][244] ;
wire   [4:0] \A[8][245] ;
wire   [4:0] \A[8][246] ;
wire   [4:0] \A[8][247] ;
wire   [4:0] \A[8][248] ;
wire   [4:0] \A[8][249] ;
wire   [4:0] \A[8][250] ;
wire   [4:0] \A[8][251] ;
wire   [4:0] \A[8][252] ;
wire   [4:0] \A[8][253] ;
wire   [4:0] \A[8][254] ;
wire   [4:0] \A[8][255] ;
wire   [4:0] \A[9][0] ;
wire   [4:0] \A[9][1] ;
wire   [4:0] \A[9][2] ;
wire   [4:0] \A[9][3] ;
wire   [4:0] \A[9][4] ;
wire   [4:0] \A[9][5] ;
wire   [4:0] \A[9][6] ;
wire   [4:0] \A[9][7] ;
wire   [4:0] \A[9][8] ;
wire   [4:0] \A[9][9] ;
wire   [4:0] \A[9][10] ;
wire   [4:0] \A[9][11] ;
wire   [4:0] \A[9][12] ;
wire   [4:0] \A[9][13] ;
wire   [4:0] \A[9][14] ;
wire   [4:0] \A[9][15] ;
wire   [4:0] \A[9][16] ;
wire   [4:0] \A[9][17] ;
wire   [4:0] \A[9][18] ;
wire   [4:0] \A[9][19] ;
wire   [4:0] \A[9][20] ;
wire   [4:0] \A[9][21] ;
wire   [4:0] \A[9][22] ;
wire   [4:0] \A[9][23] ;
wire   [4:0] \A[9][24] ;
wire   [4:0] \A[9][25] ;
wire   [4:0] \A[9][26] ;
wire   [4:0] \A[9][27] ;
wire   [4:0] \A[9][28] ;
wire   [4:0] \A[9][29] ;
wire   [4:0] \A[9][30] ;
wire   [4:0] \A[9][31] ;
wire   [4:0] \A[9][32] ;
wire   [4:0] \A[9][33] ;
wire   [4:0] \A[9][34] ;
wire   [4:0] \A[9][35] ;
wire   [4:0] \A[9][36] ;
wire   [4:0] \A[9][37] ;
wire   [4:0] \A[9][38] ;
wire   [4:0] \A[9][39] ;
wire   [4:0] \A[9][40] ;
wire   [4:0] \A[9][41] ;
wire   [4:0] \A[9][42] ;
wire   [4:0] \A[9][43] ;
wire   [4:0] \A[9][44] ;
wire   [4:0] \A[9][45] ;
wire   [4:0] \A[9][46] ;
wire   [4:0] \A[9][47] ;
wire   [4:0] \A[9][48] ;
wire   [4:0] \A[9][49] ;
wire   [4:0] \A[9][50] ;
wire   [4:0] \A[9][51] ;
wire   [4:0] \A[9][52] ;
wire   [4:0] \A[9][53] ;
wire   [4:0] \A[9][54] ;
wire   [4:0] \A[9][55] ;
wire   [4:0] \A[9][56] ;
wire   [4:0] \A[9][57] ;
wire   [4:0] \A[9][58] ;
wire   [4:0] \A[9][59] ;
wire   [4:0] \A[9][60] ;
wire   [4:0] \A[9][61] ;
wire   [4:0] \A[9][62] ;
wire   [4:0] \A[9][63] ;
wire   [4:0] \A[9][64] ;
wire   [4:0] \A[9][65] ;
wire   [4:0] \A[9][66] ;
wire   [4:0] \A[9][67] ;
wire   [4:0] \A[9][68] ;
wire   [4:0] \A[9][69] ;
wire   [4:0] \A[9][70] ;
wire   [4:0] \A[9][71] ;
wire   [4:0] \A[9][72] ;
wire   [4:0] \A[9][73] ;
wire   [4:0] \A[9][74] ;
wire   [4:0] \A[9][75] ;
wire   [4:0] \A[9][76] ;
wire   [4:0] \A[9][77] ;
wire   [4:0] \A[9][78] ;
wire   [4:0] \A[9][79] ;
wire   [4:0] \A[9][80] ;
wire   [4:0] \A[9][81] ;
wire   [4:0] \A[9][82] ;
wire   [4:0] \A[9][83] ;
wire   [4:0] \A[9][84] ;
wire   [4:0] \A[9][85] ;
wire   [4:0] \A[9][86] ;
wire   [4:0] \A[9][87] ;
wire   [4:0] \A[9][88] ;
wire   [4:0] \A[9][89] ;
wire   [4:0] \A[9][90] ;
wire   [4:0] \A[9][91] ;
wire   [4:0] \A[9][92] ;
wire   [4:0] \A[9][93] ;
wire   [4:0] \A[9][94] ;
wire   [4:0] \A[9][95] ;
wire   [4:0] \A[9][96] ;
wire   [4:0] \A[9][97] ;
wire   [4:0] \A[9][98] ;
wire   [4:0] \A[9][99] ;
wire   [4:0] \A[9][100] ;
wire   [4:0] \A[9][101] ;
wire   [4:0] \A[9][102] ;
wire   [4:0] \A[9][103] ;
wire   [4:0] \A[9][104] ;
wire   [4:0] \A[9][105] ;
wire   [4:0] \A[9][106] ;
wire   [4:0] \A[9][107] ;
wire   [4:0] \A[9][108] ;
wire   [4:0] \A[9][109] ;
wire   [4:0] \A[9][110] ;
wire   [4:0] \A[9][111] ;
wire   [4:0] \A[9][112] ;
wire   [4:0] \A[9][113] ;
wire   [4:0] \A[9][114] ;
wire   [4:0] \A[9][115] ;
wire   [4:0] \A[9][116] ;
wire   [4:0] \A[9][117] ;
wire   [4:0] \A[9][118] ;
wire   [4:0] \A[9][119] ;
wire   [4:0] \A[9][120] ;
wire   [4:0] \A[9][121] ;
wire   [4:0] \A[9][122] ;
wire   [4:0] \A[9][123] ;
wire   [4:0] \A[9][124] ;
wire   [4:0] \A[9][125] ;
wire   [4:0] \A[9][126] ;
wire   [4:0] \A[9][127] ;
wire   [4:0] \A[9][128] ;
wire   [4:0] \A[9][129] ;
wire   [4:0] \A[9][130] ;
wire   [4:0] \A[9][131] ;
wire   [4:0] \A[9][132] ;
wire   [4:0] \A[9][133] ;
wire   [4:0] \A[9][134] ;
wire   [4:0] \A[9][135] ;
wire   [4:0] \A[9][136] ;
wire   [4:0] \A[9][137] ;
wire   [4:0] \A[9][138] ;
wire   [4:0] \A[9][139] ;
wire   [4:0] \A[9][140] ;
wire   [4:0] \A[9][141] ;
wire   [4:0] \A[9][142] ;
wire   [4:0] \A[9][143] ;
wire   [4:0] \A[9][144] ;
wire   [4:0] \A[9][145] ;
wire   [4:0] \A[9][146] ;
wire   [4:0] \A[9][147] ;
wire   [4:0] \A[9][148] ;
wire   [4:0] \A[9][149] ;
wire   [4:0] \A[9][150] ;
wire   [4:0] \A[9][151] ;
wire   [4:0] \A[9][152] ;
wire   [4:0] \A[9][153] ;
wire   [4:0] \A[9][154] ;
wire   [4:0] \A[9][155] ;
wire   [4:0] \A[9][156] ;
wire   [4:0] \A[9][157] ;
wire   [4:0] \A[9][158] ;
wire   [4:0] \A[9][159] ;
wire   [4:0] \A[9][160] ;
wire   [4:0] \A[9][161] ;
wire   [4:0] \A[9][162] ;
wire   [4:0] \A[9][163] ;
wire   [4:0] \A[9][164] ;
wire   [4:0] \A[9][165] ;
wire   [4:0] \A[9][166] ;
wire   [4:0] \A[9][167] ;
wire   [4:0] \A[9][168] ;
wire   [4:0] \A[9][169] ;
wire   [4:0] \A[9][170] ;
wire   [4:0] \A[9][171] ;
wire   [4:0] \A[9][172] ;
wire   [4:0] \A[9][173] ;
wire   [4:0] \A[9][174] ;
wire   [4:0] \A[9][175] ;
wire   [4:0] \A[9][176] ;
wire   [4:0] \A[9][177] ;
wire   [4:0] \A[9][178] ;
wire   [4:0] \A[9][179] ;
wire   [4:0] \A[9][180] ;
wire   [4:0] \A[9][181] ;
wire   [4:0] \A[9][182] ;
wire   [4:0] \A[9][183] ;
wire   [4:0] \A[9][184] ;
wire   [4:0] \A[9][185] ;
wire   [4:0] \A[9][186] ;
wire   [4:0] \A[9][187] ;
wire   [4:0] \A[9][188] ;
wire   [4:0] \A[9][189] ;
wire   [4:0] \A[9][190] ;
wire   [4:0] \A[9][191] ;
wire   [4:0] \A[9][192] ;
wire   [4:0] \A[9][193] ;
wire   [4:0] \A[9][194] ;
wire   [4:0] \A[9][195] ;
wire   [4:0] \A[9][196] ;
wire   [4:0] \A[9][197] ;
wire   [4:0] \A[9][198] ;
wire   [4:0] \A[9][199] ;
wire   [4:0] \A[9][200] ;
wire   [4:0] \A[9][201] ;
wire   [4:0] \A[9][202] ;
wire   [4:0] \A[9][203] ;
wire   [4:0] \A[9][204] ;
wire   [4:0] \A[9][205] ;
wire   [4:0] \A[9][206] ;
wire   [4:0] \A[9][207] ;
wire   [4:0] \A[9][208] ;
wire   [4:0] \A[9][209] ;
wire   [4:0] \A[9][210] ;
wire   [4:0] \A[9][211] ;
wire   [4:0] \A[9][212] ;
wire   [4:0] \A[9][213] ;
wire   [4:0] \A[9][214] ;
wire   [4:0] \A[9][215] ;
wire   [4:0] \A[9][216] ;
wire   [4:0] \A[9][217] ;
wire   [4:0] \A[9][218] ;
wire   [4:0] \A[9][219] ;
wire   [4:0] \A[9][220] ;
wire   [4:0] \A[9][221] ;
wire   [4:0] \A[9][222] ;
wire   [4:0] \A[9][223] ;
wire   [4:0] \A[9][224] ;
wire   [4:0] \A[9][225] ;
wire   [4:0] \A[9][226] ;
wire   [4:0] \A[9][227] ;
wire   [4:0] \A[9][228] ;
wire   [4:0] \A[9][229] ;
wire   [4:0] \A[9][230] ;
wire   [4:0] \A[9][231] ;
wire   [4:0] \A[9][232] ;
wire   [4:0] \A[9][233] ;
wire   [4:0] \A[9][234] ;
wire   [4:0] \A[9][235] ;
wire   [4:0] \A[9][236] ;
wire   [4:0] \A[9][237] ;
wire   [4:0] \A[9][238] ;
wire   [4:0] \A[9][239] ;
wire   [4:0] \A[9][240] ;
wire   [4:0] \A[9][241] ;
wire   [4:0] \A[9][242] ;
wire   [4:0] \A[9][243] ;
wire   [4:0] \A[9][244] ;
wire   [4:0] \A[9][245] ;
wire   [4:0] \A[9][246] ;
wire   [4:0] \A[9][247] ;
wire   [4:0] \A[9][248] ;
wire   [4:0] \A[9][249] ;
wire   [4:0] \A[9][250] ;
wire   [4:0] \A[9][251] ;
wire   [4:0] \A[9][252] ;
wire   [4:0] \A[9][253] ;
wire   [4:0] \A[9][254] ;
wire   [4:0] \A[9][255] ;
wire   [4:0] \A[10][0] ;
wire   [4:0] \A[10][1] ;
wire   [4:0] \A[10][2] ;
wire   [4:0] \A[10][3] ;
wire   [4:0] \A[10][4] ;
wire   [4:0] \A[10][5] ;
wire   [4:0] \A[10][6] ;
wire   [4:0] \A[10][7] ;
wire   [4:0] \A[10][8] ;
wire   [4:0] \A[10][9] ;
wire   [4:0] \A[10][10] ;
wire   [4:0] \A[10][11] ;
wire   [4:0] \A[10][12] ;
wire   [4:0] \A[10][13] ;
wire   [4:0] \A[10][14] ;
wire   [4:0] \A[10][15] ;
wire   [4:0] \A[10][16] ;
wire   [4:0] \A[10][17] ;
wire   [4:0] \A[10][18] ;
wire   [4:0] \A[10][19] ;
wire   [4:0] \A[10][20] ;
wire   [4:0] \A[10][21] ;
wire   [4:0] \A[10][22] ;
wire   [4:0] \A[10][23] ;
wire   [4:0] \A[10][24] ;
wire   [4:0] \A[10][25] ;
wire   [4:0] \A[10][26] ;
wire   [4:0] \A[10][27] ;
wire   [4:0] \A[10][28] ;
wire   [4:0] \A[10][29] ;
wire   [4:0] \A[10][30] ;
wire   [4:0] \A[10][31] ;
wire   [4:0] \A[10][32] ;
wire   [4:0] \A[10][33] ;
wire   [4:0] \A[10][34] ;
wire   [4:0] \A[10][35] ;
wire   [4:0] \A[10][36] ;
wire   [4:0] \A[10][37] ;
wire   [4:0] \A[10][38] ;
wire   [4:0] \A[10][39] ;
wire   [4:0] \A[10][40] ;
wire   [4:0] \A[10][41] ;
wire   [4:0] \A[10][42] ;
wire   [4:0] \A[10][43] ;
wire   [4:0] \A[10][44] ;
wire   [4:0] \A[10][45] ;
wire   [4:0] \A[10][46] ;
wire   [4:0] \A[10][47] ;
wire   [4:0] \A[10][48] ;
wire   [4:0] \A[10][49] ;
wire   [4:0] \A[10][50] ;
wire   [4:0] \A[10][51] ;
wire   [4:0] \A[10][52] ;
wire   [4:0] \A[10][53] ;
wire   [4:0] \A[10][54] ;
wire   [4:0] \A[10][55] ;
wire   [4:0] \A[10][56] ;
wire   [4:0] \A[10][57] ;
wire   [4:0] \A[10][58] ;
wire   [4:0] \A[10][59] ;
wire   [4:0] \A[10][60] ;
wire   [4:0] \A[10][61] ;
wire   [4:0] \A[10][62] ;
wire   [4:0] \A[10][63] ;
wire   [4:0] \A[10][64] ;
wire   [4:0] \A[10][65] ;
wire   [4:0] \A[10][66] ;
wire   [4:0] \A[10][67] ;
wire   [4:0] \A[10][68] ;
wire   [4:0] \A[10][69] ;
wire   [4:0] \A[10][70] ;
wire   [4:0] \A[10][71] ;
wire   [4:0] \A[10][72] ;
wire   [4:0] \A[10][73] ;
wire   [4:0] \A[10][74] ;
wire   [4:0] \A[10][75] ;
wire   [4:0] \A[10][76] ;
wire   [4:0] \A[10][77] ;
wire   [4:0] \A[10][78] ;
wire   [4:0] \A[10][79] ;
wire   [4:0] \A[10][80] ;
wire   [4:0] \A[10][81] ;
wire   [4:0] \A[10][82] ;
wire   [4:0] \A[10][83] ;
wire   [4:0] \A[10][84] ;
wire   [4:0] \A[10][85] ;
wire   [4:0] \A[10][86] ;
wire   [4:0] \A[10][87] ;
wire   [4:0] \A[10][88] ;
wire   [4:0] \A[10][89] ;
wire   [4:0] \A[10][90] ;
wire   [4:0] \A[10][91] ;
wire   [4:0] \A[10][92] ;
wire   [4:0] \A[10][93] ;
wire   [4:0] \A[10][94] ;
wire   [4:0] \A[10][95] ;
wire   [4:0] \A[10][96] ;
wire   [4:0] \A[10][97] ;
wire   [4:0] \A[10][98] ;
wire   [4:0] \A[10][99] ;
wire   [4:0] \A[10][100] ;
wire   [4:0] \A[10][101] ;
wire   [4:0] \A[10][102] ;
wire   [4:0] \A[10][103] ;
wire   [4:0] \A[10][104] ;
wire   [4:0] \A[10][105] ;
wire   [4:0] \A[10][106] ;
wire   [4:0] \A[10][107] ;
wire   [4:0] \A[10][108] ;
wire   [4:0] \A[10][109] ;
wire   [4:0] \A[10][110] ;
wire   [4:0] \A[10][111] ;
wire   [4:0] \A[10][112] ;
wire   [4:0] \A[10][113] ;
wire   [4:0] \A[10][114] ;
wire   [4:0] \A[10][115] ;
wire   [4:0] \A[10][116] ;
wire   [4:0] \A[10][117] ;
wire   [4:0] \A[10][118] ;
wire   [4:0] \A[10][119] ;
wire   [4:0] \A[10][120] ;
wire   [4:0] \A[10][121] ;
wire   [4:0] \A[10][122] ;
wire   [4:0] \A[10][123] ;
wire   [4:0] \A[10][124] ;
wire   [4:0] \A[10][125] ;
wire   [4:0] \A[10][126] ;
wire   [4:0] \A[10][127] ;
wire   [4:0] \A[10][128] ;
wire   [4:0] \A[10][129] ;
wire   [4:0] \A[10][130] ;
wire   [4:0] \A[10][131] ;
wire   [4:0] \A[10][132] ;
wire   [4:0] \A[10][133] ;
wire   [4:0] \A[10][134] ;
wire   [4:0] \A[10][135] ;
wire   [4:0] \A[10][136] ;
wire   [4:0] \A[10][137] ;
wire   [4:0] \A[10][138] ;
wire   [4:0] \A[10][139] ;
wire   [4:0] \A[10][140] ;
wire   [4:0] \A[10][141] ;
wire   [4:0] \A[10][142] ;
wire   [4:0] \A[10][143] ;
wire   [4:0] \A[10][144] ;
wire   [4:0] \A[10][145] ;
wire   [4:0] \A[10][146] ;
wire   [4:0] \A[10][147] ;
wire   [4:0] \A[10][148] ;
wire   [4:0] \A[10][149] ;
wire   [4:0] \A[10][150] ;
wire   [4:0] \A[10][151] ;
wire   [4:0] \A[10][152] ;
wire   [4:0] \A[10][153] ;
wire   [4:0] \A[10][154] ;
wire   [4:0] \A[10][155] ;
wire   [4:0] \A[10][156] ;
wire   [4:0] \A[10][157] ;
wire   [4:0] \A[10][158] ;
wire   [4:0] \A[10][159] ;
wire   [4:0] \A[10][160] ;
wire   [4:0] \A[10][161] ;
wire   [4:0] \A[10][162] ;
wire   [4:0] \A[10][163] ;
wire   [4:0] \A[10][164] ;
wire   [4:0] \A[10][165] ;
wire   [4:0] \A[10][166] ;
wire   [4:0] \A[10][167] ;
wire   [4:0] \A[10][168] ;
wire   [4:0] \A[10][169] ;
wire   [4:0] \A[10][170] ;
wire   [4:0] \A[10][171] ;
wire   [4:0] \A[10][172] ;
wire   [4:0] \A[10][173] ;
wire   [4:0] \A[10][174] ;
wire   [4:0] \A[10][175] ;
wire   [4:0] \A[10][176] ;
wire   [4:0] \A[10][177] ;
wire   [4:0] \A[10][178] ;
wire   [4:0] \A[10][179] ;
wire   [4:0] \A[10][180] ;
wire   [4:0] \A[10][181] ;
wire   [4:0] \A[10][182] ;
wire   [4:0] \A[10][183] ;
wire   [4:0] \A[10][184] ;
wire   [4:0] \A[10][185] ;
wire   [4:0] \A[10][186] ;
wire   [4:0] \A[10][187] ;
wire   [4:0] \A[10][188] ;
wire   [4:0] \A[10][189] ;
wire   [4:0] \A[10][190] ;
wire   [4:0] \A[10][191] ;
wire   [4:0] \A[10][192] ;
wire   [4:0] \A[10][193] ;
wire   [4:0] \A[10][194] ;
wire   [4:0] \A[10][195] ;
wire   [4:0] \A[10][196] ;
wire   [4:0] \A[10][197] ;
wire   [4:0] \A[10][198] ;
wire   [4:0] \A[10][199] ;
wire   [4:0] \A[10][200] ;
wire   [4:0] \A[10][201] ;
wire   [4:0] \A[10][202] ;
wire   [4:0] \A[10][203] ;
wire   [4:0] \A[10][204] ;
wire   [4:0] \A[10][205] ;
wire   [4:0] \A[10][206] ;
wire   [4:0] \A[10][207] ;
wire   [4:0] \A[10][208] ;
wire   [4:0] \A[10][209] ;
wire   [4:0] \A[10][210] ;
wire   [4:0] \A[10][211] ;
wire   [4:0] \A[10][212] ;
wire   [4:0] \A[10][213] ;
wire   [4:0] \A[10][214] ;
wire   [4:0] \A[10][215] ;
wire   [4:0] \A[10][216] ;
wire   [4:0] \A[10][217] ;
wire   [4:0] \A[10][218] ;
wire   [4:0] \A[10][219] ;
wire   [4:0] \A[10][220] ;
wire   [4:0] \A[10][221] ;
wire   [4:0] \A[10][222] ;
wire   [4:0] \A[10][223] ;
wire   [4:0] \A[10][224] ;
wire   [4:0] \A[10][225] ;
wire   [4:0] \A[10][226] ;
wire   [4:0] \A[10][227] ;
wire   [4:0] \A[10][228] ;
wire   [4:0] \A[10][229] ;
wire   [4:0] \A[10][230] ;
wire   [4:0] \A[10][231] ;
wire   [4:0] \A[10][232] ;
wire   [4:0] \A[10][233] ;
wire   [4:0] \A[10][234] ;
wire   [4:0] \A[10][235] ;
wire   [4:0] \A[10][236] ;
wire   [4:0] \A[10][237] ;
wire   [4:0] \A[10][238] ;
wire   [4:0] \A[10][239] ;
wire   [4:0] \A[10][240] ;
wire   [4:0] \A[10][241] ;
wire   [4:0] \A[10][242] ;
wire   [4:0] \A[10][243] ;
wire   [4:0] \A[10][244] ;
wire   [4:0] \A[10][245] ;
wire   [4:0] \A[10][246] ;
wire   [4:0] \A[10][247] ;
wire   [4:0] \A[10][248] ;
wire   [4:0] \A[10][249] ;
wire   [4:0] \A[10][250] ;
wire   [4:0] \A[10][251] ;
wire   [4:0] \A[10][252] ;
wire   [4:0] \A[10][253] ;
wire   [4:0] \A[10][254] ;
wire   [4:0] \A[10][255] ;
wire   [4:0] \A[11][0] ;
wire   [4:0] \A[11][1] ;
wire   [4:0] \A[11][2] ;
wire   [4:0] \A[11][3] ;
wire   [4:0] \A[11][4] ;
wire   [4:0] \A[11][5] ;
wire   [4:0] \A[11][6] ;
wire   [4:0] \A[11][7] ;
wire   [4:0] \A[11][8] ;
wire   [4:0] \A[11][9] ;
wire   [4:0] \A[11][10] ;
wire   [4:0] \A[11][11] ;
wire   [4:0] \A[11][12] ;
wire   [4:0] \A[11][13] ;
wire   [4:0] \A[11][14] ;
wire   [4:0] \A[11][15] ;
wire   [4:0] \A[11][16] ;
wire   [4:0] \A[11][17] ;
wire   [4:0] \A[11][18] ;
wire   [4:0] \A[11][19] ;
wire   [4:0] \A[11][20] ;
wire   [4:0] \A[11][21] ;
wire   [4:0] \A[11][22] ;
wire   [4:0] \A[11][23] ;
wire   [4:0] \A[11][24] ;
wire   [4:0] \A[11][25] ;
wire   [4:0] \A[11][26] ;
wire   [4:0] \A[11][27] ;
wire   [4:0] \A[11][28] ;
wire   [4:0] \A[11][29] ;
wire   [4:0] \A[11][30] ;
wire   [4:0] \A[11][31] ;
wire   [4:0] \A[11][32] ;
wire   [4:0] \A[11][33] ;
wire   [4:0] \A[11][34] ;
wire   [4:0] \A[11][35] ;
wire   [4:0] \A[11][36] ;
wire   [4:0] \A[11][37] ;
wire   [4:0] \A[11][38] ;
wire   [4:0] \A[11][39] ;
wire   [4:0] \A[11][40] ;
wire   [4:0] \A[11][41] ;
wire   [4:0] \A[11][42] ;
wire   [4:0] \A[11][43] ;
wire   [4:0] \A[11][44] ;
wire   [4:0] \A[11][45] ;
wire   [4:0] \A[11][46] ;
wire   [4:0] \A[11][47] ;
wire   [4:0] \A[11][48] ;
wire   [4:0] \A[11][49] ;
wire   [4:0] \A[11][50] ;
wire   [4:0] \A[11][51] ;
wire   [4:0] \A[11][52] ;
wire   [4:0] \A[11][53] ;
wire   [4:0] \A[11][54] ;
wire   [4:0] \A[11][55] ;
wire   [4:0] \A[11][56] ;
wire   [4:0] \A[11][57] ;
wire   [4:0] \A[11][58] ;
wire   [4:0] \A[11][59] ;
wire   [4:0] \A[11][60] ;
wire   [4:0] \A[11][61] ;
wire   [4:0] \A[11][62] ;
wire   [4:0] \A[11][63] ;
wire   [4:0] \A[11][64] ;
wire   [4:0] \A[11][65] ;
wire   [4:0] \A[11][66] ;
wire   [4:0] \A[11][67] ;
wire   [4:0] \A[11][68] ;
wire   [4:0] \A[11][69] ;
wire   [4:0] \A[11][70] ;
wire   [4:0] \A[11][71] ;
wire   [4:0] \A[11][72] ;
wire   [4:0] \A[11][73] ;
wire   [4:0] \A[11][74] ;
wire   [4:0] \A[11][75] ;
wire   [4:0] \A[11][76] ;
wire   [4:0] \A[11][77] ;
wire   [4:0] \A[11][78] ;
wire   [4:0] \A[11][79] ;
wire   [4:0] \A[11][80] ;
wire   [4:0] \A[11][81] ;
wire   [4:0] \A[11][82] ;
wire   [4:0] \A[11][83] ;
wire   [4:0] \A[11][84] ;
wire   [4:0] \A[11][85] ;
wire   [4:0] \A[11][86] ;
wire   [4:0] \A[11][87] ;
wire   [4:0] \A[11][88] ;
wire   [4:0] \A[11][89] ;
wire   [4:0] \A[11][90] ;
wire   [4:0] \A[11][91] ;
wire   [4:0] \A[11][92] ;
wire   [4:0] \A[11][93] ;
wire   [4:0] \A[11][94] ;
wire   [4:0] \A[11][95] ;
wire   [4:0] \A[11][96] ;
wire   [4:0] \A[11][97] ;
wire   [4:0] \A[11][98] ;
wire   [4:0] \A[11][99] ;
wire   [4:0] \A[11][100] ;
wire   [4:0] \A[11][101] ;
wire   [4:0] \A[11][102] ;
wire   [4:0] \A[11][103] ;
wire   [4:0] \A[11][104] ;
wire   [4:0] \A[11][105] ;
wire   [4:0] \A[11][106] ;
wire   [4:0] \A[11][107] ;
wire   [4:0] \A[11][108] ;
wire   [4:0] \A[11][109] ;
wire   [4:0] \A[11][110] ;
wire   [4:0] \A[11][111] ;
wire   [4:0] \A[11][112] ;
wire   [4:0] \A[11][113] ;
wire   [4:0] \A[11][114] ;
wire   [4:0] \A[11][115] ;
wire   [4:0] \A[11][116] ;
wire   [4:0] \A[11][117] ;
wire   [4:0] \A[11][118] ;
wire   [4:0] \A[11][119] ;
wire   [4:0] \A[11][120] ;
wire   [4:0] \A[11][121] ;
wire   [4:0] \A[11][122] ;
wire   [4:0] \A[11][123] ;
wire   [4:0] \A[11][124] ;
wire   [4:0] \A[11][125] ;
wire   [4:0] \A[11][126] ;
wire   [4:0] \A[11][127] ;
wire   [4:0] \A[11][128] ;
wire   [4:0] \A[11][129] ;
wire   [4:0] \A[11][130] ;
wire   [4:0] \A[11][131] ;
wire   [4:0] \A[11][132] ;
wire   [4:0] \A[11][133] ;
wire   [4:0] \A[11][134] ;
wire   [4:0] \A[11][135] ;
wire   [4:0] \A[11][136] ;
wire   [4:0] \A[11][137] ;
wire   [4:0] \A[11][138] ;
wire   [4:0] \A[11][139] ;
wire   [4:0] \A[11][140] ;
wire   [4:0] \A[11][141] ;
wire   [4:0] \A[11][142] ;
wire   [4:0] \A[11][143] ;
wire   [4:0] \A[11][144] ;
wire   [4:0] \A[11][145] ;
wire   [4:0] \A[11][146] ;
wire   [4:0] \A[11][147] ;
wire   [4:0] \A[11][148] ;
wire   [4:0] \A[11][149] ;
wire   [4:0] \A[11][150] ;
wire   [4:0] \A[11][151] ;
wire   [4:0] \A[11][152] ;
wire   [4:0] \A[11][153] ;
wire   [4:0] \A[11][154] ;
wire   [4:0] \A[11][155] ;
wire   [4:0] \A[11][156] ;
wire   [4:0] \A[11][157] ;
wire   [4:0] \A[11][158] ;
wire   [4:0] \A[11][159] ;
wire   [4:0] \A[11][160] ;
wire   [4:0] \A[11][161] ;
wire   [4:0] \A[11][162] ;
wire   [4:0] \A[11][163] ;
wire   [4:0] \A[11][164] ;
wire   [4:0] \A[11][165] ;
wire   [4:0] \A[11][166] ;
wire   [4:0] \A[11][167] ;
wire   [4:0] \A[11][168] ;
wire   [4:0] \A[11][169] ;
wire   [4:0] \A[11][170] ;
wire   [4:0] \A[11][171] ;
wire   [4:0] \A[11][172] ;
wire   [4:0] \A[11][173] ;
wire   [4:0] \A[11][174] ;
wire   [4:0] \A[11][175] ;
wire   [4:0] \A[11][176] ;
wire   [4:0] \A[11][177] ;
wire   [4:0] \A[11][178] ;
wire   [4:0] \A[11][179] ;
wire   [4:0] \A[11][180] ;
wire   [4:0] \A[11][181] ;
wire   [4:0] \A[11][182] ;
wire   [4:0] \A[11][183] ;
wire   [4:0] \A[11][184] ;
wire   [4:0] \A[11][185] ;
wire   [4:0] \A[11][186] ;
wire   [4:0] \A[11][187] ;
wire   [4:0] \A[11][188] ;
wire   [4:0] \A[11][189] ;
wire   [4:0] \A[11][190] ;
wire   [4:0] \A[11][191] ;
wire   [4:0] \A[11][192] ;
wire   [4:0] \A[11][193] ;
wire   [4:0] \A[11][194] ;
wire   [4:0] \A[11][195] ;
wire   [4:0] \A[11][196] ;
wire   [4:0] \A[11][197] ;
wire   [4:0] \A[11][198] ;
wire   [4:0] \A[11][199] ;
wire   [4:0] \A[11][200] ;
wire   [4:0] \A[11][201] ;
wire   [4:0] \A[11][202] ;
wire   [4:0] \A[11][203] ;
wire   [4:0] \A[11][204] ;
wire   [4:0] \A[11][205] ;
wire   [4:0] \A[11][206] ;
wire   [4:0] \A[11][207] ;
wire   [4:0] \A[11][208] ;
wire   [4:0] \A[11][209] ;
wire   [4:0] \A[11][210] ;
wire   [4:0] \A[11][211] ;
wire   [4:0] \A[11][212] ;
wire   [4:0] \A[11][213] ;
wire   [4:0] \A[11][214] ;
wire   [4:0] \A[11][215] ;
wire   [4:0] \A[11][216] ;
wire   [4:0] \A[11][217] ;
wire   [4:0] \A[11][218] ;
wire   [4:0] \A[11][219] ;
wire   [4:0] \A[11][220] ;
wire   [4:0] \A[11][221] ;
wire   [4:0] \A[11][222] ;
wire   [4:0] \A[11][223] ;
wire   [4:0] \A[11][224] ;
wire   [4:0] \A[11][225] ;
wire   [4:0] \A[11][226] ;
wire   [4:0] \A[11][227] ;
wire   [4:0] \A[11][228] ;
wire   [4:0] \A[11][229] ;
wire   [4:0] \A[11][230] ;
wire   [4:0] \A[11][231] ;
wire   [4:0] \A[11][232] ;
wire   [4:0] \A[11][233] ;
wire   [4:0] \A[11][234] ;
wire   [4:0] \A[11][235] ;
wire   [4:0] \A[11][236] ;
wire   [4:0] \A[11][237] ;
wire   [4:0] \A[11][238] ;
wire   [4:0] \A[11][239] ;
wire   [4:0] \A[11][240] ;
wire   [4:0] \A[11][241] ;
wire   [4:0] \A[11][242] ;
wire   [4:0] \A[11][243] ;
wire   [4:0] \A[11][244] ;
wire   [4:0] \A[11][245] ;
wire   [4:0] \A[11][246] ;
wire   [4:0] \A[11][247] ;
wire   [4:0] \A[11][248] ;
wire   [4:0] \A[11][249] ;
wire   [4:0] \A[11][250] ;
wire   [4:0] \A[11][251] ;
wire   [4:0] \A[11][252] ;
wire   [4:0] \A[11][253] ;
wire   [4:0] \A[11][254] ;
wire   [4:0] \A[11][255] ;
wire   [4:0] \A[12][0] ;
wire   [4:0] \A[12][1] ;
wire   [4:0] \A[12][2] ;
wire   [4:0] \A[12][3] ;
wire   [4:0] \A[12][4] ;
wire   [4:0] \A[12][5] ;
wire   [4:0] \A[12][6] ;
wire   [4:0] \A[12][7] ;
wire   [4:0] \A[12][8] ;
wire   [4:0] \A[12][9] ;
wire   [4:0] \A[12][10] ;
wire   [4:0] \A[12][11] ;
wire   [4:0] \A[12][12] ;
wire   [4:0] \A[12][13] ;
wire   [4:0] \A[12][14] ;
wire   [4:0] \A[12][15] ;
wire   [4:0] \A[12][16] ;
wire   [4:0] \A[12][17] ;
wire   [4:0] \A[12][18] ;
wire   [4:0] \A[12][19] ;
wire   [4:0] \A[12][20] ;
wire   [4:0] \A[12][21] ;
wire   [4:0] \A[12][22] ;
wire   [4:0] \A[12][23] ;
wire   [4:0] \A[12][24] ;
wire   [4:0] \A[12][25] ;
wire   [4:0] \A[12][26] ;
wire   [4:0] \A[12][27] ;
wire   [4:0] \A[12][28] ;
wire   [4:0] \A[12][29] ;
wire   [4:0] \A[12][30] ;
wire   [4:0] \A[12][31] ;
wire   [4:0] \A[12][32] ;
wire   [4:0] \A[12][33] ;
wire   [4:0] \A[12][34] ;
wire   [4:0] \A[12][35] ;
wire   [4:0] \A[12][36] ;
wire   [4:0] \A[12][37] ;
wire   [4:0] \A[12][38] ;
wire   [4:0] \A[12][39] ;
wire   [4:0] \A[12][40] ;
wire   [4:0] \A[12][41] ;
wire   [4:0] \A[12][42] ;
wire   [4:0] \A[12][43] ;
wire   [4:0] \A[12][44] ;
wire   [4:0] \A[12][45] ;
wire   [4:0] \A[12][46] ;
wire   [4:0] \A[12][47] ;
wire   [4:0] \A[12][48] ;
wire   [4:0] \A[12][49] ;
wire   [4:0] \A[12][50] ;
wire   [4:0] \A[12][51] ;
wire   [4:0] \A[12][52] ;
wire   [4:0] \A[12][53] ;
wire   [4:0] \A[12][54] ;
wire   [4:0] \A[12][55] ;
wire   [4:0] \A[12][56] ;
wire   [4:0] \A[12][57] ;
wire   [4:0] \A[12][58] ;
wire   [4:0] \A[12][59] ;
wire   [4:0] \A[12][60] ;
wire   [4:0] \A[12][61] ;
wire   [4:0] \A[12][62] ;
wire   [4:0] \A[12][63] ;
wire   [4:0] \A[12][64] ;
wire   [4:0] \A[12][65] ;
wire   [4:0] \A[12][66] ;
wire   [4:0] \A[12][67] ;
wire   [4:0] \A[12][68] ;
wire   [4:0] \A[12][69] ;
wire   [4:0] \A[12][70] ;
wire   [4:0] \A[12][71] ;
wire   [4:0] \A[12][72] ;
wire   [4:0] \A[12][73] ;
wire   [4:0] \A[12][74] ;
wire   [4:0] \A[12][75] ;
wire   [4:0] \A[12][76] ;
wire   [4:0] \A[12][77] ;
wire   [4:0] \A[12][78] ;
wire   [4:0] \A[12][79] ;
wire   [4:0] \A[12][80] ;
wire   [4:0] \A[12][81] ;
wire   [4:0] \A[12][82] ;
wire   [4:0] \A[12][83] ;
wire   [4:0] \A[12][84] ;
wire   [4:0] \A[12][85] ;
wire   [4:0] \A[12][86] ;
wire   [4:0] \A[12][87] ;
wire   [4:0] \A[12][88] ;
wire   [4:0] \A[12][89] ;
wire   [4:0] \A[12][90] ;
wire   [4:0] \A[12][91] ;
wire   [4:0] \A[12][92] ;
wire   [4:0] \A[12][93] ;
wire   [4:0] \A[12][94] ;
wire   [4:0] \A[12][95] ;
wire   [4:0] \A[12][96] ;
wire   [4:0] \A[12][97] ;
wire   [4:0] \A[12][98] ;
wire   [4:0] \A[12][99] ;
wire   [4:0] \A[12][100] ;
wire   [4:0] \A[12][101] ;
wire   [4:0] \A[12][102] ;
wire   [4:0] \A[12][103] ;
wire   [4:0] \A[12][104] ;
wire   [4:0] \A[12][105] ;
wire   [4:0] \A[12][106] ;
wire   [4:0] \A[12][107] ;
wire   [4:0] \A[12][108] ;
wire   [4:0] \A[12][109] ;
wire   [4:0] \A[12][110] ;
wire   [4:0] \A[12][111] ;
wire   [4:0] \A[12][112] ;
wire   [4:0] \A[12][113] ;
wire   [4:0] \A[12][114] ;
wire   [4:0] \A[12][115] ;
wire   [4:0] \A[12][116] ;
wire   [4:0] \A[12][117] ;
wire   [4:0] \A[12][118] ;
wire   [4:0] \A[12][119] ;
wire   [4:0] \A[12][120] ;
wire   [4:0] \A[12][121] ;
wire   [4:0] \A[12][122] ;
wire   [4:0] \A[12][123] ;
wire   [4:0] \A[12][124] ;
wire   [4:0] \A[12][125] ;
wire   [4:0] \A[12][126] ;
wire   [4:0] \A[12][127] ;
wire   [4:0] \A[12][128] ;
wire   [4:0] \A[12][129] ;
wire   [4:0] \A[12][130] ;
wire   [4:0] \A[12][131] ;
wire   [4:0] \A[12][132] ;
wire   [4:0] \A[12][133] ;
wire   [4:0] \A[12][134] ;
wire   [4:0] \A[12][135] ;
wire   [4:0] \A[12][136] ;
wire   [4:0] \A[12][137] ;
wire   [4:0] \A[12][138] ;
wire   [4:0] \A[12][139] ;
wire   [4:0] \A[12][140] ;
wire   [4:0] \A[12][141] ;
wire   [4:0] \A[12][142] ;
wire   [4:0] \A[12][143] ;
wire   [4:0] \A[12][144] ;
wire   [4:0] \A[12][145] ;
wire   [4:0] \A[12][146] ;
wire   [4:0] \A[12][147] ;
wire   [4:0] \A[12][148] ;
wire   [4:0] \A[12][149] ;
wire   [4:0] \A[12][150] ;
wire   [4:0] \A[12][151] ;
wire   [4:0] \A[12][152] ;
wire   [4:0] \A[12][153] ;
wire   [4:0] \A[12][154] ;
wire   [4:0] \A[12][155] ;
wire   [4:0] \A[12][156] ;
wire   [4:0] \A[12][157] ;
wire   [4:0] \A[12][158] ;
wire   [4:0] \A[12][159] ;
wire   [4:0] \A[12][160] ;
wire   [4:0] \A[12][161] ;
wire   [4:0] \A[12][162] ;
wire   [4:0] \A[12][163] ;
wire   [4:0] \A[12][164] ;
wire   [4:0] \A[12][165] ;
wire   [4:0] \A[12][166] ;
wire   [4:0] \A[12][167] ;
wire   [4:0] \A[12][168] ;
wire   [4:0] \A[12][169] ;
wire   [4:0] \A[12][170] ;
wire   [4:0] \A[12][171] ;
wire   [4:0] \A[12][172] ;
wire   [4:0] \A[12][173] ;
wire   [4:0] \A[12][174] ;
wire   [4:0] \A[12][175] ;
wire   [4:0] \A[12][176] ;
wire   [4:0] \A[12][177] ;
wire   [4:0] \A[12][178] ;
wire   [4:0] \A[12][179] ;
wire   [4:0] \A[12][180] ;
wire   [4:0] \A[12][181] ;
wire   [4:0] \A[12][182] ;
wire   [4:0] \A[12][183] ;
wire   [4:0] \A[12][184] ;
wire   [4:0] \A[12][185] ;
wire   [4:0] \A[12][186] ;
wire   [4:0] \A[12][187] ;
wire   [4:0] \A[12][188] ;
wire   [4:0] \A[12][189] ;
wire   [4:0] \A[12][190] ;
wire   [4:0] \A[12][191] ;
wire   [4:0] \A[12][192] ;
wire   [4:0] \A[12][193] ;
wire   [4:0] \A[12][194] ;
wire   [4:0] \A[12][195] ;
wire   [4:0] \A[12][196] ;
wire   [4:0] \A[12][197] ;
wire   [4:0] \A[12][198] ;
wire   [4:0] \A[12][199] ;
wire   [4:0] \A[12][200] ;
wire   [4:0] \A[12][201] ;
wire   [4:0] \A[12][202] ;
wire   [4:0] \A[12][203] ;
wire   [4:0] \A[12][204] ;
wire   [4:0] \A[12][205] ;
wire   [4:0] \A[12][206] ;
wire   [4:0] \A[12][207] ;
wire   [4:0] \A[12][208] ;
wire   [4:0] \A[12][209] ;
wire   [4:0] \A[12][210] ;
wire   [4:0] \A[12][211] ;
wire   [4:0] \A[12][212] ;
wire   [4:0] \A[12][213] ;
wire   [4:0] \A[12][214] ;
wire   [4:0] \A[12][215] ;
wire   [4:0] \A[12][216] ;
wire   [4:0] \A[12][217] ;
wire   [4:0] \A[12][218] ;
wire   [4:0] \A[12][219] ;
wire   [4:0] \A[12][220] ;
wire   [4:0] \A[12][221] ;
wire   [4:0] \A[12][222] ;
wire   [4:0] \A[12][223] ;
wire   [4:0] \A[12][224] ;
wire   [4:0] \A[12][225] ;
wire   [4:0] \A[12][226] ;
wire   [4:0] \A[12][227] ;
wire   [4:0] \A[12][228] ;
wire   [4:0] \A[12][229] ;
wire   [4:0] \A[12][230] ;
wire   [4:0] \A[12][231] ;
wire   [4:0] \A[12][232] ;
wire   [4:0] \A[12][233] ;
wire   [4:0] \A[12][234] ;
wire   [4:0] \A[12][235] ;
wire   [4:0] \A[12][236] ;
wire   [4:0] \A[12][237] ;
wire   [4:0] \A[12][238] ;
wire   [4:0] \A[12][239] ;
wire   [4:0] \A[12][240] ;
wire   [4:0] \A[12][241] ;
wire   [4:0] \A[12][242] ;
wire   [4:0] \A[12][243] ;
wire   [4:0] \A[12][244] ;
wire   [4:0] \A[12][245] ;
wire   [4:0] \A[12][246] ;
wire   [4:0] \A[12][247] ;
wire   [4:0] \A[12][248] ;
wire   [4:0] \A[12][249] ;
wire   [4:0] \A[12][250] ;
wire   [4:0] \A[12][251] ;
wire   [4:0] \A[12][252] ;
wire   [4:0] \A[12][253] ;
wire   [4:0] \A[12][254] ;
wire   [4:0] \A[12][255] ;
wire   [4:0] \A[13][0] ;
wire   [4:0] \A[13][1] ;
wire   [4:0] \A[13][2] ;
wire   [4:0] \A[13][3] ;
wire   [4:0] \A[13][4] ;
wire   [4:0] \A[13][5] ;
wire   [4:0] \A[13][6] ;
wire   [4:0] \A[13][7] ;
wire   [4:0] \A[13][8] ;
wire   [4:0] \A[13][9] ;
wire   [4:0] \A[13][10] ;
wire   [4:0] \A[13][11] ;
wire   [4:0] \A[13][12] ;
wire   [4:0] \A[13][13] ;
wire   [4:0] \A[13][14] ;
wire   [4:0] \A[13][15] ;
wire   [4:0] \A[13][16] ;
wire   [4:0] \A[13][17] ;
wire   [4:0] \A[13][18] ;
wire   [4:0] \A[13][19] ;
wire   [4:0] \A[13][20] ;
wire   [4:0] \A[13][21] ;
wire   [4:0] \A[13][22] ;
wire   [4:0] \A[13][23] ;
wire   [4:0] \A[13][24] ;
wire   [4:0] \A[13][25] ;
wire   [4:0] \A[13][26] ;
wire   [4:0] \A[13][27] ;
wire   [4:0] \A[13][28] ;
wire   [4:0] \A[13][29] ;
wire   [4:0] \A[13][30] ;
wire   [4:0] \A[13][31] ;
wire   [4:0] \A[13][32] ;
wire   [4:0] \A[13][33] ;
wire   [4:0] \A[13][34] ;
wire   [4:0] \A[13][35] ;
wire   [4:0] \A[13][36] ;
wire   [4:0] \A[13][37] ;
wire   [4:0] \A[13][38] ;
wire   [4:0] \A[13][39] ;
wire   [4:0] \A[13][40] ;
wire   [4:0] \A[13][41] ;
wire   [4:0] \A[13][42] ;
wire   [4:0] \A[13][43] ;
wire   [4:0] \A[13][44] ;
wire   [4:0] \A[13][45] ;
wire   [4:0] \A[13][46] ;
wire   [4:0] \A[13][47] ;
wire   [4:0] \A[13][48] ;
wire   [4:0] \A[13][49] ;
wire   [4:0] \A[13][50] ;
wire   [4:0] \A[13][51] ;
wire   [4:0] \A[13][52] ;
wire   [4:0] \A[13][53] ;
wire   [4:0] \A[13][54] ;
wire   [4:0] \A[13][55] ;
wire   [4:0] \A[13][56] ;
wire   [4:0] \A[13][57] ;
wire   [4:0] \A[13][58] ;
wire   [4:0] \A[13][59] ;
wire   [4:0] \A[13][60] ;
wire   [4:0] \A[13][61] ;
wire   [4:0] \A[13][62] ;
wire   [4:0] \A[13][63] ;
wire   [4:0] \A[13][64] ;
wire   [4:0] \A[13][65] ;
wire   [4:0] \A[13][66] ;
wire   [4:0] \A[13][67] ;
wire   [4:0] \A[13][68] ;
wire   [4:0] \A[13][69] ;
wire   [4:0] \A[13][70] ;
wire   [4:0] \A[13][71] ;
wire   [4:0] \A[13][72] ;
wire   [4:0] \A[13][73] ;
wire   [4:0] \A[13][74] ;
wire   [4:0] \A[13][75] ;
wire   [4:0] \A[13][76] ;
wire   [4:0] \A[13][77] ;
wire   [4:0] \A[13][78] ;
wire   [4:0] \A[13][79] ;
wire   [4:0] \A[13][80] ;
wire   [4:0] \A[13][81] ;
wire   [4:0] \A[13][82] ;
wire   [4:0] \A[13][83] ;
wire   [4:0] \A[13][84] ;
wire   [4:0] \A[13][85] ;
wire   [4:0] \A[13][86] ;
wire   [4:0] \A[13][87] ;
wire   [4:0] \A[13][88] ;
wire   [4:0] \A[13][89] ;
wire   [4:0] \A[13][90] ;
wire   [4:0] \A[13][91] ;
wire   [4:0] \A[13][92] ;
wire   [4:0] \A[13][93] ;
wire   [4:0] \A[13][94] ;
wire   [4:0] \A[13][95] ;
wire   [4:0] \A[13][96] ;
wire   [4:0] \A[13][97] ;
wire   [4:0] \A[13][98] ;
wire   [4:0] \A[13][99] ;
wire   [4:0] \A[13][100] ;
wire   [4:0] \A[13][101] ;
wire   [4:0] \A[13][102] ;
wire   [4:0] \A[13][103] ;
wire   [4:0] \A[13][104] ;
wire   [4:0] \A[13][105] ;
wire   [4:0] \A[13][106] ;
wire   [4:0] \A[13][107] ;
wire   [4:0] \A[13][108] ;
wire   [4:0] \A[13][109] ;
wire   [4:0] \A[13][110] ;
wire   [4:0] \A[13][111] ;
wire   [4:0] \A[13][112] ;
wire   [4:0] \A[13][113] ;
wire   [4:0] \A[13][114] ;
wire   [4:0] \A[13][115] ;
wire   [4:0] \A[13][116] ;
wire   [4:0] \A[13][117] ;
wire   [4:0] \A[13][118] ;
wire   [4:0] \A[13][119] ;
wire   [4:0] \A[13][120] ;
wire   [4:0] \A[13][121] ;
wire   [4:0] \A[13][122] ;
wire   [4:0] \A[13][123] ;
wire   [4:0] \A[13][124] ;
wire   [4:0] \A[13][125] ;
wire   [4:0] \A[13][126] ;
wire   [4:0] \A[13][127] ;
wire   [4:0] \A[13][128] ;
wire   [4:0] \A[13][129] ;
wire   [4:0] \A[13][130] ;
wire   [4:0] \A[13][131] ;
wire   [4:0] \A[13][132] ;
wire   [4:0] \A[13][133] ;
wire   [4:0] \A[13][134] ;
wire   [4:0] \A[13][135] ;
wire   [4:0] \A[13][136] ;
wire   [4:0] \A[13][137] ;
wire   [4:0] \A[13][138] ;
wire   [4:0] \A[13][139] ;
wire   [4:0] \A[13][140] ;
wire   [4:0] \A[13][141] ;
wire   [4:0] \A[13][142] ;
wire   [4:0] \A[13][143] ;
wire   [4:0] \A[13][144] ;
wire   [4:0] \A[13][145] ;
wire   [4:0] \A[13][146] ;
wire   [4:0] \A[13][147] ;
wire   [4:0] \A[13][148] ;
wire   [4:0] \A[13][149] ;
wire   [4:0] \A[13][150] ;
wire   [4:0] \A[13][151] ;
wire   [4:0] \A[13][152] ;
wire   [4:0] \A[13][153] ;
wire   [4:0] \A[13][154] ;
wire   [4:0] \A[13][155] ;
wire   [4:0] \A[13][156] ;
wire   [4:0] \A[13][157] ;
wire   [4:0] \A[13][158] ;
wire   [4:0] \A[13][159] ;
wire   [4:0] \A[13][160] ;
wire   [4:0] \A[13][161] ;
wire   [4:0] \A[13][162] ;
wire   [4:0] \A[13][163] ;
wire   [4:0] \A[13][164] ;
wire   [4:0] \A[13][165] ;
wire   [4:0] \A[13][166] ;
wire   [4:0] \A[13][167] ;
wire   [4:0] \A[13][168] ;
wire   [4:0] \A[13][169] ;
wire   [4:0] \A[13][170] ;
wire   [4:0] \A[13][171] ;
wire   [4:0] \A[13][172] ;
wire   [4:0] \A[13][173] ;
wire   [4:0] \A[13][174] ;
wire   [4:0] \A[13][175] ;
wire   [4:0] \A[13][176] ;
wire   [4:0] \A[13][177] ;
wire   [4:0] \A[13][178] ;
wire   [4:0] \A[13][179] ;
wire   [4:0] \A[13][180] ;
wire   [4:0] \A[13][181] ;
wire   [4:0] \A[13][182] ;
wire   [4:0] \A[13][183] ;
wire   [4:0] \A[13][184] ;
wire   [4:0] \A[13][185] ;
wire   [4:0] \A[13][186] ;
wire   [4:0] \A[13][187] ;
wire   [4:0] \A[13][188] ;
wire   [4:0] \A[13][189] ;
wire   [4:0] \A[13][190] ;
wire   [4:0] \A[13][191] ;
wire   [4:0] \A[13][192] ;
wire   [4:0] \A[13][193] ;
wire   [4:0] \A[13][194] ;
wire   [4:0] \A[13][195] ;
wire   [4:0] \A[13][196] ;
wire   [4:0] \A[13][197] ;
wire   [4:0] \A[13][198] ;
wire   [4:0] \A[13][199] ;
wire   [4:0] \A[13][200] ;
wire   [4:0] \A[13][201] ;
wire   [4:0] \A[13][202] ;
wire   [4:0] \A[13][203] ;
wire   [4:0] \A[13][204] ;
wire   [4:0] \A[13][205] ;
wire   [4:0] \A[13][206] ;
wire   [4:0] \A[13][207] ;
wire   [4:0] \A[13][208] ;
wire   [4:0] \A[13][209] ;
wire   [4:0] \A[13][210] ;
wire   [4:0] \A[13][211] ;
wire   [4:0] \A[13][212] ;
wire   [4:0] \A[13][213] ;
wire   [4:0] \A[13][214] ;
wire   [4:0] \A[13][215] ;
wire   [4:0] \A[13][216] ;
wire   [4:0] \A[13][217] ;
wire   [4:0] \A[13][218] ;
wire   [4:0] \A[13][219] ;
wire   [4:0] \A[13][220] ;
wire   [4:0] \A[13][221] ;
wire   [4:0] \A[13][222] ;
wire   [4:0] \A[13][223] ;
wire   [4:0] \A[13][224] ;
wire   [4:0] \A[13][225] ;
wire   [4:0] \A[13][226] ;
wire   [4:0] \A[13][227] ;
wire   [4:0] \A[13][228] ;
wire   [4:0] \A[13][229] ;
wire   [4:0] \A[13][230] ;
wire   [4:0] \A[13][231] ;
wire   [4:0] \A[13][232] ;
wire   [4:0] \A[13][233] ;
wire   [4:0] \A[13][234] ;
wire   [4:0] \A[13][235] ;
wire   [4:0] \A[13][236] ;
wire   [4:0] \A[13][237] ;
wire   [4:0] \A[13][238] ;
wire   [4:0] \A[13][239] ;
wire   [4:0] \A[13][240] ;
wire   [4:0] \A[13][241] ;
wire   [4:0] \A[13][242] ;
wire   [4:0] \A[13][243] ;
wire   [4:0] \A[13][244] ;
wire   [4:0] \A[13][245] ;
wire   [4:0] \A[13][246] ;
wire   [4:0] \A[13][247] ;
wire   [4:0] \A[13][248] ;
wire   [4:0] \A[13][249] ;
wire   [4:0] \A[13][250] ;
wire   [4:0] \A[13][251] ;
wire   [4:0] \A[13][252] ;
wire   [4:0] \A[13][253] ;
wire   [4:0] \A[13][254] ;
wire   [4:0] \A[13][255] ;
wire   [4:0] \A[14][0] ;
wire   [4:0] \A[14][1] ;
wire   [4:0] \A[14][2] ;
wire   [4:0] \A[14][3] ;
wire   [4:0] \A[14][4] ;
wire   [4:0] \A[14][5] ;
wire   [4:0] \A[14][6] ;
wire   [4:0] \A[14][7] ;
wire   [4:0] \A[14][8] ;
wire   [4:0] \A[14][9] ;
wire   [4:0] \A[14][10] ;
wire   [4:0] \A[14][11] ;
wire   [4:0] \A[14][12] ;
wire   [4:0] \A[14][13] ;
wire   [4:0] \A[14][14] ;
wire   [4:0] \A[14][15] ;
wire   [4:0] \A[14][16] ;
wire   [4:0] \A[14][17] ;
wire   [4:0] \A[14][18] ;
wire   [4:0] \A[14][19] ;
wire   [4:0] \A[14][20] ;
wire   [4:0] \A[14][21] ;
wire   [4:0] \A[14][22] ;
wire   [4:0] \A[14][23] ;
wire   [4:0] \A[14][24] ;
wire   [4:0] \A[14][25] ;
wire   [4:0] \A[14][26] ;
wire   [4:0] \A[14][27] ;
wire   [4:0] \A[14][28] ;
wire   [4:0] \A[14][29] ;
wire   [4:0] \A[14][30] ;
wire   [4:0] \A[14][31] ;
wire   [4:0] \A[14][32] ;
wire   [4:0] \A[14][33] ;
wire   [4:0] \A[14][34] ;
wire   [4:0] \A[14][35] ;
wire   [4:0] \A[14][36] ;
wire   [4:0] \A[14][37] ;
wire   [4:0] \A[14][38] ;
wire   [4:0] \A[14][39] ;
wire   [4:0] \A[14][40] ;
wire   [4:0] \A[14][41] ;
wire   [4:0] \A[14][42] ;
wire   [4:0] \A[14][43] ;
wire   [4:0] \A[14][44] ;
wire   [4:0] \A[14][45] ;
wire   [4:0] \A[14][46] ;
wire   [4:0] \A[14][47] ;
wire   [4:0] \A[14][48] ;
wire   [4:0] \A[14][49] ;
wire   [4:0] \A[14][50] ;
wire   [4:0] \A[14][51] ;
wire   [4:0] \A[14][52] ;
wire   [4:0] \A[14][53] ;
wire   [4:0] \A[14][54] ;
wire   [4:0] \A[14][55] ;
wire   [4:0] \A[14][56] ;
wire   [4:0] \A[14][57] ;
wire   [4:0] \A[14][58] ;
wire   [4:0] \A[14][59] ;
wire   [4:0] \A[14][60] ;
wire   [4:0] \A[14][61] ;
wire   [4:0] \A[14][62] ;
wire   [4:0] \A[14][63] ;
wire   [4:0] \A[14][64] ;
wire   [4:0] \A[14][65] ;
wire   [4:0] \A[14][66] ;
wire   [4:0] \A[14][67] ;
wire   [4:0] \A[14][68] ;
wire   [4:0] \A[14][69] ;
wire   [4:0] \A[14][70] ;
wire   [4:0] \A[14][71] ;
wire   [4:0] \A[14][72] ;
wire   [4:0] \A[14][73] ;
wire   [4:0] \A[14][74] ;
wire   [4:0] \A[14][75] ;
wire   [4:0] \A[14][76] ;
wire   [4:0] \A[14][77] ;
wire   [4:0] \A[14][78] ;
wire   [4:0] \A[14][79] ;
wire   [4:0] \A[14][80] ;
wire   [4:0] \A[14][81] ;
wire   [4:0] \A[14][82] ;
wire   [4:0] \A[14][83] ;
wire   [4:0] \A[14][84] ;
wire   [4:0] \A[14][85] ;
wire   [4:0] \A[14][86] ;
wire   [4:0] \A[14][87] ;
wire   [4:0] \A[14][88] ;
wire   [4:0] \A[14][89] ;
wire   [4:0] \A[14][90] ;
wire   [4:0] \A[14][91] ;
wire   [4:0] \A[14][92] ;
wire   [4:0] \A[14][93] ;
wire   [4:0] \A[14][94] ;
wire   [4:0] \A[14][95] ;
wire   [4:0] \A[14][96] ;
wire   [4:0] \A[14][97] ;
wire   [4:0] \A[14][98] ;
wire   [4:0] \A[14][99] ;
wire   [4:0] \A[14][100] ;
wire   [4:0] \A[14][101] ;
wire   [4:0] \A[14][102] ;
wire   [4:0] \A[14][103] ;
wire   [4:0] \A[14][104] ;
wire   [4:0] \A[14][105] ;
wire   [4:0] \A[14][106] ;
wire   [4:0] \A[14][107] ;
wire   [4:0] \A[14][108] ;
wire   [4:0] \A[14][109] ;
wire   [4:0] \A[14][110] ;
wire   [4:0] \A[14][111] ;
wire   [4:0] \A[14][112] ;
wire   [4:0] \A[14][113] ;
wire   [4:0] \A[14][114] ;
wire   [4:0] \A[14][115] ;
wire   [4:0] \A[14][116] ;
wire   [4:0] \A[14][117] ;
wire   [4:0] \A[14][118] ;
wire   [4:0] \A[14][119] ;
wire   [4:0] \A[14][120] ;
wire   [4:0] \A[14][121] ;
wire   [4:0] \A[14][122] ;
wire   [4:0] \A[14][123] ;
wire   [4:0] \A[14][124] ;
wire   [4:0] \A[14][125] ;
wire   [4:0] \A[14][126] ;
wire   [4:0] \A[14][127] ;
wire   [4:0] \A[14][128] ;
wire   [4:0] \A[14][129] ;
wire   [4:0] \A[14][130] ;
wire   [4:0] \A[14][131] ;
wire   [4:0] \A[14][132] ;
wire   [4:0] \A[14][133] ;
wire   [4:0] \A[14][134] ;
wire   [4:0] \A[14][135] ;
wire   [4:0] \A[14][136] ;
wire   [4:0] \A[14][137] ;
wire   [4:0] \A[14][138] ;
wire   [4:0] \A[14][139] ;
wire   [4:0] \A[14][140] ;
wire   [4:0] \A[14][141] ;
wire   [4:0] \A[14][142] ;
wire   [4:0] \A[14][143] ;
wire   [4:0] \A[14][144] ;
wire   [4:0] \A[14][145] ;
wire   [4:0] \A[14][146] ;
wire   [4:0] \A[14][147] ;
wire   [4:0] \A[14][148] ;
wire   [4:0] \A[14][149] ;
wire   [4:0] \A[14][150] ;
wire   [4:0] \A[14][151] ;
wire   [4:0] \A[14][152] ;
wire   [4:0] \A[14][153] ;
wire   [4:0] \A[14][154] ;
wire   [4:0] \A[14][155] ;
wire   [4:0] \A[14][156] ;
wire   [4:0] \A[14][157] ;
wire   [4:0] \A[14][158] ;
wire   [4:0] \A[14][159] ;
wire   [4:0] \A[14][160] ;
wire   [4:0] \A[14][161] ;
wire   [4:0] \A[14][162] ;
wire   [4:0] \A[14][163] ;
wire   [4:0] \A[14][164] ;
wire   [4:0] \A[14][165] ;
wire   [4:0] \A[14][166] ;
wire   [4:0] \A[14][167] ;
wire   [4:0] \A[14][168] ;
wire   [4:0] \A[14][169] ;
wire   [4:0] \A[14][170] ;
wire   [4:0] \A[14][171] ;
wire   [4:0] \A[14][172] ;
wire   [4:0] \A[14][173] ;
wire   [4:0] \A[14][174] ;
wire   [4:0] \A[14][175] ;
wire   [4:0] \A[14][176] ;
wire   [4:0] \A[14][177] ;
wire   [4:0] \A[14][178] ;
wire   [4:0] \A[14][179] ;
wire   [4:0] \A[14][180] ;
wire   [4:0] \A[14][181] ;
wire   [4:0] \A[14][182] ;
wire   [4:0] \A[14][183] ;
wire   [4:0] \A[14][184] ;
wire   [4:0] \A[14][185] ;
wire   [4:0] \A[14][186] ;
wire   [4:0] \A[14][187] ;
wire   [4:0] \A[14][188] ;
wire   [4:0] \A[14][189] ;
wire   [4:0] \A[14][190] ;
wire   [4:0] \A[14][191] ;
wire   [4:0] \A[14][192] ;
wire   [4:0] \A[14][193] ;
wire   [4:0] \A[14][194] ;
wire   [4:0] \A[14][195] ;
wire   [4:0] \A[14][196] ;
wire   [4:0] \A[14][197] ;
wire   [4:0] \A[14][198] ;
wire   [4:0] \A[14][199] ;
wire   [4:0] \A[14][200] ;
wire   [4:0] \A[14][201] ;
wire   [4:0] \A[14][202] ;
wire   [4:0] \A[14][203] ;
wire   [4:0] \A[14][204] ;
wire   [4:0] \A[14][205] ;
wire   [4:0] \A[14][206] ;
wire   [4:0] \A[14][207] ;
wire   [4:0] \A[14][208] ;
wire   [4:0] \A[14][209] ;
wire   [4:0] \A[14][210] ;
wire   [4:0] \A[14][211] ;
wire   [4:0] \A[14][212] ;
wire   [4:0] \A[14][213] ;
wire   [4:0] \A[14][214] ;
wire   [4:0] \A[14][215] ;
wire   [4:0] \A[14][216] ;
wire   [4:0] \A[14][217] ;
wire   [4:0] \A[14][218] ;
wire   [4:0] \A[14][219] ;
wire   [4:0] \A[14][220] ;
wire   [4:0] \A[14][221] ;
wire   [4:0] \A[14][222] ;
wire   [4:0] \A[14][223] ;
wire   [4:0] \A[14][224] ;
wire   [4:0] \A[14][225] ;
wire   [4:0] \A[14][226] ;
wire   [4:0] \A[14][227] ;
wire   [4:0] \A[14][228] ;
wire   [4:0] \A[14][229] ;
wire   [4:0] \A[14][230] ;
wire   [4:0] \A[14][231] ;
wire   [4:0] \A[14][232] ;
wire   [4:0] \A[14][233] ;
wire   [4:0] \A[14][234] ;
wire   [4:0] \A[14][235] ;
wire   [4:0] \A[14][236] ;
wire   [4:0] \A[14][237] ;
wire   [4:0] \A[14][238] ;
wire   [4:0] \A[14][239] ;
wire   [4:0] \A[14][240] ;
wire   [4:0] \A[14][241] ;
wire   [4:0] \A[14][242] ;
wire   [4:0] \A[14][243] ;
wire   [4:0] \A[14][244] ;
wire   [4:0] \A[14][245] ;
wire   [4:0] \A[14][246] ;
wire   [4:0] \A[14][247] ;
wire   [4:0] \A[14][248] ;
wire   [4:0] \A[14][249] ;
wire   [4:0] \A[14][250] ;
wire   [4:0] \A[14][251] ;
wire   [4:0] \A[14][252] ;
wire   [4:0] \A[14][253] ;
wire   [4:0] \A[14][254] ;
wire   [4:0] \A[14][255] ;
wire   [4:0] \A[15][0] ;
wire   [4:0] \A[15][1] ;
wire   [4:0] \A[15][2] ;
wire   [4:0] \A[15][3] ;
wire   [4:0] \A[15][4] ;
wire   [4:0] \A[15][5] ;
wire   [4:0] \A[15][6] ;
wire   [4:0] \A[15][7] ;
wire   [4:0] \A[15][8] ;
wire   [4:0] \A[15][9] ;
wire   [4:0] \A[15][10] ;
wire   [4:0] \A[15][11] ;
wire   [4:0] \A[15][12] ;
wire   [4:0] \A[15][13] ;
wire   [4:0] \A[15][14] ;
wire   [4:0] \A[15][15] ;
wire   [4:0] \A[15][16] ;
wire   [4:0] \A[15][17] ;
wire   [4:0] \A[15][18] ;
wire   [4:0] \A[15][19] ;
wire   [4:0] \A[15][20] ;
wire   [4:0] \A[15][21] ;
wire   [4:0] \A[15][22] ;
wire   [4:0] \A[15][23] ;
wire   [4:0] \A[15][24] ;
wire   [4:0] \A[15][25] ;
wire   [4:0] \A[15][26] ;
wire   [4:0] \A[15][27] ;
wire   [4:0] \A[15][28] ;
wire   [4:0] \A[15][29] ;
wire   [4:0] \A[15][30] ;
wire   [4:0] \A[15][31] ;
wire   [4:0] \A[15][32] ;
wire   [4:0] \A[15][33] ;
wire   [4:0] \A[15][34] ;
wire   [4:0] \A[15][35] ;
wire   [4:0] \A[15][36] ;
wire   [4:0] \A[15][37] ;
wire   [4:0] \A[15][38] ;
wire   [4:0] \A[15][39] ;
wire   [4:0] \A[15][40] ;
wire   [4:0] \A[15][41] ;
wire   [4:0] \A[15][42] ;
wire   [4:0] \A[15][43] ;
wire   [4:0] \A[15][44] ;
wire   [4:0] \A[15][45] ;
wire   [4:0] \A[15][46] ;
wire   [4:0] \A[15][47] ;
wire   [4:0] \A[15][48] ;
wire   [4:0] \A[15][49] ;
wire   [4:0] \A[15][50] ;
wire   [4:0] \A[15][51] ;
wire   [4:0] \A[15][52] ;
wire   [4:0] \A[15][53] ;
wire   [4:0] \A[15][54] ;
wire   [4:0] \A[15][55] ;
wire   [4:0] \A[15][56] ;
wire   [4:0] \A[15][57] ;
wire   [4:0] \A[15][58] ;
wire   [4:0] \A[15][59] ;
wire   [4:0] \A[15][60] ;
wire   [4:0] \A[15][61] ;
wire   [4:0] \A[15][62] ;
wire   [4:0] \A[15][63] ;
wire   [4:0] \A[15][64] ;
wire   [4:0] \A[15][65] ;
wire   [4:0] \A[15][66] ;
wire   [4:0] \A[15][67] ;
wire   [4:0] \A[15][68] ;
wire   [4:0] \A[15][69] ;
wire   [4:0] \A[15][70] ;
wire   [4:0] \A[15][71] ;
wire   [4:0] \A[15][72] ;
wire   [4:0] \A[15][73] ;
wire   [4:0] \A[15][74] ;
wire   [4:0] \A[15][75] ;
wire   [4:0] \A[15][76] ;
wire   [4:0] \A[15][77] ;
wire   [4:0] \A[15][78] ;
wire   [4:0] \A[15][79] ;
wire   [4:0] \A[15][80] ;
wire   [4:0] \A[15][81] ;
wire   [4:0] \A[15][82] ;
wire   [4:0] \A[15][83] ;
wire   [4:0] \A[15][84] ;
wire   [4:0] \A[15][85] ;
wire   [4:0] \A[15][86] ;
wire   [4:0] \A[15][87] ;
wire   [4:0] \A[15][88] ;
wire   [4:0] \A[15][89] ;
wire   [4:0] \A[15][90] ;
wire   [4:0] \A[15][91] ;
wire   [4:0] \A[15][92] ;
wire   [4:0] \A[15][93] ;
wire   [4:0] \A[15][94] ;
wire   [4:0] \A[15][95] ;
wire   [4:0] \A[15][96] ;
wire   [4:0] \A[15][97] ;
wire   [4:0] \A[15][98] ;
wire   [4:0] \A[15][99] ;
wire   [4:0] \A[15][100] ;
wire   [4:0] \A[15][101] ;
wire   [4:0] \A[15][102] ;
wire   [4:0] \A[15][103] ;
wire   [4:0] \A[15][104] ;
wire   [4:0] \A[15][105] ;
wire   [4:0] \A[15][106] ;
wire   [4:0] \A[15][107] ;
wire   [4:0] \A[15][108] ;
wire   [4:0] \A[15][109] ;
wire   [4:0] \A[15][110] ;
wire   [4:0] \A[15][111] ;
wire   [4:0] \A[15][112] ;
wire   [4:0] \A[15][113] ;
wire   [4:0] \A[15][114] ;
wire   [4:0] \A[15][115] ;
wire   [4:0] \A[15][116] ;
wire   [4:0] \A[15][117] ;
wire   [4:0] \A[15][118] ;
wire   [4:0] \A[15][119] ;
wire   [4:0] \A[15][120] ;
wire   [4:0] \A[15][121] ;
wire   [4:0] \A[15][122] ;
wire   [4:0] \A[15][123] ;
wire   [4:0] \A[15][124] ;
wire   [4:0] \A[15][125] ;
wire   [4:0] \A[15][126] ;
wire   [4:0] \A[15][127] ;
wire   [4:0] \A[15][128] ;
wire   [4:0] \A[15][129] ;
wire   [4:0] \A[15][130] ;
wire   [4:0] \A[15][131] ;
wire   [4:0] \A[15][132] ;
wire   [4:0] \A[15][133] ;
wire   [4:0] \A[15][134] ;
wire   [4:0] \A[15][135] ;
wire   [4:0] \A[15][136] ;
wire   [4:0] \A[15][137] ;
wire   [4:0] \A[15][138] ;
wire   [4:0] \A[15][139] ;
wire   [4:0] \A[15][140] ;
wire   [4:0] \A[15][141] ;
wire   [4:0] \A[15][142] ;
wire   [4:0] \A[15][143] ;
wire   [4:0] \A[15][144] ;
wire   [4:0] \A[15][145] ;
wire   [4:0] \A[15][146] ;
wire   [4:0] \A[15][147] ;
wire   [4:0] \A[15][148] ;
wire   [4:0] \A[15][149] ;
wire   [4:0] \A[15][150] ;
wire   [4:0] \A[15][151] ;
wire   [4:0] \A[15][152] ;
wire   [4:0] \A[15][153] ;
wire   [4:0] \A[15][154] ;
wire   [4:0] \A[15][155] ;
wire   [4:0] \A[15][156] ;
wire   [4:0] \A[15][157] ;
wire   [4:0] \A[15][158] ;
wire   [4:0] \A[15][159] ;
wire   [4:0] \A[15][160] ;
wire   [4:0] \A[15][161] ;
wire   [4:0] \A[15][162] ;
wire   [4:0] \A[15][163] ;
wire   [4:0] \A[15][164] ;
wire   [4:0] \A[15][165] ;
wire   [4:0] \A[15][166] ;
wire   [4:0] \A[15][167] ;
wire   [4:0] \A[15][168] ;
wire   [4:0] \A[15][169] ;
wire   [4:0] \A[15][170] ;
wire   [4:0] \A[15][171] ;
wire   [4:0] \A[15][172] ;
wire   [4:0] \A[15][173] ;
wire   [4:0] \A[15][174] ;
wire   [4:0] \A[15][175] ;
wire   [4:0] \A[15][176] ;
wire   [4:0] \A[15][177] ;
wire   [4:0] \A[15][178] ;
wire   [4:0] \A[15][179] ;
wire   [4:0] \A[15][180] ;
wire   [4:0] \A[15][181] ;
wire   [4:0] \A[15][182] ;
wire   [4:0] \A[15][183] ;
wire   [4:0] \A[15][184] ;
wire   [4:0] \A[15][185] ;
wire   [4:0] \A[15][186] ;
wire   [4:0] \A[15][187] ;
wire   [4:0] \A[15][188] ;
wire   [4:0] \A[15][189] ;
wire   [4:0] \A[15][190] ;
wire   [4:0] \A[15][191] ;
wire   [4:0] \A[15][192] ;
wire   [4:0] \A[15][193] ;
wire   [4:0] \A[15][194] ;
wire   [4:0] \A[15][195] ;
wire   [4:0] \A[15][196] ;
wire   [4:0] \A[15][197] ;
wire   [4:0] \A[15][198] ;
wire   [4:0] \A[15][199] ;
wire   [4:0] \A[15][200] ;
wire   [4:0] \A[15][201] ;
wire   [4:0] \A[15][202] ;
wire   [4:0] \A[15][203] ;
wire   [4:0] \A[15][204] ;
wire   [4:0] \A[15][205] ;
wire   [4:0] \A[15][206] ;
wire   [4:0] \A[15][207] ;
wire   [4:0] \A[15][208] ;
wire   [4:0] \A[15][209] ;
wire   [4:0] \A[15][210] ;
wire   [4:0] \A[15][211] ;
wire   [4:0] \A[15][212] ;
wire   [4:0] \A[15][213] ;
wire   [4:0] \A[15][214] ;
wire   [4:0] \A[15][215] ;
wire   [4:0] \A[15][216] ;
wire   [4:0] \A[15][217] ;
wire   [4:0] \A[15][218] ;
wire   [4:0] \A[15][219] ;
wire   [4:0] \A[15][220] ;
wire   [4:0] \A[15][221] ;
wire   [4:0] \A[15][222] ;
wire   [4:0] \A[15][223] ;
wire   [4:0] \A[15][224] ;
wire   [4:0] \A[15][225] ;
wire   [4:0] \A[15][226] ;
wire   [4:0] \A[15][227] ;
wire   [4:0] \A[15][228] ;
wire   [4:0] \A[15][229] ;
wire   [4:0] \A[15][230] ;
wire   [4:0] \A[15][231] ;
wire   [4:0] \A[15][232] ;
wire   [4:0] \A[15][233] ;
wire   [4:0] \A[15][234] ;
wire   [4:0] \A[15][235] ;
wire   [4:0] \A[15][236] ;
wire   [4:0] \A[15][237] ;
wire   [4:0] \A[15][238] ;
wire   [4:0] \A[15][239] ;
wire   [4:0] \A[15][240] ;
wire   [4:0] \A[15][241] ;
wire   [4:0] \A[15][242] ;
wire   [4:0] \A[15][243] ;
wire   [4:0] \A[15][244] ;
wire   [4:0] \A[15][245] ;
wire   [4:0] \A[15][246] ;
wire   [4:0] \A[15][247] ;
wire   [4:0] \A[15][248] ;
wire   [4:0] \A[15][249] ;
wire   [4:0] \A[15][250] ;
wire   [4:0] \A[15][251] ;
wire   [4:0] \A[15][252] ;
wire   [4:0] \A[15][253] ;
wire   [4:0] \A[15][254] ;
wire   [4:0] \A[15][255] ;
wire   [4:0] \A[16][0] ;
wire   [4:0] \A[16][1] ;
wire   [4:0] \A[16][2] ;
wire   [4:0] \A[16][3] ;
wire   [4:0] \A[16][4] ;
wire   [4:0] \A[16][5] ;
wire   [4:0] \A[16][6] ;
wire   [4:0] \A[16][7] ;
wire   [4:0] \A[16][8] ;
wire   [4:0] \A[16][9] ;
wire   [4:0] \A[16][10] ;
wire   [4:0] \A[16][11] ;
wire   [4:0] \A[16][12] ;
wire   [4:0] \A[16][13] ;
wire   [4:0] \A[16][14] ;
wire   [4:0] \A[16][15] ;
wire   [4:0] \A[16][16] ;
wire   [4:0] \A[16][17] ;
wire   [4:0] \A[16][18] ;
wire   [4:0] \A[16][19] ;
wire   [4:0] \A[16][20] ;
wire   [4:0] \A[16][21] ;
wire   [4:0] \A[16][22] ;
wire   [4:0] \A[16][23] ;
wire   [4:0] \A[16][24] ;
wire   [4:0] \A[16][25] ;
wire   [4:0] \A[16][26] ;
wire   [4:0] \A[16][27] ;
wire   [4:0] \A[16][28] ;
wire   [4:0] \A[16][29] ;
wire   [4:0] \A[16][30] ;
wire   [4:0] \A[16][31] ;
wire   [4:0] \A[16][32] ;
wire   [4:0] \A[16][33] ;
wire   [4:0] \A[16][34] ;
wire   [4:0] \A[16][35] ;
wire   [4:0] \A[16][36] ;
wire   [4:0] \A[16][37] ;
wire   [4:0] \A[16][38] ;
wire   [4:0] \A[16][39] ;
wire   [4:0] \A[16][40] ;
wire   [4:0] \A[16][41] ;
wire   [4:0] \A[16][42] ;
wire   [4:0] \A[16][43] ;
wire   [4:0] \A[16][44] ;
wire   [4:0] \A[16][45] ;
wire   [4:0] \A[16][46] ;
wire   [4:0] \A[16][47] ;
wire   [4:0] \A[16][48] ;
wire   [4:0] \A[16][49] ;
wire   [4:0] \A[16][50] ;
wire   [4:0] \A[16][51] ;
wire   [4:0] \A[16][52] ;
wire   [4:0] \A[16][53] ;
wire   [4:0] \A[16][54] ;
wire   [4:0] \A[16][55] ;
wire   [4:0] \A[16][56] ;
wire   [4:0] \A[16][57] ;
wire   [4:0] \A[16][58] ;
wire   [4:0] \A[16][59] ;
wire   [4:0] \A[16][60] ;
wire   [4:0] \A[16][61] ;
wire   [4:0] \A[16][62] ;
wire   [4:0] \A[16][63] ;
wire   [4:0] \A[16][64] ;
wire   [4:0] \A[16][65] ;
wire   [4:0] \A[16][66] ;
wire   [4:0] \A[16][67] ;
wire   [4:0] \A[16][68] ;
wire   [4:0] \A[16][69] ;
wire   [4:0] \A[16][70] ;
wire   [4:0] \A[16][71] ;
wire   [4:0] \A[16][72] ;
wire   [4:0] \A[16][73] ;
wire   [4:0] \A[16][74] ;
wire   [4:0] \A[16][75] ;
wire   [4:0] \A[16][76] ;
wire   [4:0] \A[16][77] ;
wire   [4:0] \A[16][78] ;
wire   [4:0] \A[16][79] ;
wire   [4:0] \A[16][80] ;
wire   [4:0] \A[16][81] ;
wire   [4:0] \A[16][82] ;
wire   [4:0] \A[16][83] ;
wire   [4:0] \A[16][84] ;
wire   [4:0] \A[16][85] ;
wire   [4:0] \A[16][86] ;
wire   [4:0] \A[16][87] ;
wire   [4:0] \A[16][88] ;
wire   [4:0] \A[16][89] ;
wire   [4:0] \A[16][90] ;
wire   [4:0] \A[16][91] ;
wire   [4:0] \A[16][92] ;
wire   [4:0] \A[16][93] ;
wire   [4:0] \A[16][94] ;
wire   [4:0] \A[16][95] ;
wire   [4:0] \A[16][96] ;
wire   [4:0] \A[16][97] ;
wire   [4:0] \A[16][98] ;
wire   [4:0] \A[16][99] ;
wire   [4:0] \A[16][100] ;
wire   [4:0] \A[16][101] ;
wire   [4:0] \A[16][102] ;
wire   [4:0] \A[16][103] ;
wire   [4:0] \A[16][104] ;
wire   [4:0] \A[16][105] ;
wire   [4:0] \A[16][106] ;
wire   [4:0] \A[16][107] ;
wire   [4:0] \A[16][108] ;
wire   [4:0] \A[16][109] ;
wire   [4:0] \A[16][110] ;
wire   [4:0] \A[16][111] ;
wire   [4:0] \A[16][112] ;
wire   [4:0] \A[16][113] ;
wire   [4:0] \A[16][114] ;
wire   [4:0] \A[16][115] ;
wire   [4:0] \A[16][116] ;
wire   [4:0] \A[16][117] ;
wire   [4:0] \A[16][118] ;
wire   [4:0] \A[16][119] ;
wire   [4:0] \A[16][120] ;
wire   [4:0] \A[16][121] ;
wire   [4:0] \A[16][122] ;
wire   [4:0] \A[16][123] ;
wire   [4:0] \A[16][124] ;
wire   [4:0] \A[16][125] ;
wire   [4:0] \A[16][126] ;
wire   [4:0] \A[16][127] ;
wire   [4:0] \A[16][128] ;
wire   [4:0] \A[16][129] ;
wire   [4:0] \A[16][130] ;
wire   [4:0] \A[16][131] ;
wire   [4:0] \A[16][132] ;
wire   [4:0] \A[16][133] ;
wire   [4:0] \A[16][134] ;
wire   [4:0] \A[16][135] ;
wire   [4:0] \A[16][136] ;
wire   [4:0] \A[16][137] ;
wire   [4:0] \A[16][138] ;
wire   [4:0] \A[16][139] ;
wire   [4:0] \A[16][140] ;
wire   [4:0] \A[16][141] ;
wire   [4:0] \A[16][142] ;
wire   [4:0] \A[16][143] ;
wire   [4:0] \A[16][144] ;
wire   [4:0] \A[16][145] ;
wire   [4:0] \A[16][146] ;
wire   [4:0] \A[16][147] ;
wire   [4:0] \A[16][148] ;
wire   [4:0] \A[16][149] ;
wire   [4:0] \A[16][150] ;
wire   [4:0] \A[16][151] ;
wire   [4:0] \A[16][152] ;
wire   [4:0] \A[16][153] ;
wire   [4:0] \A[16][154] ;
wire   [4:0] \A[16][155] ;
wire   [4:0] \A[16][156] ;
wire   [4:0] \A[16][157] ;
wire   [4:0] \A[16][158] ;
wire   [4:0] \A[16][159] ;
wire   [4:0] \A[16][160] ;
wire   [4:0] \A[16][161] ;
wire   [4:0] \A[16][162] ;
wire   [4:0] \A[16][163] ;
wire   [4:0] \A[16][164] ;
wire   [4:0] \A[16][165] ;
wire   [4:0] \A[16][166] ;
wire   [4:0] \A[16][167] ;
wire   [4:0] \A[16][168] ;
wire   [4:0] \A[16][169] ;
wire   [4:0] \A[16][170] ;
wire   [4:0] \A[16][171] ;
wire   [4:0] \A[16][172] ;
wire   [4:0] \A[16][173] ;
wire   [4:0] \A[16][174] ;
wire   [4:0] \A[16][175] ;
wire   [4:0] \A[16][176] ;
wire   [4:0] \A[16][177] ;
wire   [4:0] \A[16][178] ;
wire   [4:0] \A[16][179] ;
wire   [4:0] \A[16][180] ;
wire   [4:0] \A[16][181] ;
wire   [4:0] \A[16][182] ;
wire   [4:0] \A[16][183] ;
wire   [4:0] \A[16][184] ;
wire   [4:0] \A[16][185] ;
wire   [4:0] \A[16][186] ;
wire   [4:0] \A[16][187] ;
wire   [4:0] \A[16][188] ;
wire   [4:0] \A[16][189] ;
wire   [4:0] \A[16][190] ;
wire   [4:0] \A[16][191] ;
wire   [4:0] \A[16][192] ;
wire   [4:0] \A[16][193] ;
wire   [4:0] \A[16][194] ;
wire   [4:0] \A[16][195] ;
wire   [4:0] \A[16][196] ;
wire   [4:0] \A[16][197] ;
wire   [4:0] \A[16][198] ;
wire   [4:0] \A[16][199] ;
wire   [4:0] \A[16][200] ;
wire   [4:0] \A[16][201] ;
wire   [4:0] \A[16][202] ;
wire   [4:0] \A[16][203] ;
wire   [4:0] \A[16][204] ;
wire   [4:0] \A[16][205] ;
wire   [4:0] \A[16][206] ;
wire   [4:0] \A[16][207] ;
wire   [4:0] \A[16][208] ;
wire   [4:0] \A[16][209] ;
wire   [4:0] \A[16][210] ;
wire   [4:0] \A[16][211] ;
wire   [4:0] \A[16][212] ;
wire   [4:0] \A[16][213] ;
wire   [4:0] \A[16][214] ;
wire   [4:0] \A[16][215] ;
wire   [4:0] \A[16][216] ;
wire   [4:0] \A[16][217] ;
wire   [4:0] \A[16][218] ;
wire   [4:0] \A[16][219] ;
wire   [4:0] \A[16][220] ;
wire   [4:0] \A[16][221] ;
wire   [4:0] \A[16][222] ;
wire   [4:0] \A[16][223] ;
wire   [4:0] \A[16][224] ;
wire   [4:0] \A[16][225] ;
wire   [4:0] \A[16][226] ;
wire   [4:0] \A[16][227] ;
wire   [4:0] \A[16][228] ;
wire   [4:0] \A[16][229] ;
wire   [4:0] \A[16][230] ;
wire   [4:0] \A[16][231] ;
wire   [4:0] \A[16][232] ;
wire   [4:0] \A[16][233] ;
wire   [4:0] \A[16][234] ;
wire   [4:0] \A[16][235] ;
wire   [4:0] \A[16][236] ;
wire   [4:0] \A[16][237] ;
wire   [4:0] \A[16][238] ;
wire   [4:0] \A[16][239] ;
wire   [4:0] \A[16][240] ;
wire   [4:0] \A[16][241] ;
wire   [4:0] \A[16][242] ;
wire   [4:0] \A[16][243] ;
wire   [4:0] \A[16][244] ;
wire   [4:0] \A[16][245] ;
wire   [4:0] \A[16][246] ;
wire   [4:0] \A[16][247] ;
wire   [4:0] \A[16][248] ;
wire   [4:0] \A[16][249] ;
wire   [4:0] \A[16][250] ;
wire   [4:0] \A[16][251] ;
wire   [4:0] \A[16][252] ;
wire   [4:0] \A[16][253] ;
wire   [4:0] \A[16][254] ;
wire   [4:0] \A[16][255] ;
wire   [4:0] \A[17][0] ;
wire   [4:0] \A[17][1] ;
wire   [4:0] \A[17][2] ;
wire   [4:0] \A[17][3] ;
wire   [4:0] \A[17][4] ;
wire   [4:0] \A[17][5] ;
wire   [4:0] \A[17][6] ;
wire   [4:0] \A[17][7] ;
wire   [4:0] \A[17][8] ;
wire   [4:0] \A[17][9] ;
wire   [4:0] \A[17][10] ;
wire   [4:0] \A[17][11] ;
wire   [4:0] \A[17][12] ;
wire   [4:0] \A[17][13] ;
wire   [4:0] \A[17][14] ;
wire   [4:0] \A[17][15] ;
wire   [4:0] \A[17][16] ;
wire   [4:0] \A[17][17] ;
wire   [4:0] \A[17][18] ;
wire   [4:0] \A[17][19] ;
wire   [4:0] \A[17][20] ;
wire   [4:0] \A[17][21] ;
wire   [4:0] \A[17][22] ;
wire   [4:0] \A[17][23] ;
wire   [4:0] \A[17][24] ;
wire   [4:0] \A[17][25] ;
wire   [4:0] \A[17][26] ;
wire   [4:0] \A[17][27] ;
wire   [4:0] \A[17][28] ;
wire   [4:0] \A[17][29] ;
wire   [4:0] \A[17][30] ;
wire   [4:0] \A[17][31] ;
wire   [4:0] \A[17][32] ;
wire   [4:0] \A[17][33] ;
wire   [4:0] \A[17][34] ;
wire   [4:0] \A[17][35] ;
wire   [4:0] \A[17][36] ;
wire   [4:0] \A[17][37] ;
wire   [4:0] \A[17][38] ;
wire   [4:0] \A[17][39] ;
wire   [4:0] \A[17][40] ;
wire   [4:0] \A[17][41] ;
wire   [4:0] \A[17][42] ;
wire   [4:0] \A[17][43] ;
wire   [4:0] \A[17][44] ;
wire   [4:0] \A[17][45] ;
wire   [4:0] \A[17][46] ;
wire   [4:0] \A[17][47] ;
wire   [4:0] \A[17][48] ;
wire   [4:0] \A[17][49] ;
wire   [4:0] \A[17][50] ;
wire   [4:0] \A[17][51] ;
wire   [4:0] \A[17][52] ;
wire   [4:0] \A[17][53] ;
wire   [4:0] \A[17][54] ;
wire   [4:0] \A[17][55] ;
wire   [4:0] \A[17][56] ;
wire   [4:0] \A[17][57] ;
wire   [4:0] \A[17][58] ;
wire   [4:0] \A[17][59] ;
wire   [4:0] \A[17][60] ;
wire   [4:0] \A[17][61] ;
wire   [4:0] \A[17][62] ;
wire   [4:0] \A[17][63] ;
wire   [4:0] \A[17][64] ;
wire   [4:0] \A[17][65] ;
wire   [4:0] \A[17][66] ;
wire   [4:0] \A[17][67] ;
wire   [4:0] \A[17][68] ;
wire   [4:0] \A[17][69] ;
wire   [4:0] \A[17][70] ;
wire   [4:0] \A[17][71] ;
wire   [4:0] \A[17][72] ;
wire   [4:0] \A[17][73] ;
wire   [4:0] \A[17][74] ;
wire   [4:0] \A[17][75] ;
wire   [4:0] \A[17][76] ;
wire   [4:0] \A[17][77] ;
wire   [4:0] \A[17][78] ;
wire   [4:0] \A[17][79] ;
wire   [4:0] \A[17][80] ;
wire   [4:0] \A[17][81] ;
wire   [4:0] \A[17][82] ;
wire   [4:0] \A[17][83] ;
wire   [4:0] \A[17][84] ;
wire   [4:0] \A[17][85] ;
wire   [4:0] \A[17][86] ;
wire   [4:0] \A[17][87] ;
wire   [4:0] \A[17][88] ;
wire   [4:0] \A[17][89] ;
wire   [4:0] \A[17][90] ;
wire   [4:0] \A[17][91] ;
wire   [4:0] \A[17][92] ;
wire   [4:0] \A[17][93] ;
wire   [4:0] \A[17][94] ;
wire   [4:0] \A[17][95] ;
wire   [4:0] \A[17][96] ;
wire   [4:0] \A[17][97] ;
wire   [4:0] \A[17][98] ;
wire   [4:0] \A[17][99] ;
wire   [4:0] \A[17][100] ;
wire   [4:0] \A[17][101] ;
wire   [4:0] \A[17][102] ;
wire   [4:0] \A[17][103] ;
wire   [4:0] \A[17][104] ;
wire   [4:0] \A[17][105] ;
wire   [4:0] \A[17][106] ;
wire   [4:0] \A[17][107] ;
wire   [4:0] \A[17][108] ;
wire   [4:0] \A[17][109] ;
wire   [4:0] \A[17][110] ;
wire   [4:0] \A[17][111] ;
wire   [4:0] \A[17][112] ;
wire   [4:0] \A[17][113] ;
wire   [4:0] \A[17][114] ;
wire   [4:0] \A[17][115] ;
wire   [4:0] \A[17][116] ;
wire   [4:0] \A[17][117] ;
wire   [4:0] \A[17][118] ;
wire   [4:0] \A[17][119] ;
wire   [4:0] \A[17][120] ;
wire   [4:0] \A[17][121] ;
wire   [4:0] \A[17][122] ;
wire   [4:0] \A[17][123] ;
wire   [4:0] \A[17][124] ;
wire   [4:0] \A[17][125] ;
wire   [4:0] \A[17][126] ;
wire   [4:0] \A[17][127] ;
wire   [4:0] \A[17][128] ;
wire   [4:0] \A[17][129] ;
wire   [4:0] \A[17][130] ;
wire   [4:0] \A[17][131] ;
wire   [4:0] \A[17][132] ;
wire   [4:0] \A[17][133] ;
wire   [4:0] \A[17][134] ;
wire   [4:0] \A[17][135] ;
wire   [4:0] \A[17][136] ;
wire   [4:0] \A[17][137] ;
wire   [4:0] \A[17][138] ;
wire   [4:0] \A[17][139] ;
wire   [4:0] \A[17][140] ;
wire   [4:0] \A[17][141] ;
wire   [4:0] \A[17][142] ;
wire   [4:0] \A[17][143] ;
wire   [4:0] \A[17][144] ;
wire   [4:0] \A[17][145] ;
wire   [4:0] \A[17][146] ;
wire   [4:0] \A[17][147] ;
wire   [4:0] \A[17][148] ;
wire   [4:0] \A[17][149] ;
wire   [4:0] \A[17][150] ;
wire   [4:0] \A[17][151] ;
wire   [4:0] \A[17][152] ;
wire   [4:0] \A[17][153] ;
wire   [4:0] \A[17][154] ;
wire   [4:0] \A[17][155] ;
wire   [4:0] \A[17][156] ;
wire   [4:0] \A[17][157] ;
wire   [4:0] \A[17][158] ;
wire   [4:0] \A[17][159] ;
wire   [4:0] \A[17][160] ;
wire   [4:0] \A[17][161] ;
wire   [4:0] \A[17][162] ;
wire   [4:0] \A[17][163] ;
wire   [4:0] \A[17][164] ;
wire   [4:0] \A[17][165] ;
wire   [4:0] \A[17][166] ;
wire   [4:0] \A[17][167] ;
wire   [4:0] \A[17][168] ;
wire   [4:0] \A[17][169] ;
wire   [4:0] \A[17][170] ;
wire   [4:0] \A[17][171] ;
wire   [4:0] \A[17][172] ;
wire   [4:0] \A[17][173] ;
wire   [4:0] \A[17][174] ;
wire   [4:0] \A[17][175] ;
wire   [4:0] \A[17][176] ;
wire   [4:0] \A[17][177] ;
wire   [4:0] \A[17][178] ;
wire   [4:0] \A[17][179] ;
wire   [4:0] \A[17][180] ;
wire   [4:0] \A[17][181] ;
wire   [4:0] \A[17][182] ;
wire   [4:0] \A[17][183] ;
wire   [4:0] \A[17][184] ;
wire   [4:0] \A[17][185] ;
wire   [4:0] \A[17][186] ;
wire   [4:0] \A[17][187] ;
wire   [4:0] \A[17][188] ;
wire   [4:0] \A[17][189] ;
wire   [4:0] \A[17][190] ;
wire   [4:0] \A[17][191] ;
wire   [4:0] \A[17][192] ;
wire   [4:0] \A[17][193] ;
wire   [4:0] \A[17][194] ;
wire   [4:0] \A[17][195] ;
wire   [4:0] \A[17][196] ;
wire   [4:0] \A[17][197] ;
wire   [4:0] \A[17][198] ;
wire   [4:0] \A[17][199] ;
wire   [4:0] \A[17][200] ;
wire   [4:0] \A[17][201] ;
wire   [4:0] \A[17][202] ;
wire   [4:0] \A[17][203] ;
wire   [4:0] \A[17][204] ;
wire   [4:0] \A[17][205] ;
wire   [4:0] \A[17][206] ;
wire   [4:0] \A[17][207] ;
wire   [4:0] \A[17][208] ;
wire   [4:0] \A[17][209] ;
wire   [4:0] \A[17][210] ;
wire   [4:0] \A[17][211] ;
wire   [4:0] \A[17][212] ;
wire   [4:0] \A[17][213] ;
wire   [4:0] \A[17][214] ;
wire   [4:0] \A[17][215] ;
wire   [4:0] \A[17][216] ;
wire   [4:0] \A[17][217] ;
wire   [4:0] \A[17][218] ;
wire   [4:0] \A[17][219] ;
wire   [4:0] \A[17][220] ;
wire   [4:0] \A[17][221] ;
wire   [4:0] \A[17][222] ;
wire   [4:0] \A[17][223] ;
wire   [4:0] \A[17][224] ;
wire   [4:0] \A[17][225] ;
wire   [4:0] \A[17][226] ;
wire   [4:0] \A[17][227] ;
wire   [4:0] \A[17][228] ;
wire   [4:0] \A[17][229] ;
wire   [4:0] \A[17][230] ;
wire   [4:0] \A[17][231] ;
wire   [4:0] \A[17][232] ;
wire   [4:0] \A[17][233] ;
wire   [4:0] \A[17][234] ;
wire   [4:0] \A[17][235] ;
wire   [4:0] \A[17][236] ;
wire   [4:0] \A[17][237] ;
wire   [4:0] \A[17][238] ;
wire   [4:0] \A[17][239] ;
wire   [4:0] \A[17][240] ;
wire   [4:0] \A[17][241] ;
wire   [4:0] \A[17][242] ;
wire   [4:0] \A[17][243] ;
wire   [4:0] \A[17][244] ;
wire   [4:0] \A[17][245] ;
wire   [4:0] \A[17][246] ;
wire   [4:0] \A[17][247] ;
wire   [4:0] \A[17][248] ;
wire   [4:0] \A[17][249] ;
wire   [4:0] \A[17][250] ;
wire   [4:0] \A[17][251] ;
wire   [4:0] \A[17][252] ;
wire   [4:0] \A[17][253] ;
wire   [4:0] \A[17][254] ;
wire   [4:0] \A[17][255] ;
wire   [4:0] \A[18][0] ;
wire   [4:0] \A[18][1] ;
wire   [4:0] \A[18][2] ;
wire   [4:0] \A[18][3] ;
wire   [4:0] \A[18][4] ;
wire   [4:0] \A[18][5] ;
wire   [4:0] \A[18][6] ;
wire   [4:0] \A[18][7] ;
wire   [4:0] \A[18][8] ;
wire   [4:0] \A[18][9] ;
wire   [4:0] \A[18][10] ;
wire   [4:0] \A[18][11] ;
wire   [4:0] \A[18][12] ;
wire   [4:0] \A[18][13] ;
wire   [4:0] \A[18][14] ;
wire   [4:0] \A[18][15] ;
wire   [4:0] \A[18][16] ;
wire   [4:0] \A[18][17] ;
wire   [4:0] \A[18][18] ;
wire   [4:0] \A[18][19] ;
wire   [4:0] \A[18][20] ;
wire   [4:0] \A[18][21] ;
wire   [4:0] \A[18][22] ;
wire   [4:0] \A[18][23] ;
wire   [4:0] \A[18][24] ;
wire   [4:0] \A[18][25] ;
wire   [4:0] \A[18][26] ;
wire   [4:0] \A[18][27] ;
wire   [4:0] \A[18][28] ;
wire   [4:0] \A[18][29] ;
wire   [4:0] \A[18][30] ;
wire   [4:0] \A[18][31] ;
wire   [4:0] \A[18][32] ;
wire   [4:0] \A[18][33] ;
wire   [4:0] \A[18][34] ;
wire   [4:0] \A[18][35] ;
wire   [4:0] \A[18][36] ;
wire   [4:0] \A[18][37] ;
wire   [4:0] \A[18][38] ;
wire   [4:0] \A[18][39] ;
wire   [4:0] \A[18][40] ;
wire   [4:0] \A[18][41] ;
wire   [4:0] \A[18][42] ;
wire   [4:0] \A[18][43] ;
wire   [4:0] \A[18][44] ;
wire   [4:0] \A[18][45] ;
wire   [4:0] \A[18][46] ;
wire   [4:0] \A[18][47] ;
wire   [4:0] \A[18][48] ;
wire   [4:0] \A[18][49] ;
wire   [4:0] \A[18][50] ;
wire   [4:0] \A[18][51] ;
wire   [4:0] \A[18][52] ;
wire   [4:0] \A[18][53] ;
wire   [4:0] \A[18][54] ;
wire   [4:0] \A[18][55] ;
wire   [4:0] \A[18][56] ;
wire   [4:0] \A[18][57] ;
wire   [4:0] \A[18][58] ;
wire   [4:0] \A[18][59] ;
wire   [4:0] \A[18][60] ;
wire   [4:0] \A[18][61] ;
wire   [4:0] \A[18][62] ;
wire   [4:0] \A[18][63] ;
wire   [4:0] \A[18][64] ;
wire   [4:0] \A[18][65] ;
wire   [4:0] \A[18][66] ;
wire   [4:0] \A[18][67] ;
wire   [4:0] \A[18][68] ;
wire   [4:0] \A[18][69] ;
wire   [4:0] \A[18][70] ;
wire   [4:0] \A[18][71] ;
wire   [4:0] \A[18][72] ;
wire   [4:0] \A[18][73] ;
wire   [4:0] \A[18][74] ;
wire   [4:0] \A[18][75] ;
wire   [4:0] \A[18][76] ;
wire   [4:0] \A[18][77] ;
wire   [4:0] \A[18][78] ;
wire   [4:0] \A[18][79] ;
wire   [4:0] \A[18][80] ;
wire   [4:0] \A[18][81] ;
wire   [4:0] \A[18][82] ;
wire   [4:0] \A[18][83] ;
wire   [4:0] \A[18][84] ;
wire   [4:0] \A[18][85] ;
wire   [4:0] \A[18][86] ;
wire   [4:0] \A[18][87] ;
wire   [4:0] \A[18][88] ;
wire   [4:0] \A[18][89] ;
wire   [4:0] \A[18][90] ;
wire   [4:0] \A[18][91] ;
wire   [4:0] \A[18][92] ;
wire   [4:0] \A[18][93] ;
wire   [4:0] \A[18][94] ;
wire   [4:0] \A[18][95] ;
wire   [4:0] \A[18][96] ;
wire   [4:0] \A[18][97] ;
wire   [4:0] \A[18][98] ;
wire   [4:0] \A[18][99] ;
wire   [4:0] \A[18][100] ;
wire   [4:0] \A[18][101] ;
wire   [4:0] \A[18][102] ;
wire   [4:0] \A[18][103] ;
wire   [4:0] \A[18][104] ;
wire   [4:0] \A[18][105] ;
wire   [4:0] \A[18][106] ;
wire   [4:0] \A[18][107] ;
wire   [4:0] \A[18][108] ;
wire   [4:0] \A[18][109] ;
wire   [4:0] \A[18][110] ;
wire   [4:0] \A[18][111] ;
wire   [4:0] \A[18][112] ;
wire   [4:0] \A[18][113] ;
wire   [4:0] \A[18][114] ;
wire   [4:0] \A[18][115] ;
wire   [4:0] \A[18][116] ;
wire   [4:0] \A[18][117] ;
wire   [4:0] \A[18][118] ;
wire   [4:0] \A[18][119] ;
wire   [4:0] \A[18][120] ;
wire   [4:0] \A[18][121] ;
wire   [4:0] \A[18][122] ;
wire   [4:0] \A[18][123] ;
wire   [4:0] \A[18][124] ;
wire   [4:0] \A[18][125] ;
wire   [4:0] \A[18][126] ;
wire   [4:0] \A[18][127] ;
wire   [4:0] \A[18][128] ;
wire   [4:0] \A[18][129] ;
wire   [4:0] \A[18][130] ;
wire   [4:0] \A[18][131] ;
wire   [4:0] \A[18][132] ;
wire   [4:0] \A[18][133] ;
wire   [4:0] \A[18][134] ;
wire   [4:0] \A[18][135] ;
wire   [4:0] \A[18][136] ;
wire   [4:0] \A[18][137] ;
wire   [4:0] \A[18][138] ;
wire   [4:0] \A[18][139] ;
wire   [4:0] \A[18][140] ;
wire   [4:0] \A[18][141] ;
wire   [4:0] \A[18][142] ;
wire   [4:0] \A[18][143] ;
wire   [4:0] \A[18][144] ;
wire   [4:0] \A[18][145] ;
wire   [4:0] \A[18][146] ;
wire   [4:0] \A[18][147] ;
wire   [4:0] \A[18][148] ;
wire   [4:0] \A[18][149] ;
wire   [4:0] \A[18][150] ;
wire   [4:0] \A[18][151] ;
wire   [4:0] \A[18][152] ;
wire   [4:0] \A[18][153] ;
wire   [4:0] \A[18][154] ;
wire   [4:0] \A[18][155] ;
wire   [4:0] \A[18][156] ;
wire   [4:0] \A[18][157] ;
wire   [4:0] \A[18][158] ;
wire   [4:0] \A[18][159] ;
wire   [4:0] \A[18][160] ;
wire   [4:0] \A[18][161] ;
wire   [4:0] \A[18][162] ;
wire   [4:0] \A[18][163] ;
wire   [4:0] \A[18][164] ;
wire   [4:0] \A[18][165] ;
wire   [4:0] \A[18][166] ;
wire   [4:0] \A[18][167] ;
wire   [4:0] \A[18][168] ;
wire   [4:0] \A[18][169] ;
wire   [4:0] \A[18][170] ;
wire   [4:0] \A[18][171] ;
wire   [4:0] \A[18][172] ;
wire   [4:0] \A[18][173] ;
wire   [4:0] \A[18][174] ;
wire   [4:0] \A[18][175] ;
wire   [4:0] \A[18][176] ;
wire   [4:0] \A[18][177] ;
wire   [4:0] \A[18][178] ;
wire   [4:0] \A[18][179] ;
wire   [4:0] \A[18][180] ;
wire   [4:0] \A[18][181] ;
wire   [4:0] \A[18][182] ;
wire   [4:0] \A[18][183] ;
wire   [4:0] \A[18][184] ;
wire   [4:0] \A[18][185] ;
wire   [4:0] \A[18][186] ;
wire   [4:0] \A[18][187] ;
wire   [4:0] \A[18][188] ;
wire   [4:0] \A[18][189] ;
wire   [4:0] \A[18][190] ;
wire   [4:0] \A[18][191] ;
wire   [4:0] \A[18][192] ;
wire   [4:0] \A[18][193] ;
wire   [4:0] \A[18][194] ;
wire   [4:0] \A[18][195] ;
wire   [4:0] \A[18][196] ;
wire   [4:0] \A[18][197] ;
wire   [4:0] \A[18][198] ;
wire   [4:0] \A[18][199] ;
wire   [4:0] \A[18][200] ;
wire   [4:0] \A[18][201] ;
wire   [4:0] \A[18][202] ;
wire   [4:0] \A[18][203] ;
wire   [4:0] \A[18][204] ;
wire   [4:0] \A[18][205] ;
wire   [4:0] \A[18][206] ;
wire   [4:0] \A[18][207] ;
wire   [4:0] \A[18][208] ;
wire   [4:0] \A[18][209] ;
wire   [4:0] \A[18][210] ;
wire   [4:0] \A[18][211] ;
wire   [4:0] \A[18][212] ;
wire   [4:0] \A[18][213] ;
wire   [4:0] \A[18][214] ;
wire   [4:0] \A[18][215] ;
wire   [4:0] \A[18][216] ;
wire   [4:0] \A[18][217] ;
wire   [4:0] \A[18][218] ;
wire   [4:0] \A[18][219] ;
wire   [4:0] \A[18][220] ;
wire   [4:0] \A[18][221] ;
wire   [4:0] \A[18][222] ;
wire   [4:0] \A[18][223] ;
wire   [4:0] \A[18][224] ;
wire   [4:0] \A[18][225] ;
wire   [4:0] \A[18][226] ;
wire   [4:0] \A[18][227] ;
wire   [4:0] \A[18][228] ;
wire   [4:0] \A[18][229] ;
wire   [4:0] \A[18][230] ;
wire   [4:0] \A[18][231] ;
wire   [4:0] \A[18][232] ;
wire   [4:0] \A[18][233] ;
wire   [4:0] \A[18][234] ;
wire   [4:0] \A[18][235] ;
wire   [4:0] \A[18][236] ;
wire   [4:0] \A[18][237] ;
wire   [4:0] \A[18][238] ;
wire   [4:0] \A[18][239] ;
wire   [4:0] \A[18][240] ;
wire   [4:0] \A[18][241] ;
wire   [4:0] \A[18][242] ;
wire   [4:0] \A[18][243] ;
wire   [4:0] \A[18][244] ;
wire   [4:0] \A[18][245] ;
wire   [4:0] \A[18][246] ;
wire   [4:0] \A[18][247] ;
wire   [4:0] \A[18][248] ;
wire   [4:0] \A[18][249] ;
wire   [4:0] \A[18][250] ;
wire   [4:0] \A[18][251] ;
wire   [4:0] \A[18][252] ;
wire   [4:0] \A[18][253] ;
wire   [4:0] \A[18][254] ;
wire   [4:0] \A[18][255] ;
wire   [4:0] \A[19][0] ;
wire   [4:0] \A[19][1] ;
wire   [4:0] \A[19][2] ;
wire   [4:0] \A[19][3] ;
wire   [4:0] \A[19][4] ;
wire   [4:0] \A[19][5] ;
wire   [4:0] \A[19][6] ;
wire   [4:0] \A[19][7] ;
wire   [4:0] \A[19][8] ;
wire   [4:0] \A[19][9] ;
wire   [4:0] \A[19][10] ;
wire   [4:0] \A[19][11] ;
wire   [4:0] \A[19][12] ;
wire   [4:0] \A[19][13] ;
wire   [4:0] \A[19][14] ;
wire   [4:0] \A[19][15] ;
wire   [4:0] \A[19][16] ;
wire   [4:0] \A[19][17] ;
wire   [4:0] \A[19][18] ;
wire   [4:0] \A[19][19] ;
wire   [4:0] \A[19][20] ;
wire   [4:0] \A[19][21] ;
wire   [4:0] \A[19][22] ;
wire   [4:0] \A[19][23] ;
wire   [4:0] \A[19][24] ;
wire   [4:0] \A[19][25] ;
wire   [4:0] \A[19][26] ;
wire   [4:0] \A[19][27] ;
wire   [4:0] \A[19][28] ;
wire   [4:0] \A[19][29] ;
wire   [4:0] \A[19][30] ;
wire   [4:0] \A[19][31] ;
wire   [4:0] \A[19][32] ;
wire   [4:0] \A[19][33] ;
wire   [4:0] \A[19][34] ;
wire   [4:0] \A[19][35] ;
wire   [4:0] \A[19][36] ;
wire   [4:0] \A[19][37] ;
wire   [4:0] \A[19][38] ;
wire   [4:0] \A[19][39] ;
wire   [4:0] \A[19][40] ;
wire   [4:0] \A[19][41] ;
wire   [4:0] \A[19][42] ;
wire   [4:0] \A[19][43] ;
wire   [4:0] \A[19][44] ;
wire   [4:0] \A[19][45] ;
wire   [4:0] \A[19][46] ;
wire   [4:0] \A[19][47] ;
wire   [4:0] \A[19][48] ;
wire   [4:0] \A[19][49] ;
wire   [4:0] \A[19][50] ;
wire   [4:0] \A[19][51] ;
wire   [4:0] \A[19][52] ;
wire   [4:0] \A[19][53] ;
wire   [4:0] \A[19][54] ;
wire   [4:0] \A[19][55] ;
wire   [4:0] \A[19][56] ;
wire   [4:0] \A[19][57] ;
wire   [4:0] \A[19][58] ;
wire   [4:0] \A[19][59] ;
wire   [4:0] \A[19][60] ;
wire   [4:0] \A[19][61] ;
wire   [4:0] \A[19][62] ;
wire   [4:0] \A[19][63] ;
wire   [4:0] \A[19][64] ;
wire   [4:0] \A[19][65] ;
wire   [4:0] \A[19][66] ;
wire   [4:0] \A[19][67] ;
wire   [4:0] \A[19][68] ;
wire   [4:0] \A[19][69] ;
wire   [4:0] \A[19][70] ;
wire   [4:0] \A[19][71] ;
wire   [4:0] \A[19][72] ;
wire   [4:0] \A[19][73] ;
wire   [4:0] \A[19][74] ;
wire   [4:0] \A[19][75] ;
wire   [4:0] \A[19][76] ;
wire   [4:0] \A[19][77] ;
wire   [4:0] \A[19][78] ;
wire   [4:0] \A[19][79] ;
wire   [4:0] \A[19][80] ;
wire   [4:0] \A[19][81] ;
wire   [4:0] \A[19][82] ;
wire   [4:0] \A[19][83] ;
wire   [4:0] \A[19][84] ;
wire   [4:0] \A[19][85] ;
wire   [4:0] \A[19][86] ;
wire   [4:0] \A[19][87] ;
wire   [4:0] \A[19][88] ;
wire   [4:0] \A[19][89] ;
wire   [4:0] \A[19][90] ;
wire   [4:0] \A[19][91] ;
wire   [4:0] \A[19][92] ;
wire   [4:0] \A[19][93] ;
wire   [4:0] \A[19][94] ;
wire   [4:0] \A[19][95] ;
wire   [4:0] \A[19][96] ;
wire   [4:0] \A[19][97] ;
wire   [4:0] \A[19][98] ;
wire   [4:0] \A[19][99] ;
wire   [4:0] \A[19][100] ;
wire   [4:0] \A[19][101] ;
wire   [4:0] \A[19][102] ;
wire   [4:0] \A[19][103] ;
wire   [4:0] \A[19][104] ;
wire   [4:0] \A[19][105] ;
wire   [4:0] \A[19][106] ;
wire   [4:0] \A[19][107] ;
wire   [4:0] \A[19][108] ;
wire   [4:0] \A[19][109] ;
wire   [4:0] \A[19][110] ;
wire   [4:0] \A[19][111] ;
wire   [4:0] \A[19][112] ;
wire   [4:0] \A[19][113] ;
wire   [4:0] \A[19][114] ;
wire   [4:0] \A[19][115] ;
wire   [4:0] \A[19][116] ;
wire   [4:0] \A[19][117] ;
wire   [4:0] \A[19][118] ;
wire   [4:0] \A[19][119] ;
wire   [4:0] \A[19][120] ;
wire   [4:0] \A[19][121] ;
wire   [4:0] \A[19][122] ;
wire   [4:0] \A[19][123] ;
wire   [4:0] \A[19][124] ;
wire   [4:0] \A[19][125] ;
wire   [4:0] \A[19][126] ;
wire   [4:0] \A[19][127] ;
wire   [4:0] \A[19][128] ;
wire   [4:0] \A[19][129] ;
wire   [4:0] \A[19][130] ;
wire   [4:0] \A[19][131] ;
wire   [4:0] \A[19][132] ;
wire   [4:0] \A[19][133] ;
wire   [4:0] \A[19][134] ;
wire   [4:0] \A[19][135] ;
wire   [4:0] \A[19][136] ;
wire   [4:0] \A[19][137] ;
wire   [4:0] \A[19][138] ;
wire   [4:0] \A[19][139] ;
wire   [4:0] \A[19][140] ;
wire   [4:0] \A[19][141] ;
wire   [4:0] \A[19][142] ;
wire   [4:0] \A[19][143] ;
wire   [4:0] \A[19][144] ;
wire   [4:0] \A[19][145] ;
wire   [4:0] \A[19][146] ;
wire   [4:0] \A[19][147] ;
wire   [4:0] \A[19][148] ;
wire   [4:0] \A[19][149] ;
wire   [4:0] \A[19][150] ;
wire   [4:0] \A[19][151] ;
wire   [4:0] \A[19][152] ;
wire   [4:0] \A[19][153] ;
wire   [4:0] \A[19][154] ;
wire   [4:0] \A[19][155] ;
wire   [4:0] \A[19][156] ;
wire   [4:0] \A[19][157] ;
wire   [4:0] \A[19][158] ;
wire   [4:0] \A[19][159] ;
wire   [4:0] \A[19][160] ;
wire   [4:0] \A[19][161] ;
wire   [4:0] \A[19][162] ;
wire   [4:0] \A[19][163] ;
wire   [4:0] \A[19][164] ;
wire   [4:0] \A[19][165] ;
wire   [4:0] \A[19][166] ;
wire   [4:0] \A[19][167] ;
wire   [4:0] \A[19][168] ;
wire   [4:0] \A[19][169] ;
wire   [4:0] \A[19][170] ;
wire   [4:0] \A[19][171] ;
wire   [4:0] \A[19][172] ;
wire   [4:0] \A[19][173] ;
wire   [4:0] \A[19][174] ;
wire   [4:0] \A[19][175] ;
wire   [4:0] \A[19][176] ;
wire   [4:0] \A[19][177] ;
wire   [4:0] \A[19][178] ;
wire   [4:0] \A[19][179] ;
wire   [4:0] \A[19][180] ;
wire   [4:0] \A[19][181] ;
wire   [4:0] \A[19][182] ;
wire   [4:0] \A[19][183] ;
wire   [4:0] \A[19][184] ;
wire   [4:0] \A[19][185] ;
wire   [4:0] \A[19][186] ;
wire   [4:0] \A[19][187] ;
wire   [4:0] \A[19][188] ;
wire   [4:0] \A[19][189] ;
wire   [4:0] \A[19][190] ;
wire   [4:0] \A[19][191] ;
wire   [4:0] \A[19][192] ;
wire   [4:0] \A[19][193] ;
wire   [4:0] \A[19][194] ;
wire   [4:0] \A[19][195] ;
wire   [4:0] \A[19][196] ;
wire   [4:0] \A[19][197] ;
wire   [4:0] \A[19][198] ;
wire   [4:0] \A[19][199] ;
wire   [4:0] \A[19][200] ;
wire   [4:0] \A[19][201] ;
wire   [4:0] \A[19][202] ;
wire   [4:0] \A[19][203] ;
wire   [4:0] \A[19][204] ;
wire   [4:0] \A[19][205] ;
wire   [4:0] \A[19][206] ;
wire   [4:0] \A[19][207] ;
wire   [4:0] \A[19][208] ;
wire   [4:0] \A[19][209] ;
wire   [4:0] \A[19][210] ;
wire   [4:0] \A[19][211] ;
wire   [4:0] \A[19][212] ;
wire   [4:0] \A[19][213] ;
wire   [4:0] \A[19][214] ;
wire   [4:0] \A[19][215] ;
wire   [4:0] \A[19][216] ;
wire   [4:0] \A[19][217] ;
wire   [4:0] \A[19][218] ;
wire   [4:0] \A[19][219] ;
wire   [4:0] \A[19][220] ;
wire   [4:0] \A[19][221] ;
wire   [4:0] \A[19][222] ;
wire   [4:0] \A[19][223] ;
wire   [4:0] \A[19][224] ;
wire   [4:0] \A[19][225] ;
wire   [4:0] \A[19][226] ;
wire   [4:0] \A[19][227] ;
wire   [4:0] \A[19][228] ;
wire   [4:0] \A[19][229] ;
wire   [4:0] \A[19][230] ;
wire   [4:0] \A[19][231] ;
wire   [4:0] \A[19][232] ;
wire   [4:0] \A[19][233] ;
wire   [4:0] \A[19][234] ;
wire   [4:0] \A[19][235] ;
wire   [4:0] \A[19][236] ;
wire   [4:0] \A[19][237] ;
wire   [4:0] \A[19][238] ;
wire   [4:0] \A[19][239] ;
wire   [4:0] \A[19][240] ;
wire   [4:0] \A[19][241] ;
wire   [4:0] \A[19][242] ;
wire   [4:0] \A[19][243] ;
wire   [4:0] \A[19][244] ;
wire   [4:0] \A[19][245] ;
wire   [4:0] \A[19][246] ;
wire   [4:0] \A[19][247] ;
wire   [4:0] \A[19][248] ;
wire   [4:0] \A[19][249] ;
wire   [4:0] \A[19][250] ;
wire   [4:0] \A[19][251] ;
wire   [4:0] \A[19][252] ;
wire   [4:0] \A[19][253] ;
wire   [4:0] \A[19][254] ;
wire   [4:0] \A[19][255] ;
wire   [0:255] B;
wire   [179:0] out;
wire   [0:127] in;
  assign N$1 = 1'b0;
  assign N$2 = 1'b0;
  assign N$3 = 1'b0;
  assign N$4 = 1'b0;
  assign N$5 = 1'b0;
  assign N$6 = 1'b0;
  assign N$7 = 1'b0;
  assign N$8 = 1'b0;
  assign N$9 = 1'b0;
  assign N$10 = 1'b0;
  assign N$11 = 1'b0;
  assign N$12 = 1'b0;
  assign N$13 = 1'b0;
  assign N$14 = 1'b0;
  assign N$15 = 1'b0;
  assign N$16 = 1'b0;
  assign N$17 = 1'b0;
  assign N$18 = 1'b0;
  assign N$19 = 1'b0;
  assign N$20 = 1'b0;
  assign N$21 = 1'b0;
  assign N$22 = 1'b0;
  assign N$23 = 1'b0;
  assign N$24 = 1'b0;
  assign N$25 = 1'b0;
  assign N$26 = 1'b0;
  assign N$27 = 1'b0;
  assign N$28 = 1'b0;
  assign N$29 = 1'b0;
  assign N$30 = 1'b0;
  assign N$31 = 1'b0;
  assign N$32 = 1'b0;
  assign N$33 = 1'b0;
  assign N$34 = 1'b0;
  assign N$35 = 1'b0;
  assign N$36 = 1'b0;
  assign N$37 = 1'b0;
  assign N$38 = 1'b0;
  assign N$39 = 1'b0;
  assign N$40 = 1'b0;
  assign N$41 = 1'b0;
  assign N$42 = 1'b0;
  assign N$43 = 1'b0;
  assign N$44 = 1'b0;
  assign N$45 = 1'b0;
  assign N$46 = 1'b0;
  assign N$47 = 1'b0;
  assign N$48 = 1'b0;
  assign N$49 = 1'b0;
  assign N$50 = 1'b0;
  assign N$51 = 1'b0;
  assign N$52 = 1'b0;
  assign N$53 = 1'b0;
  assign N$54 = 1'b0;
  assign N$55 = 1'b0;
  assign N$56 = 1'b0;
  assign N$57 = 1'b0;
  assign N$58 = 1'b0;
  assign N$59 = 1'b0;
  assign N$60 = 1'b0;
  assign N$61 = 1'b0;
  assign N$62 = 1'b0;
  assign N$63 = 1'b0;
  assign N$64 = 1'b0;
  assign N$65 = 1'b0;
  assign N$66 = 1'b0;
  assign N$67 = 1'b0;
  assign N$68 = 1'b0;
  assign N$69 = 1'b0;
  assign N$70 = 1'b0;
  assign N$71 = 1'b0;
  assign N$72 = 1'b0;
  assign N$73 = 1'b0;
  assign N$74 = 1'b0;
  assign N$75 = 1'b0;
  assign N$76 = 1'b0;
  assign N$77 = 1'b0;
  assign N$78 = 1'b0;
  assign N$79 = 1'b0;
  assign N$80 = 1'b0;
  assign N$81 = 1'b0;
  assign N$82 = 1'b0;
  assign N$83 = 1'b0;
  assign N$84 = 1'b0;
  assign N$85 = 1'b0;
  assign N$86 = 1'b0;
  assign N$87 = 1'b0;
  assign N$88 = 1'b0;
  assign N$89 = 1'b0;
  assign N$90 = 1'b0;
  assign N$91 = 1'b0;
  assign N$92 = 1'b0;
  assign N$93 = 1'b0;
  assign N$94 = 1'b0;
  assign N$95 = 1'b0;
  assign N$96 = 1'b0;
  assign N$97 = 1'b0;
  assign N$98 = 1'b0;
  assign N$99 = 1'b0;
  assign N$100 = 1'b0;
  assign N$101 = 1'b0;
  assign N$102 = 1'b0;
  assign N$103 = 1'b0;
  assign N$104 = 1'b0;
  assign N$105 = 1'b0;
  assign N$106 = 1'b0;
  assign N$107 = 1'b0;
  assign N$108 = 1'b0;
  assign N$109 = 1'b0;
  assign N$110 = 1'b0;
  assign N$111 = 1'b0;
  assign N$112 = 1'b0;
  assign N$113 = 1'b0;
  assign N$114 = 1'b0;
  assign N$115 = 1'b0;
  assign N$116 = 1'b0;
  assign N$117 = 1'b0;
  assign N$118 = 1'b0;
  assign N$119 = 1'b0;
  assign N$120 = 1'b0;
  assign N$121 = 1'b0;
  assign N$122 = 1'b0;
  assign N$123 = 1'b0;
  assign N$124 = 1'b0;
  assign N$125 = 1'b0;
  assign N$126 = 1'b0;
  assign N$127 = 1'b0;
  assign N$128 = 1'b0;
  assign N$129 = 1'b0;
  assign N$130 = 1'b0;
  assign N$131 = 1'b0;
  assign N$132 = 1'b0;
  assign N$133 = 1'b0;
  assign N$134 = 1'b0;
  assign N$135 = 1'b0;
  assign N$136 = 1'b0;
  assign N$137 = 1'b0;
  assign N$138 = 1'b0;
  assign N$139 = 1'b0;
  assign N$140 = 1'b0;
  assign N$141 = 1'b0;
  assign N$142 = 1'b0;
  assign N$143 = 1'b0;
  assign N$144 = 1'b0;
  assign N$145 = 1'b0;
  assign N$146 = 1'b0;
  assign N$147 = 1'b0;
  assign N$148 = 1'b0;
  assign N$149 = 1'b0;
  assign N$150 = 1'b0;
  assign N$151 = 1'b0;
  assign N$152 = 1'b0;
  assign N$153 = 1'b0;
  assign N$154 = 1'b0;
  assign N$155 = 1'b0;
  assign N$156 = 1'b0;
  assign N$157 = 1'b0;
  assign N$158 = 1'b0;
  assign N$159 = 1'b0;
  assign N$160 = 1'b0;
  assign N$161 = 1'b0;
  assign N$162 = 1'b0;
  assign N$163 = 1'b0;
  assign N$164 = 1'b0;
  assign N$165 = 1'b0;
  assign N$166 = 1'b0;
  assign N$167 = 1'b0;
  assign N$168 = 1'b0;
  assign N$169 = 1'b0;
  assign N$170 = 1'b0;
  assign N$171 = 1'b0;
  assign N$172 = 1'b0;
  assign N$173 = 1'b0;
  assign N$174 = 1'b0;
  assign N$175 = 1'b0;
  assign N$176 = 1'b0;
  assign N$177 = 1'b0;
  assign N$178 = 1'b0;
  assign N$179 = 1'b0;
  assign N$180 = 1'b0;
  assign N$181 = 1'b0;
  assign N$182 = 1'b0;
  assign N$183 = 1'b0;
  assign N$184 = 1'b0;
  assign N$185 = 1'b0;
  assign N$186 = 1'b0;
  assign N$187 = 1'b0;
  assign N$188 = 1'b0;
  assign N$189 = 1'b0;
  assign N$190 = 1'b0;
  assign N$191 = 1'b0;
  assign N$192 = 1'b0;
  assign N$193 = 1'b0;
  assign N$194 = 1'b0;
  assign N$195 = 1'b0;
  assign N$196 = 1'b0;
  assign N$197 = 1'b0;
  assign N$198 = 1'b0;
  assign N$199 = 1'b0;
  assign N$200 = 1'b0;
  assign N$201 = 1'b0;
  assign N$202 = 1'b0;
  assign N$203 = 1'b0;
  assign N$204 = 1'b0;
  assign N$205 = 1'b0;
  assign N$206 = 1'b0;
  assign N$207 = 1'b0;
  assign N$208 = 1'b0;
  assign N$209 = 1'b0;
  assign N$210 = 1'b0;
  assign N$211 = 1'b0;
  assign N$212 = 1'b0;
  assign N$213 = 1'b0;
  assign N$214 = 1'b0;
  assign N$215 = 1'b0;
  assign N$216 = 1'b0;
  assign N$217 = 1'b0;
  assign N$218 = 1'b0;
  assign N$219 = 1'b0;
  assign N$220 = 1'b0;
  assign N$221 = 1'b0;
  assign N$222 = 1'b0;
  assign N$223 = 1'b0;
  assign N$224 = 1'b0;
  assign N$225 = 1'b0;
  assign N$226 = 1'b0;
  assign N$227 = 1'b0;
  assign N$228 = 1'b0;
  assign N$229 = 1'b0;
  assign N$230 = 1'b0;
  assign N$231 = 1'b0;
  assign N$232 = 1'b0;
  assign N$233 = 1'b0;
  assign N$234 = 1'b0;
  assign N$235 = 1'b0;
  assign N$236 = 1'b0;
  assign N$237 = 1'b0;
  assign N$238 = 1'b0;
  assign N$239 = 1'b0;
  assign N$240 = 1'b0;
  assign N$241 = 1'b0;
  assign N$242 = 1'b0;
  assign N$243 = 1'b0;
  assign N$244 = 1'b0;
  assign N$245 = 1'b0;
  assign N$246 = 1'b0;
  assign N$247 = 1'b0;
  assign N$248 = 1'b0;
  assign N$249 = 1'b0;
  assign N$250 = 1'b0;
  assign N$251 = 1'b0;
  assign N$252 = 1'b0;
  assign N$253 = 1'b0;
  assign N$254 = 1'b0;
  assign N$255 = 1'b0;
  assign N$256 = 1'b0;
  assign N$257 = 1'b0;
  assign N$258 = 1'b0;
  assign N$259 = 1'b0;
  assign N$260 = 1'b0;
  assign N$261 = 1'b0;
  assign N$262 = 1'b0;
  assign N$263 = 1'b0;
  assign N$264 = 1'b0;
  assign N$265 = 1'b0;
  assign \biases_l1[0] [3] = 1'b0;
  assign \biases_l1[0] [2] = 1'b0;
  assign \biases_l1[1] [2] = 1'b0;
  assign \biases_l1[1] [1] = 1'b0;
  assign \biases_l1[2] [6] = 1'b0;
  assign \biases_l1[2] [5] = 1'b0;
  assign \biases_l1[2] [3] = 1'b0;
  assign \biases_l1[2] [2] = 1'b0;
  assign \biases_l1[3] [2] = 1'b0;
  assign \biases_l1[3] [1] = 1'b0;
  assign \biases_l1[3] [0] = 1'b0;
  assign \biases_l1[4] [6] = 1'b0;
  assign \biases_l1[4] [5] = 1'b0;
  assign \biases_l1[4] [4] = 1'b0;
  assign \biases_l1[4] [2] = 1'b0;
  assign \biases_l1[5] [6] = 1'b0;
  assign \biases_l1[5] [5] = 1'b0;
  assign \biases_l1[5] [4] = 1'b0;
  assign \biases_l1[5] [3] = 1'b0;
  assign \biases_l1[5] [1] = 1'b0;
  assign \biases_l1[6] [6] = 1'b0;
  assign \biases_l1[6] [5] = 1'b0;
  assign \biases_l1[6] [4] = 1'b0;
  assign \biases_l1[6] [3] = 1'b0;
  assign \biases_l1[6] [2] = 1'b0;
  assign \biases_l1[7] [6] = 1'b0;
  assign \biases_l1[7] [5] = 1'b0;
  assign \biases_l1[7] [4] = 1'b0;
  assign \biases_l1[7] [2] = 1'b0;
  assign \biases_l1[7] [1] = 1'b0;
  assign \biases_l1[8] [6] = 1'b0;
  assign \biases_l1[8] [5] = 1'b0;
  assign \biases_l1[8] [1] = 1'b0;
  assign \biases_l1[9] [6] = 1'b0;
  assign \biases_l1[9] [5] = 1'b0;
  assign \biases_l1[9] [3] = 1'b0;
  assign \biases_l1[9] [0] = 1'b0;
  assign \biases_l1[10] [4] = 1'b0;
  assign \biases_l1[10] [3] = 1'b0;
  assign \biases_l1[11] [6] = 1'b0;
  assign \biases_l1[11] [5] = 1'b0;
  assign \biases_l1[11] [4] = 1'b0;
  assign \biases_l1[11] [3] = 1'b0;
  assign \biases_l1[11] [1] = 1'b0;
  assign \biases_l1[12] [4] = 1'b0;
  assign \biases_l1[12] [1] = 1'b0;
  assign \biases_l1[12] [0] = 1'b0;
  assign \biases_l1[13] [4] = 1'b0;
  assign \biases_l1[13] [3] = 1'b0;
  assign \biases_l1[13] [2] = 1'b0;
  assign \biases_l1[13] [1] = 1'b0;
  assign \biases_l1[13] [0] = 1'b0;
  assign \biases_l1[14] [4] = 1'b0;
  assign \biases_l1[14] [1] = 1'b0;
  assign \biases_l1[15] [5] = 1'b0;
  assign \biases_l1[15] [1] = 1'b0;
  assign \biases_l1[16] [4] = 1'b0;
  assign \biases_l1[16] [0] = 1'b0;
  assign \biases_l1[17] [6] = 1'b0;
  assign \biases_l1[17] [5] = 1'b0;
  assign \biases_l1[17] [3] = 1'b0;
  assign \biases_l1[17] [2] = 1'b0;
  assign \biases_l1[17] [0] = 1'b0;
  assign \biases_l1[18] [2] = 1'b0;
  assign \biases_l1[18] [0] = 1'b0;
  assign \biases_l1[19] [6] = 1'b0;
  assign \biases_l1[19] [4] = 1'b0;
  assign \biases_l1[19] [2] = 1'b0;
  assign \biases_l1[19] [1] = 1'b0;
  assign \A[0][0] [4] = 1'b0;
  assign \A[0][0] [3] = 1'b0;
  assign \A[0][0] [2] = 1'b0;
  assign \A[0][0] [1] = 1'b0;
  assign \A[0][1] [4] = 1'b0;
  assign \A[0][1] [3] = 1'b0;
  assign \A[0][1] [2] = 1'b0;
  assign \A[0][1] [1] = 1'b0;
  assign \A[0][2] [4] = 1'b0;
  assign \A[0][2] [3] = 1'b0;
  assign \A[0][2] [2] = 1'b0;
  assign \A[0][2] [1] = 1'b0;
  assign \A[0][2] [0] = 1'b0;
  assign \A[0][3] [0] = 1'b0;
  assign \A[0][4] [4] = 1'b0;
  assign \A[0][4] [3] = 1'b0;
  assign \A[0][4] [2] = 1'b0;
  assign \A[0][4] [1] = 1'b0;
  assign \A[0][5] [4] = 1'b0;
  assign \A[0][5] [3] = 1'b0;
  assign \A[0][5] [2] = 1'b0;
  assign \A[0][5] [1] = 1'b0;
  assign \A[0][6] [4] = 1'b0;
  assign \A[0][6] [3] = 1'b0;
  assign \A[0][6] [1] = 1'b0;
  assign \A[0][6] [0] = 1'b0;
  assign \A[0][9] [1] = 1'b0;
  assign \A[0][10] [4] = 1'b0;
  assign \A[0][10] [3] = 1'b0;
  assign \A[0][10] [2] = 1'b0;
  assign \A[0][10] [1] = 1'b0;
  assign \A[0][10] [0] = 1'b0;
  assign \A[0][11] [0] = 1'b0;
  assign \A[0][12] [0] = 1'b0;
  assign \A[0][13] [4] = 1'b0;
  assign \A[0][13] [3] = 1'b0;
  assign \A[0][13] [2] = 1'b0;
  assign \A[0][13] [1] = 1'b0;
  assign \A[0][14] [4] = 1'b0;
  assign \A[0][14] [3] = 1'b0;
  assign \A[0][14] [2] = 1'b0;
  assign \A[0][14] [1] = 1'b0;
  assign \A[0][15] [4] = 1'b0;
  assign \A[0][15] [3] = 1'b0;
  assign \A[0][15] [2] = 1'b0;
  assign \A[0][15] [1] = 1'b0;
  assign \A[0][15] [0] = 1'b0;
  assign \A[0][17] [0] = 1'b0;
  assign \A[0][19] [4] = 1'b0;
  assign \A[0][19] [3] = 1'b0;
  assign \A[0][19] [2] = 1'b0;
  assign \A[0][20] [4] = 1'b0;
  assign \A[0][20] [3] = 1'b0;
  assign \A[0][20] [2] = 1'b0;
  assign \A[0][20] [1] = 1'b0;
  assign \A[0][20] [0] = 1'b0;
  assign \A[0][22] [4] = 1'b0;
  assign \A[0][22] [3] = 1'b0;
  assign \A[0][22] [2] = 1'b0;
  assign \A[0][22] [1] = 1'b0;
  assign \A[0][24] [4] = 1'b0;
  assign \A[0][24] [3] = 1'b0;
  assign \A[0][24] [2] = 1'b0;
  assign \A[0][24] [1] = 1'b0;
  assign \A[0][24] [0] = 1'b0;
  assign \A[0][25] [4] = 1'b0;
  assign \A[0][25] [3] = 1'b0;
  assign \A[0][25] [2] = 1'b0;
  assign \A[0][25] [1] = 1'b0;
  assign \A[0][25] [0] = 1'b0;
  assign \A[0][26] [0] = 1'b0;
  assign \A[0][27] [4] = 1'b0;
  assign \A[0][27] [3] = 1'b0;
  assign \A[0][27] [2] = 1'b0;
  assign \A[0][27] [1] = 1'b0;
  assign \A[0][29] [4] = 1'b0;
  assign \A[0][29] [3] = 1'b0;
  assign \A[0][29] [2] = 1'b0;
  assign \A[0][29] [1] = 1'b0;
  assign \A[0][30] [4] = 1'b0;
  assign \A[0][30] [3] = 1'b0;
  assign \A[0][30] [2] = 1'b0;
  assign \A[0][30] [1] = 1'b0;
  assign \A[0][30] [0] = 1'b0;
  assign \A[0][31] [4] = 1'b0;
  assign \A[0][31] [3] = 1'b0;
  assign \A[0][31] [2] = 1'b0;
  assign \A[0][31] [1] = 1'b0;
  assign \A[0][33] [4] = 1'b0;
  assign \A[0][33] [3] = 1'b0;
  assign \A[0][33] [2] = 1'b0;
  assign \A[0][34] [0] = 1'b0;
  assign \A[0][35] [4] = 1'b0;
  assign \A[0][35] [3] = 1'b0;
  assign \A[0][35] [2] = 1'b0;
  assign \A[0][35] [0] = 1'b0;
  assign \A[0][36] [4] = 1'b0;
  assign \A[0][36] [3] = 1'b0;
  assign \A[0][36] [2] = 1'b0;
  assign \A[0][36] [1] = 1'b0;
  assign \A[0][36] [0] = 1'b0;
  assign \A[0][38] [4] = 1'b0;
  assign \A[0][38] [3] = 1'b0;
  assign \A[0][38] [2] = 1'b0;
  assign \A[0][38] [1] = 1'b0;
  assign \A[0][38] [0] = 1'b0;
  assign \A[0][39] [4] = 1'b0;
  assign \A[0][39] [3] = 1'b0;
  assign \A[0][39] [2] = 1'b0;
  assign \A[0][39] [1] = 1'b0;
  assign \A[0][40] [4] = 1'b0;
  assign \A[0][40] [3] = 1'b0;
  assign \A[0][40] [2] = 1'b0;
  assign \A[0][40] [1] = 1'b0;
  assign \A[0][40] [0] = 1'b0;
  assign \A[0][42] [4] = 1'b0;
  assign \A[0][42] [3] = 1'b0;
  assign \A[0][42] [2] = 1'b0;
  assign \A[0][42] [0] = 1'b0;
  assign \A[0][43] [0] = 1'b0;
  assign \A[0][44] [4] = 1'b0;
  assign \A[0][44] [3] = 1'b0;
  assign \A[0][44] [2] = 1'b0;
  assign \A[0][44] [1] = 1'b0;
  assign \A[0][44] [0] = 1'b0;
  assign \A[0][45] [4] = 1'b0;
  assign \A[0][45] [3] = 1'b0;
  assign \A[0][45] [2] = 1'b0;
  assign \A[0][45] [1] = 1'b0;
  assign \A[0][45] [0] = 1'b0;
  assign \A[0][46] [4] = 1'b0;
  assign \A[0][46] [3] = 1'b0;
  assign \A[0][46] [2] = 1'b0;
  assign \A[0][46] [0] = 1'b0;
  assign \A[0][47] [4] = 1'b0;
  assign \A[0][47] [3] = 1'b0;
  assign \A[0][47] [2] = 1'b0;
  assign \A[0][47] [0] = 1'b0;
  assign \A[0][49] [1] = 1'b0;
  assign \A[0][50] [4] = 1'b0;
  assign \A[0][50] [3] = 1'b0;
  assign \A[0][50] [2] = 1'b0;
  assign \A[0][50] [1] = 1'b0;
  assign \A[0][50] [0] = 1'b0;
  assign \A[0][51] [4] = 1'b0;
  assign \A[0][51] [3] = 1'b0;
  assign \A[0][51] [2] = 1'b0;
  assign \A[0][51] [1] = 1'b0;
  assign \A[0][51] [0] = 1'b0;
  assign \A[0][52] [4] = 1'b0;
  assign \A[0][52] [3] = 1'b0;
  assign \A[0][52] [2] = 1'b0;
  assign \A[0][52] [1] = 1'b0;
  assign \A[0][52] [0] = 1'b0;
  assign \A[0][53] [4] = 1'b0;
  assign \A[0][53] [3] = 1'b0;
  assign \A[0][53] [2] = 1'b0;
  assign \A[0][53] [1] = 1'b0;
  assign \A[0][53] [0] = 1'b0;
  assign \A[0][54] [4] = 1'b0;
  assign \A[0][54] [3] = 1'b0;
  assign \A[0][54] [2] = 1'b0;
  assign \A[0][54] [1] = 1'b0;
  assign \A[0][54] [0] = 1'b0;
  assign \A[0][55] [4] = 1'b0;
  assign \A[0][55] [3] = 1'b0;
  assign \A[0][55] [2] = 1'b0;
  assign \A[0][55] [1] = 1'b0;
  assign \A[0][55] [0] = 1'b0;
  assign \A[0][56] [4] = 1'b0;
  assign \A[0][56] [3] = 1'b0;
  assign \A[0][56] [2] = 1'b0;
  assign \A[0][56] [1] = 1'b0;
  assign \A[0][59] [4] = 1'b0;
  assign \A[0][59] [3] = 1'b0;
  assign \A[0][59] [2] = 1'b0;
  assign \A[0][59] [1] = 1'b0;
  assign \A[0][60] [4] = 1'b0;
  assign \A[0][60] [3] = 1'b0;
  assign \A[0][60] [2] = 1'b0;
  assign \A[0][60] [0] = 1'b0;
  assign \A[0][61] [4] = 1'b0;
  assign \A[0][61] [3] = 1'b0;
  assign \A[0][61] [2] = 1'b0;
  assign \A[0][61] [0] = 1'b0;
  assign \A[0][62] [4] = 1'b0;
  assign \A[0][62] [3] = 1'b0;
  assign \A[0][62] [2] = 1'b0;
  assign \A[0][62] [1] = 1'b0;
  assign \A[0][62] [0] = 1'b0;
  assign \A[0][63] [4] = 1'b0;
  assign \A[0][63] [3] = 1'b0;
  assign \A[0][63] [2] = 1'b0;
  assign \A[0][63] [0] = 1'b0;
  assign \A[0][64] [4] = 1'b0;
  assign \A[0][64] [3] = 1'b0;
  assign \A[0][64] [2] = 1'b0;
  assign \A[0][64] [1] = 1'b0;
  assign \A[0][64] [0] = 1'b0;
  assign \A[0][68] [4] = 1'b0;
  assign \A[0][68] [3] = 1'b0;
  assign \A[0][68] [2] = 1'b0;
  assign \A[0][68] [1] = 1'b0;
  assign \A[0][69] [4] = 1'b0;
  assign \A[0][69] [3] = 1'b0;
  assign \A[0][69] [2] = 1'b0;
  assign \A[0][69] [1] = 1'b0;
  assign \A[0][69] [0] = 1'b0;
  assign \A[0][70] [0] = 1'b0;
  assign \A[0][71] [4] = 1'b0;
  assign \A[0][71] [3] = 1'b0;
  assign \A[0][71] [2] = 1'b0;
  assign \A[0][71] [0] = 1'b0;
  assign \A[0][72] [4] = 1'b0;
  assign \A[0][72] [3] = 1'b0;
  assign \A[0][72] [2] = 1'b0;
  assign \A[0][72] [1] = 1'b0;
  assign \A[0][73] [4] = 1'b0;
  assign \A[0][73] [3] = 1'b0;
  assign \A[0][73] [2] = 1'b0;
  assign \A[0][73] [1] = 1'b0;
  assign \A[0][73] [0] = 1'b0;
  assign \A[0][75] [1] = 1'b0;
  assign \A[0][76] [4] = 1'b0;
  assign \A[0][76] [3] = 1'b0;
  assign \A[0][76] [2] = 1'b0;
  assign \A[0][76] [1] = 1'b0;
  assign \A[0][77] [0] = 1'b0;
  assign \A[0][78] [4] = 1'b0;
  assign \A[0][78] [3] = 1'b0;
  assign \A[0][78] [2] = 1'b0;
  assign \A[0][78] [1] = 1'b0;
  assign \A[0][78] [0] = 1'b0;
  assign \A[0][79] [4] = 1'b0;
  assign \A[0][79] [3] = 1'b0;
  assign \A[0][79] [2] = 1'b0;
  assign \A[0][79] [1] = 1'b0;
  assign \A[0][79] [0] = 1'b0;
  assign \A[0][80] [1] = 1'b0;
  assign \A[0][82] [4] = 1'b0;
  assign \A[0][82] [3] = 1'b0;
  assign \A[0][82] [2] = 1'b0;
  assign \A[0][82] [1] = 1'b0;
  assign \A[0][83] [4] = 1'b0;
  assign \A[0][83] [3] = 1'b0;
  assign \A[0][83] [2] = 1'b0;
  assign \A[0][83] [0] = 1'b0;
  assign \A[0][84] [0] = 1'b0;
  assign \A[0][87] [4] = 1'b0;
  assign \A[0][87] [3] = 1'b0;
  assign \A[0][87] [2] = 1'b0;
  assign \A[0][87] [1] = 1'b0;
  assign \A[0][87] [0] = 1'b0;
  assign \A[0][88] [4] = 1'b0;
  assign \A[0][88] [3] = 1'b0;
  assign \A[0][88] [2] = 1'b0;
  assign \A[0][88] [0] = 1'b0;
  assign \A[0][89] [0] = 1'b0;
  assign \A[0][91] [4] = 1'b0;
  assign \A[0][91] [3] = 1'b0;
  assign \A[0][91] [2] = 1'b0;
  assign \A[0][91] [1] = 1'b0;
  assign \A[0][91] [0] = 1'b0;
  assign \A[0][92] [4] = 1'b0;
  assign \A[0][92] [3] = 1'b0;
  assign \A[0][92] [2] = 1'b0;
  assign \A[0][92] [1] = 1'b0;
  assign \A[0][93] [4] = 1'b0;
  assign \A[0][93] [3] = 1'b0;
  assign \A[0][93] [2] = 1'b0;
  assign \A[0][93] [1] = 1'b0;
  assign \A[0][94] [0] = 1'b0;
  assign \A[0][95] [4] = 1'b0;
  assign \A[0][95] [3] = 1'b0;
  assign \A[0][95] [2] = 1'b0;
  assign \A[0][95] [0] = 1'b0;
  assign \A[0][99] [4] = 1'b0;
  assign \A[0][99] [3] = 1'b0;
  assign \A[0][99] [2] = 1'b0;
  assign \A[0][99] [1] = 1'b0;
  assign \A[0][99] [0] = 1'b0;
  assign \A[0][100] [4] = 1'b0;
  assign \A[0][100] [3] = 1'b0;
  assign \A[0][100] [2] = 1'b0;
  assign \A[0][100] [1] = 1'b0;
  assign \A[0][102] [4] = 1'b0;
  assign \A[0][102] [3] = 1'b0;
  assign \A[0][102] [2] = 1'b0;
  assign \A[0][102] [1] = 1'b0;
  assign \A[0][103] [4] = 1'b0;
  assign \A[0][103] [3] = 1'b0;
  assign \A[0][103] [2] = 1'b0;
  assign \A[0][103] [0] = 1'b0;
  assign \A[0][104] [1] = 1'b0;
  assign \A[0][106] [1] = 1'b0;
  assign \A[0][107] [4] = 1'b0;
  assign \A[0][107] [3] = 1'b0;
  assign \A[0][107] [2] = 1'b0;
  assign \A[0][107] [1] = 1'b0;
  assign \A[0][107] [0] = 1'b0;
  assign \A[0][108] [0] = 1'b0;
  assign \A[0][109] [4] = 1'b0;
  assign \A[0][109] [3] = 1'b0;
  assign \A[0][109] [2] = 1'b0;
  assign \A[0][109] [1] = 1'b0;
  assign \A[0][109] [0] = 1'b0;
  assign \A[0][110] [4] = 1'b0;
  assign \A[0][110] [3] = 1'b0;
  assign \A[0][110] [2] = 1'b0;
  assign \A[0][110] [1] = 1'b0;
  assign \A[0][110] [0] = 1'b0;
  assign \A[0][111] [4] = 1'b0;
  assign \A[0][111] [3] = 1'b0;
  assign \A[0][111] [2] = 1'b0;
  assign \A[0][111] [1] = 1'b0;
  assign \A[0][113] [4] = 1'b0;
  assign \A[0][113] [3] = 1'b0;
  assign \A[0][113] [2] = 1'b0;
  assign \A[0][113] [1] = 1'b0;
  assign \A[0][113] [0] = 1'b0;
  assign \A[0][114] [4] = 1'b0;
  assign \A[0][114] [3] = 1'b0;
  assign \A[0][114] [2] = 1'b0;
  assign \A[0][114] [0] = 1'b0;
  assign \A[0][115] [0] = 1'b0;
  assign \A[0][116] [4] = 1'b0;
  assign \A[0][116] [3] = 1'b0;
  assign \A[0][116] [2] = 1'b0;
  assign \A[0][116] [1] = 1'b0;
  assign \A[0][116] [0] = 1'b0;
  assign \A[0][117] [0] = 1'b0;
  assign \A[0][118] [0] = 1'b0;
  assign \A[0][119] [1] = 1'b0;
  assign \A[0][120] [4] = 1'b0;
  assign \A[0][120] [3] = 1'b0;
  assign \A[0][120] [2] = 1'b0;
  assign \A[0][120] [1] = 1'b0;
  assign \A[0][124] [4] = 1'b0;
  assign \A[0][124] [3] = 1'b0;
  assign \A[0][124] [2] = 1'b0;
  assign \A[0][124] [1] = 1'b0;
  assign \A[0][124] [0] = 1'b0;
  assign \A[0][127] [4] = 1'b0;
  assign \A[0][127] [3] = 1'b0;
  assign \A[0][127] [2] = 1'b0;
  assign \A[0][127] [1] = 1'b0;
  assign \A[0][127] [0] = 1'b0;
  assign \A[0][128] [4] = 1'b0;
  assign \A[0][128] [3] = 1'b0;
  assign \A[0][128] [2] = 1'b0;
  assign \A[0][128] [1] = 1'b0;
  assign \A[0][129] [4] = 1'b0;
  assign \A[0][129] [3] = 1'b0;
  assign \A[0][129] [2] = 1'b0;
  assign \A[0][129] [1] = 1'b0;
  assign \A[0][129] [0] = 1'b0;
  assign \A[0][130] [4] = 1'b0;
  assign \A[0][130] [3] = 1'b0;
  assign \A[0][130] [2] = 1'b0;
  assign \A[0][130] [1] = 1'b0;
  assign \A[0][131] [4] = 1'b0;
  assign \A[0][131] [3] = 1'b0;
  assign \A[0][131] [2] = 1'b0;
  assign \A[0][131] [1] = 1'b0;
  assign \A[0][131] [0] = 1'b0;
  assign \A[0][132] [4] = 1'b0;
  assign \A[0][132] [3] = 1'b0;
  assign \A[0][132] [2] = 1'b0;
  assign \A[0][132] [1] = 1'b0;
  assign \A[0][133] [4] = 1'b0;
  assign \A[0][133] [3] = 1'b0;
  assign \A[0][133] [2] = 1'b0;
  assign \A[0][133] [1] = 1'b0;
  assign \A[0][133] [0] = 1'b0;
  assign \A[0][135] [4] = 1'b0;
  assign \A[0][135] [3] = 1'b0;
  assign \A[0][135] [2] = 1'b0;
  assign \A[0][135] [1] = 1'b0;
  assign \A[0][135] [0] = 1'b0;
  assign \A[0][136] [4] = 1'b0;
  assign \A[0][136] [3] = 1'b0;
  assign \A[0][136] [2] = 1'b0;
  assign \A[0][136] [1] = 1'b0;
  assign \A[0][137] [1] = 1'b0;
  assign \A[0][137] [0] = 1'b0;
  assign \A[0][138] [4] = 1'b0;
  assign \A[0][138] [3] = 1'b0;
  assign \A[0][138] [2] = 1'b0;
  assign \A[0][138] [0] = 1'b0;
  assign \A[0][139] [4] = 1'b0;
  assign \A[0][139] [3] = 1'b0;
  assign \A[0][139] [2] = 1'b0;
  assign \A[0][139] [1] = 1'b0;
  assign \A[0][140] [4] = 1'b0;
  assign \A[0][140] [3] = 1'b0;
  assign \A[0][140] [2] = 1'b0;
  assign \A[0][140] [1] = 1'b0;
  assign \A[0][140] [0] = 1'b0;
  assign \A[0][143] [4] = 1'b0;
  assign \A[0][143] [3] = 1'b0;
  assign \A[0][143] [2] = 1'b0;
  assign \A[0][143] [1] = 1'b0;
  assign \A[0][143] [0] = 1'b0;
  assign \A[0][144] [4] = 1'b0;
  assign \A[0][144] [3] = 1'b0;
  assign \A[0][144] [2] = 1'b0;
  assign \A[0][144] [1] = 1'b0;
  assign \A[0][145] [0] = 1'b0;
  assign \A[0][146] [4] = 1'b0;
  assign \A[0][146] [3] = 1'b0;
  assign \A[0][146] [2] = 1'b0;
  assign \A[0][147] [4] = 1'b0;
  assign \A[0][147] [3] = 1'b0;
  assign \A[0][147] [2] = 1'b0;
  assign \A[0][147] [1] = 1'b0;
  assign \A[0][147] [0] = 1'b0;
  assign \A[0][148] [4] = 1'b0;
  assign \A[0][148] [3] = 1'b0;
  assign \A[0][148] [2] = 1'b0;
  assign \A[0][148] [1] = 1'b0;
  assign \A[0][148] [0] = 1'b0;
  assign \A[0][149] [0] = 1'b0;
  assign \A[0][150] [4] = 1'b0;
  assign \A[0][150] [3] = 1'b0;
  assign \A[0][150] [2] = 1'b0;
  assign \A[0][150] [1] = 1'b0;
  assign \A[0][151] [0] = 1'b0;
  assign \A[0][152] [4] = 1'b0;
  assign \A[0][152] [3] = 1'b0;
  assign \A[0][152] [2] = 1'b0;
  assign \A[0][152] [1] = 1'b0;
  assign \A[0][152] [0] = 1'b0;
  assign \A[0][153] [4] = 1'b0;
  assign \A[0][153] [3] = 1'b0;
  assign \A[0][153] [2] = 1'b0;
  assign \A[0][153] [1] = 1'b0;
  assign \A[0][154] [1] = 1'b0;
  assign \A[0][159] [4] = 1'b0;
  assign \A[0][159] [3] = 1'b0;
  assign \A[0][159] [2] = 1'b0;
  assign \A[0][159] [0] = 1'b0;
  assign \A[0][160] [4] = 1'b0;
  assign \A[0][160] [3] = 1'b0;
  assign \A[0][160] [2] = 1'b0;
  assign \A[0][160] [1] = 1'b0;
  assign \A[0][160] [0] = 1'b0;
  assign \A[0][161] [4] = 1'b0;
  assign \A[0][161] [3] = 1'b0;
  assign \A[0][161] [2] = 1'b0;
  assign \A[0][161] [1] = 1'b0;
  assign \A[0][161] [0] = 1'b0;
  assign \A[0][162] [0] = 1'b0;
  assign \A[0][163] [4] = 1'b0;
  assign \A[0][163] [3] = 1'b0;
  assign \A[0][163] [2] = 1'b0;
  assign \A[0][163] [1] = 1'b0;
  assign \A[0][163] [0] = 1'b0;
  assign \A[0][164] [0] = 1'b0;
  assign \A[0][166] [4] = 1'b0;
  assign \A[0][166] [3] = 1'b0;
  assign \A[0][166] [2] = 1'b0;
  assign \A[0][166] [1] = 1'b0;
  assign \A[0][167] [1] = 1'b0;
  assign \A[0][168] [4] = 1'b0;
  assign \A[0][168] [3] = 1'b0;
  assign \A[0][168] [2] = 1'b0;
  assign \A[0][168] [1] = 1'b0;
  assign \A[0][168] [0] = 1'b0;
  assign \A[0][171] [4] = 1'b0;
  assign \A[0][171] [3] = 1'b0;
  assign \A[0][171] [2] = 1'b0;
  assign \A[0][171] [1] = 1'b0;
  assign \A[0][173] [4] = 1'b0;
  assign \A[0][173] [3] = 1'b0;
  assign \A[0][173] [2] = 1'b0;
  assign \A[0][173] [1] = 1'b0;
  assign \A[0][173] [0] = 1'b0;
  assign \A[0][174] [4] = 1'b0;
  assign \A[0][174] [3] = 1'b0;
  assign \A[0][174] [2] = 1'b0;
  assign \A[0][174] [1] = 1'b0;
  assign \A[0][177] [1] = 1'b0;
  assign \A[0][178] [4] = 1'b0;
  assign \A[0][178] [3] = 1'b0;
  assign \A[0][178] [2] = 1'b0;
  assign \A[0][178] [1] = 1'b0;
  assign \A[0][178] [0] = 1'b0;
  assign \A[0][179] [4] = 1'b0;
  assign \A[0][179] [3] = 1'b0;
  assign \A[0][179] [2] = 1'b0;
  assign \A[0][179] [1] = 1'b0;
  assign \A[0][180] [4] = 1'b0;
  assign \A[0][180] [3] = 1'b0;
  assign \A[0][180] [2] = 1'b0;
  assign \A[0][180] [1] = 1'b0;
  assign \A[0][180] [0] = 1'b0;
  assign \A[0][181] [4] = 1'b0;
  assign \A[0][181] [3] = 1'b0;
  assign \A[0][181] [2] = 1'b0;
  assign \A[0][181] [1] = 1'b0;
  assign \A[0][181] [0] = 1'b0;
  assign \A[0][182] [4] = 1'b0;
  assign \A[0][182] [3] = 1'b0;
  assign \A[0][182] [2] = 1'b0;
  assign \A[0][182] [1] = 1'b0;
  assign \A[0][182] [0] = 1'b0;
  assign \A[0][183] [4] = 1'b0;
  assign \A[0][183] [3] = 1'b0;
  assign \A[0][183] [2] = 1'b0;
  assign \A[0][183] [1] = 1'b0;
  assign \A[0][185] [0] = 1'b0;
  assign \A[0][186] [0] = 1'b0;
  assign \A[0][187] [4] = 1'b0;
  assign \A[0][187] [3] = 1'b0;
  assign \A[0][187] [2] = 1'b0;
  assign \A[0][187] [1] = 1'b0;
  assign \A[0][188] [4] = 1'b0;
  assign \A[0][188] [3] = 1'b0;
  assign \A[0][188] [2] = 1'b0;
  assign \A[0][188] [1] = 1'b0;
  assign \A[0][188] [0] = 1'b0;
  assign \A[0][189] [4] = 1'b0;
  assign \A[0][189] [3] = 1'b0;
  assign \A[0][189] [2] = 1'b0;
  assign \A[0][189] [1] = 1'b0;
  assign \A[0][191] [4] = 1'b0;
  assign \A[0][191] [3] = 1'b0;
  assign \A[0][191] [2] = 1'b0;
  assign \A[0][191] [0] = 1'b0;
  assign \A[0][192] [4] = 1'b0;
  assign \A[0][192] [3] = 1'b0;
  assign \A[0][192] [2] = 1'b0;
  assign \A[0][192] [1] = 1'b0;
  assign \A[0][192] [0] = 1'b0;
  assign \A[0][193] [0] = 1'b0;
  assign \A[0][194] [0] = 1'b0;
  assign \A[0][196] [4] = 1'b0;
  assign \A[0][196] [3] = 1'b0;
  assign \A[0][196] [2] = 1'b0;
  assign \A[0][196] [1] = 1'b0;
  assign \A[0][197] [1] = 1'b0;
  assign \A[0][197] [0] = 1'b0;
  assign \A[0][198] [4] = 1'b0;
  assign \A[0][198] [3] = 1'b0;
  assign \A[0][198] [2] = 1'b0;
  assign \A[0][198] [1] = 1'b0;
  assign \A[0][198] [0] = 1'b0;
  assign \A[0][200] [4] = 1'b0;
  assign \A[0][200] [3] = 1'b0;
  assign \A[0][200] [2] = 1'b0;
  assign \A[0][200] [0] = 1'b0;
  assign \A[0][201] [4] = 1'b0;
  assign \A[0][201] [3] = 1'b0;
  assign \A[0][201] [2] = 1'b0;
  assign \A[0][201] [1] = 1'b0;
  assign \A[0][202] [4] = 1'b0;
  assign \A[0][202] [3] = 1'b0;
  assign \A[0][202] [2] = 1'b0;
  assign \A[0][202] [1] = 1'b0;
  assign \A[0][203] [4] = 1'b0;
  assign \A[0][203] [3] = 1'b0;
  assign \A[0][203] [2] = 1'b0;
  assign \A[0][203] [1] = 1'b0;
  assign \A[0][204] [4] = 1'b0;
  assign \A[0][204] [3] = 1'b0;
  assign \A[0][204] [2] = 1'b0;
  assign \A[0][204] [1] = 1'b0;
  assign \A[0][205] [0] = 1'b0;
  assign \A[0][206] [4] = 1'b0;
  assign \A[0][206] [3] = 1'b0;
  assign \A[0][206] [2] = 1'b0;
  assign \A[0][206] [1] = 1'b0;
  assign \A[0][206] [0] = 1'b0;
  assign \A[0][207] [4] = 1'b0;
  assign \A[0][207] [3] = 1'b0;
  assign \A[0][207] [2] = 1'b0;
  assign \A[0][207] [1] = 1'b0;
  assign \A[0][207] [0] = 1'b0;
  assign \A[0][209] [0] = 1'b0;
  assign \A[0][212] [4] = 1'b0;
  assign \A[0][212] [3] = 1'b0;
  assign \A[0][212] [2] = 1'b0;
  assign \A[0][212] [1] = 1'b0;
  assign \A[0][213] [0] = 1'b0;
  assign \A[0][214] [4] = 1'b0;
  assign \A[0][214] [3] = 1'b0;
  assign \A[0][214] [2] = 1'b0;
  assign \A[0][214] [1] = 1'b0;
  assign \A[0][214] [0] = 1'b0;
  assign \A[0][215] [4] = 1'b0;
  assign \A[0][215] [3] = 1'b0;
  assign \A[0][215] [2] = 1'b0;
  assign \A[0][215] [1] = 1'b0;
  assign \A[0][215] [0] = 1'b0;
  assign \A[0][216] [4] = 1'b0;
  assign \A[0][216] [3] = 1'b0;
  assign \A[0][216] [2] = 1'b0;
  assign \A[0][217] [4] = 1'b0;
  assign \A[0][217] [3] = 1'b0;
  assign \A[0][217] [2] = 1'b0;
  assign \A[0][217] [1] = 1'b0;
  assign \A[0][217] [0] = 1'b0;
  assign \A[0][218] [4] = 1'b0;
  assign \A[0][218] [3] = 1'b0;
  assign \A[0][218] [2] = 1'b0;
  assign \A[0][218] [1] = 1'b0;
  assign \A[0][218] [0] = 1'b0;
  assign \A[0][219] [4] = 1'b0;
  assign \A[0][219] [3] = 1'b0;
  assign \A[0][219] [2] = 1'b0;
  assign \A[0][219] [1] = 1'b0;
  assign \A[0][221] [4] = 1'b0;
  assign \A[0][221] [3] = 1'b0;
  assign \A[0][221] [2] = 1'b0;
  assign \A[0][221] [1] = 1'b0;
  assign \A[0][221] [0] = 1'b0;
  assign \A[0][222] [4] = 1'b0;
  assign \A[0][222] [3] = 1'b0;
  assign \A[0][222] [2] = 1'b0;
  assign \A[0][222] [1] = 1'b0;
  assign \A[0][223] [4] = 1'b0;
  assign \A[0][223] [3] = 1'b0;
  assign \A[0][223] [2] = 1'b0;
  assign \A[0][223] [1] = 1'b0;
  assign \A[0][223] [0] = 1'b0;
  assign \A[0][224] [4] = 1'b0;
  assign \A[0][224] [3] = 1'b0;
  assign \A[0][224] [2] = 1'b0;
  assign \A[0][225] [4] = 1'b0;
  assign \A[0][225] [3] = 1'b0;
  assign \A[0][225] [2] = 1'b0;
  assign \A[0][225] [1] = 1'b0;
  assign \A[0][225] [0] = 1'b0;
  assign \A[0][227] [4] = 1'b0;
  assign \A[0][227] [3] = 1'b0;
  assign \A[0][227] [2] = 1'b0;
  assign \A[0][227] [1] = 1'b0;
  assign \A[0][228] [4] = 1'b0;
  assign \A[0][228] [3] = 1'b0;
  assign \A[0][228] [2] = 1'b0;
  assign \A[0][228] [1] = 1'b0;
  assign \A[0][229] [4] = 1'b0;
  assign \A[0][229] [3] = 1'b0;
  assign \A[0][229] [2] = 1'b0;
  assign \A[0][229] [1] = 1'b0;
  assign \A[0][229] [0] = 1'b0;
  assign \A[0][230] [1] = 1'b0;
  assign \A[0][231] [4] = 1'b0;
  assign \A[0][231] [3] = 1'b0;
  assign \A[0][231] [2] = 1'b0;
  assign \A[0][231] [1] = 1'b0;
  assign \A[0][231] [0] = 1'b0;
  assign \A[0][232] [0] = 1'b0;
  assign \A[0][233] [4] = 1'b0;
  assign \A[0][233] [3] = 1'b0;
  assign \A[0][233] [2] = 1'b0;
  assign \A[0][233] [1] = 1'b0;
  assign \A[0][234] [0] = 1'b0;
  assign \A[0][235] [4] = 1'b0;
  assign \A[0][235] [3] = 1'b0;
  assign \A[0][235] [2] = 1'b0;
  assign \A[0][235] [1] = 1'b0;
  assign \A[0][236] [4] = 1'b0;
  assign \A[0][236] [3] = 1'b0;
  assign \A[0][236] [2] = 1'b0;
  assign \A[0][236] [1] = 1'b0;
  assign \A[0][236] [0] = 1'b0;
  assign \A[0][237] [4] = 1'b0;
  assign \A[0][237] [3] = 1'b0;
  assign \A[0][237] [2] = 1'b0;
  assign \A[0][237] [0] = 1'b0;
  assign \A[0][238] [4] = 1'b0;
  assign \A[0][238] [3] = 1'b0;
  assign \A[0][238] [2] = 1'b0;
  assign \A[0][238] [1] = 1'b0;
  assign \A[0][239] [4] = 1'b0;
  assign \A[0][239] [3] = 1'b0;
  assign \A[0][239] [2] = 1'b0;
  assign \A[0][239] [0] = 1'b0;
  assign \A[0][240] [4] = 1'b0;
  assign \A[0][240] [3] = 1'b0;
  assign \A[0][240] [2] = 1'b0;
  assign \A[0][240] [1] = 1'b0;
  assign \A[0][240] [0] = 1'b0;
  assign \A[0][244] [4] = 1'b0;
  assign \A[0][244] [3] = 1'b0;
  assign \A[0][244] [2] = 1'b0;
  assign \A[0][244] [0] = 1'b0;
  assign \A[0][245] [4] = 1'b0;
  assign \A[0][245] [3] = 1'b0;
  assign \A[0][245] [2] = 1'b0;
  assign \A[0][245] [1] = 1'b0;
  assign \A[0][246] [4] = 1'b0;
  assign \A[0][246] [3] = 1'b0;
  assign \A[0][246] [2] = 1'b0;
  assign \A[0][246] [0] = 1'b0;
  assign \A[0][247] [4] = 1'b0;
  assign \A[0][247] [3] = 1'b0;
  assign \A[0][247] [2] = 1'b0;
  assign \A[0][247] [1] = 1'b0;
  assign \A[0][248] [4] = 1'b0;
  assign \A[0][248] [3] = 1'b0;
  assign \A[0][248] [2] = 1'b0;
  assign \A[0][249] [4] = 1'b0;
  assign \A[0][249] [3] = 1'b0;
  assign \A[0][249] [2] = 1'b0;
  assign \A[0][249] [1] = 1'b0;
  assign \A[0][249] [0] = 1'b0;
  assign \A[0][251] [4] = 1'b0;
  assign \A[0][251] [3] = 1'b0;
  assign \A[0][251] [2] = 1'b0;
  assign \A[0][251] [1] = 1'b0;
  assign \A[0][251] [0] = 1'b0;
  assign \A[0][252] [0] = 1'b0;
  assign \A[0][253] [4] = 1'b0;
  assign \A[0][253] [3] = 1'b0;
  assign \A[0][253] [2] = 1'b0;
  assign \A[0][253] [1] = 1'b0;
  assign \A[0][254] [0] = 1'b0;
  assign \A[1][0] [4] = 1'b0;
  assign \A[1][0] [3] = 1'b0;
  assign \A[1][0] [2] = 1'b0;
  assign \A[1][0] [0] = 1'b0;
  assign \A[1][1] [0] = 1'b0;
  assign \A[1][3] [4] = 1'b0;
  assign \A[1][3] [3] = 1'b0;
  assign \A[1][3] [2] = 1'b0;
  assign \A[1][3] [1] = 1'b0;
  assign \A[1][3] [0] = 1'b0;
  assign \A[1][4] [4] = 1'b0;
  assign \A[1][4] [3] = 1'b0;
  assign \A[1][4] [2] = 1'b0;
  assign \A[1][4] [1] = 1'b0;
  assign \A[1][4] [0] = 1'b0;
  assign \A[1][5] [0] = 1'b0;
  assign \A[1][6] [4] = 1'b0;
  assign \A[1][6] [3] = 1'b0;
  assign \A[1][6] [2] = 1'b0;
  assign \A[1][6] [1] = 1'b0;
  assign \A[1][9] [4] = 1'b0;
  assign \A[1][9] [3] = 1'b0;
  assign \A[1][9] [2] = 1'b0;
  assign \A[1][9] [1] = 1'b0;
  assign \A[1][9] [0] = 1'b0;
  assign \A[1][10] [0] = 1'b0;
  assign \A[1][11] [4] = 1'b0;
  assign \A[1][11] [3] = 1'b0;
  assign \A[1][11] [2] = 1'b0;
  assign \A[1][11] [0] = 1'b0;
  assign \A[1][12] [4] = 1'b0;
  assign \A[1][12] [3] = 1'b0;
  assign \A[1][12] [2] = 1'b0;
  assign \A[1][12] [1] = 1'b0;
  assign \A[1][13] [1] = 1'b0;
  assign \A[1][14] [4] = 1'b0;
  assign \A[1][14] [3] = 1'b0;
  assign \A[1][14] [2] = 1'b0;
  assign \A[1][14] [1] = 1'b0;
  assign \A[1][15] [4] = 1'b0;
  assign \A[1][15] [3] = 1'b0;
  assign \A[1][15] [2] = 1'b0;
  assign \A[1][15] [1] = 1'b0;
  assign \A[1][15] [0] = 1'b0;
  assign \A[1][18] [4] = 1'b0;
  assign \A[1][18] [3] = 1'b0;
  assign \A[1][18] [2] = 1'b0;
  assign \A[1][18] [1] = 1'b0;
  assign \A[1][18] [0] = 1'b0;
  assign \A[1][19] [4] = 1'b0;
  assign \A[1][19] [3] = 1'b0;
  assign \A[1][19] [2] = 1'b0;
  assign \A[1][19] [0] = 1'b0;
  assign \A[1][20] [4] = 1'b0;
  assign \A[1][20] [3] = 1'b0;
  assign \A[1][20] [2] = 1'b0;
  assign \A[1][20] [1] = 1'b0;
  assign \A[1][20] [0] = 1'b0;
  assign \A[1][22] [4] = 1'b0;
  assign \A[1][22] [3] = 1'b0;
  assign \A[1][22] [2] = 1'b0;
  assign \A[1][22] [1] = 1'b0;
  assign \A[1][22] [0] = 1'b0;
  assign \A[1][23] [4] = 1'b0;
  assign \A[1][23] [3] = 1'b0;
  assign \A[1][23] [2] = 1'b0;
  assign \A[1][23] [0] = 1'b0;
  assign \A[1][25] [4] = 1'b0;
  assign \A[1][25] [3] = 1'b0;
  assign \A[1][25] [2] = 1'b0;
  assign \A[1][25] [1] = 1'b0;
  assign \A[1][25] [0] = 1'b0;
  assign \A[1][26] [1] = 1'b0;
  assign \A[1][27] [4] = 1'b0;
  assign \A[1][27] [3] = 1'b0;
  assign \A[1][27] [2] = 1'b0;
  assign \A[1][27] [1] = 1'b0;
  assign \A[1][27] [0] = 1'b0;
  assign \A[1][30] [4] = 1'b0;
  assign \A[1][30] [3] = 1'b0;
  assign \A[1][30] [2] = 1'b0;
  assign \A[1][30] [0] = 1'b0;
  assign \A[1][31] [4] = 1'b0;
  assign \A[1][31] [3] = 1'b0;
  assign \A[1][31] [2] = 1'b0;
  assign \A[1][31] [1] = 1'b0;
  assign \A[1][31] [0] = 1'b0;
  assign \A[1][32] [0] = 1'b0;
  assign \A[1][33] [1] = 1'b0;
  assign \A[1][34] [4] = 1'b0;
  assign \A[1][34] [3] = 1'b0;
  assign \A[1][34] [2] = 1'b0;
  assign \A[1][34] [1] = 1'b0;
  assign \A[1][34] [0] = 1'b0;
  assign \A[1][35] [4] = 1'b0;
  assign \A[1][35] [3] = 1'b0;
  assign \A[1][35] [2] = 1'b0;
  assign \A[1][35] [1] = 1'b0;
  assign \A[1][35] [0] = 1'b0;
  assign \A[1][36] [4] = 1'b0;
  assign \A[1][36] [3] = 1'b0;
  assign \A[1][36] [2] = 1'b0;
  assign \A[1][36] [1] = 1'b0;
  assign \A[1][36] [0] = 1'b0;
  assign \A[1][37] [4] = 1'b0;
  assign \A[1][37] [3] = 1'b0;
  assign \A[1][37] [2] = 1'b0;
  assign \A[1][37] [1] = 1'b0;
  assign \A[1][37] [0] = 1'b0;
  assign \A[1][38] [4] = 1'b0;
  assign \A[1][38] [3] = 1'b0;
  assign \A[1][38] [2] = 1'b0;
  assign \A[1][38] [1] = 1'b0;
  assign \A[1][38] [0] = 1'b0;
  assign \A[1][40] [0] = 1'b0;
  assign \A[1][42] [4] = 1'b0;
  assign \A[1][42] [3] = 1'b0;
  assign \A[1][42] [2] = 1'b0;
  assign \A[1][42] [1] = 1'b0;
  assign \A[1][42] [0] = 1'b0;
  assign \A[1][43] [4] = 1'b0;
  assign \A[1][43] [3] = 1'b0;
  assign \A[1][43] [2] = 1'b0;
  assign \A[1][43] [1] = 1'b0;
  assign \A[1][43] [0] = 1'b0;
  assign \A[1][46] [4] = 1'b0;
  assign \A[1][46] [3] = 1'b0;
  assign \A[1][46] [2] = 1'b0;
  assign \A[1][46] [1] = 1'b0;
  assign \A[1][46] [0] = 1'b0;
  assign \A[1][47] [4] = 1'b0;
  assign \A[1][47] [3] = 1'b0;
  assign \A[1][47] [2] = 1'b0;
  assign \A[1][47] [1] = 1'b0;
  assign \A[1][47] [0] = 1'b0;
  assign \A[1][49] [4] = 1'b0;
  assign \A[1][49] [3] = 1'b0;
  assign \A[1][49] [2] = 1'b0;
  assign \A[1][52] [1] = 1'b0;
  assign \A[1][53] [4] = 1'b0;
  assign \A[1][53] [3] = 1'b0;
  assign \A[1][53] [2] = 1'b0;
  assign \A[1][53] [1] = 1'b0;
  assign \A[1][53] [0] = 1'b0;
  assign \A[1][54] [4] = 1'b0;
  assign \A[1][54] [3] = 1'b0;
  assign \A[1][54] [2] = 1'b0;
  assign \A[1][54] [1] = 1'b0;
  assign \A[1][56] [0] = 1'b0;
  assign \A[1][57] [4] = 1'b0;
  assign \A[1][57] [3] = 1'b0;
  assign \A[1][57] [2] = 1'b0;
  assign \A[1][57] [1] = 1'b0;
  assign \A[1][57] [0] = 1'b0;
  assign \A[1][59] [0] = 1'b0;
  assign \A[1][61] [4] = 1'b0;
  assign \A[1][61] [3] = 1'b0;
  assign \A[1][61] [2] = 1'b0;
  assign \A[1][61] [1] = 1'b0;
  assign \A[1][62] [1] = 1'b0;
  assign \A[1][63] [4] = 1'b0;
  assign \A[1][63] [3] = 1'b0;
  assign \A[1][63] [2] = 1'b0;
  assign \A[1][63] [1] = 1'b0;
  assign \A[1][63] [0] = 1'b0;
  assign \A[1][64] [4] = 1'b0;
  assign \A[1][64] [3] = 1'b0;
  assign \A[1][64] [2] = 1'b0;
  assign \A[1][64] [1] = 1'b0;
  assign \A[1][64] [0] = 1'b0;
  assign \A[1][65] [4] = 1'b0;
  assign \A[1][65] [3] = 1'b0;
  assign \A[1][65] [2] = 1'b0;
  assign \A[1][65] [1] = 1'b0;
  assign \A[1][66] [0] = 1'b0;
  assign \A[1][67] [0] = 1'b0;
  assign \A[1][68] [1] = 1'b0;
  assign \A[1][69] [4] = 1'b0;
  assign \A[1][69] [3] = 1'b0;
  assign \A[1][69] [2] = 1'b0;
  assign \A[1][69] [0] = 1'b0;
  assign \A[1][70] [4] = 1'b0;
  assign \A[1][70] [3] = 1'b0;
  assign \A[1][70] [2] = 1'b0;
  assign \A[1][70] [1] = 1'b0;
  assign \A[1][71] [0] = 1'b0;
  assign \A[1][72] [4] = 1'b0;
  assign \A[1][72] [3] = 1'b0;
  assign \A[1][72] [2] = 1'b0;
  assign \A[1][72] [1] = 1'b0;
  assign \A[1][72] [0] = 1'b0;
  assign \A[1][74] [0] = 1'b0;
  assign \A[1][75] [4] = 1'b0;
  assign \A[1][75] [3] = 1'b0;
  assign \A[1][75] [2] = 1'b0;
  assign \A[1][75] [1] = 1'b0;
  assign \A[1][76] [0] = 1'b0;
  assign \A[1][79] [1] = 1'b0;
  assign \A[1][80] [4] = 1'b0;
  assign \A[1][80] [3] = 1'b0;
  assign \A[1][80] [2] = 1'b0;
  assign \A[1][80] [1] = 1'b0;
  assign \A[1][80] [0] = 1'b0;
  assign \A[1][81] [1] = 1'b0;
  assign \A[1][82] [4] = 1'b0;
  assign \A[1][82] [3] = 1'b0;
  assign \A[1][82] [2] = 1'b0;
  assign \A[1][82] [1] = 1'b0;
  assign \A[1][83] [0] = 1'b0;
  assign \A[1][84] [0] = 1'b0;
  assign \A[1][85] [4] = 1'b0;
  assign \A[1][85] [3] = 1'b0;
  assign \A[1][85] [2] = 1'b0;
  assign \A[1][85] [1] = 1'b0;
  assign \A[1][86] [4] = 1'b0;
  assign \A[1][86] [3] = 1'b0;
  assign \A[1][86] [2] = 1'b0;
  assign \A[1][86] [1] = 1'b0;
  assign \A[1][86] [0] = 1'b0;
  assign \A[1][87] [4] = 1'b0;
  assign \A[1][87] [3] = 1'b0;
  assign \A[1][87] [2] = 1'b0;
  assign \A[1][87] [1] = 1'b0;
  assign \A[1][87] [0] = 1'b0;
  assign \A[1][89] [0] = 1'b0;
  assign \A[1][90] [4] = 1'b0;
  assign \A[1][90] [3] = 1'b0;
  assign \A[1][90] [2] = 1'b0;
  assign \A[1][90] [1] = 1'b0;
  assign \A[1][91] [4] = 1'b0;
  assign \A[1][91] [3] = 1'b0;
  assign \A[1][91] [2] = 1'b0;
  assign \A[1][91] [1] = 1'b0;
  assign \A[1][92] [4] = 1'b0;
  assign \A[1][92] [3] = 1'b0;
  assign \A[1][92] [2] = 1'b0;
  assign \A[1][92] [1] = 1'b0;
  assign \A[1][92] [0] = 1'b0;
  assign \A[1][93] [4] = 1'b0;
  assign \A[1][93] [3] = 1'b0;
  assign \A[1][93] [2] = 1'b0;
  assign \A[1][93] [1] = 1'b0;
  assign \A[1][95] [4] = 1'b0;
  assign \A[1][95] [3] = 1'b0;
  assign \A[1][95] [2] = 1'b0;
  assign \A[1][95] [0] = 1'b0;
  assign \A[1][97] [4] = 1'b0;
  assign \A[1][97] [3] = 1'b0;
  assign \A[1][97] [2] = 1'b0;
  assign \A[1][97] [1] = 1'b0;
  assign \A[1][97] [0] = 1'b0;
  assign \A[1][98] [4] = 1'b0;
  assign \A[1][98] [3] = 1'b0;
  assign \A[1][98] [2] = 1'b0;
  assign \A[1][98] [1] = 1'b0;
  assign \A[1][98] [0] = 1'b0;
  assign \A[1][99] [4] = 1'b0;
  assign \A[1][99] [3] = 1'b0;
  assign \A[1][99] [2] = 1'b0;
  assign \A[1][99] [1] = 1'b0;
  assign \A[1][100] [4] = 1'b0;
  assign \A[1][100] [3] = 1'b0;
  assign \A[1][100] [2] = 1'b0;
  assign \A[1][100] [0] = 1'b0;
  assign \A[1][101] [4] = 1'b0;
  assign \A[1][101] [3] = 1'b0;
  assign \A[1][101] [2] = 1'b0;
  assign \A[1][101] [1] = 1'b0;
  assign \A[1][101] [0] = 1'b0;
  assign \A[1][102] [4] = 1'b0;
  assign \A[1][102] [3] = 1'b0;
  assign \A[1][102] [2] = 1'b0;
  assign \A[1][102] [0] = 1'b0;
  assign \A[1][103] [4] = 1'b0;
  assign \A[1][103] [3] = 1'b0;
  assign \A[1][103] [2] = 1'b0;
  assign \A[1][103] [0] = 1'b0;
  assign \A[1][104] [4] = 1'b0;
  assign \A[1][104] [3] = 1'b0;
  assign \A[1][104] [2] = 1'b0;
  assign \A[1][105] [0] = 1'b0;
  assign \A[1][106] [4] = 1'b0;
  assign \A[1][106] [3] = 1'b0;
  assign \A[1][106] [2] = 1'b0;
  assign \A[1][106] [1] = 1'b0;
  assign \A[1][107] [0] = 1'b0;
  assign \A[1][108] [4] = 1'b0;
  assign \A[1][108] [3] = 1'b0;
  assign \A[1][108] [2] = 1'b0;
  assign \A[1][108] [1] = 1'b0;
  assign \A[1][114] [0] = 1'b0;
  assign \A[1][116] [4] = 1'b0;
  assign \A[1][116] [3] = 1'b0;
  assign \A[1][116] [2] = 1'b0;
  assign \A[1][116] [1] = 1'b0;
  assign \A[1][116] [0] = 1'b0;
  assign \A[1][117] [4] = 1'b0;
  assign \A[1][117] [3] = 1'b0;
  assign \A[1][117] [2] = 1'b0;
  assign \A[1][117] [1] = 1'b0;
  assign \A[1][117] [0] = 1'b0;
  assign \A[1][118] [4] = 1'b0;
  assign \A[1][118] [3] = 1'b0;
  assign \A[1][118] [2] = 1'b0;
  assign \A[1][118] [1] = 1'b0;
  assign \A[1][119] [4] = 1'b0;
  assign \A[1][119] [3] = 1'b0;
  assign \A[1][119] [2] = 1'b0;
  assign \A[1][119] [1] = 1'b0;
  assign \A[1][120] [4] = 1'b0;
  assign \A[1][120] [3] = 1'b0;
  assign \A[1][120] [2] = 1'b0;
  assign \A[1][120] [1] = 1'b0;
  assign \A[1][120] [0] = 1'b0;
  assign \A[1][121] [4] = 1'b0;
  assign \A[1][121] [3] = 1'b0;
  assign \A[1][121] [2] = 1'b0;
  assign \A[1][121] [1] = 1'b0;
  assign \A[1][121] [0] = 1'b0;
  assign \A[1][122] [4] = 1'b0;
  assign \A[1][122] [3] = 1'b0;
  assign \A[1][122] [2] = 1'b0;
  assign \A[1][122] [1] = 1'b0;
  assign \A[1][123] [0] = 1'b0;
  assign \A[1][124] [4] = 1'b0;
  assign \A[1][124] [3] = 1'b0;
  assign \A[1][124] [2] = 1'b0;
  assign \A[1][124] [1] = 1'b0;
  assign \A[1][124] [0] = 1'b0;
  assign \A[1][125] [4] = 1'b0;
  assign \A[1][125] [3] = 1'b0;
  assign \A[1][125] [2] = 1'b0;
  assign \A[1][125] [1] = 1'b0;
  assign \A[1][125] [0] = 1'b0;
  assign \A[1][126] [4] = 1'b0;
  assign \A[1][126] [3] = 1'b0;
  assign \A[1][126] [2] = 1'b0;
  assign \A[1][126] [1] = 1'b0;
  assign \A[1][126] [0] = 1'b0;
  assign \A[1][127] [4] = 1'b0;
  assign \A[1][127] [3] = 1'b0;
  assign \A[1][127] [2] = 1'b0;
  assign \A[1][127] [1] = 1'b0;
  assign \A[1][127] [0] = 1'b0;
  assign \A[1][128] [4] = 1'b0;
  assign \A[1][128] [3] = 1'b0;
  assign \A[1][128] [2] = 1'b0;
  assign \A[1][128] [1] = 1'b0;
  assign \A[1][128] [0] = 1'b0;
  assign \A[1][129] [4] = 1'b0;
  assign \A[1][129] [3] = 1'b0;
  assign \A[1][129] [2] = 1'b0;
  assign \A[1][129] [1] = 1'b0;
  assign \A[1][129] [0] = 1'b0;
  assign \A[1][130] [4] = 1'b0;
  assign \A[1][130] [3] = 1'b0;
  assign \A[1][130] [2] = 1'b0;
  assign \A[1][130] [1] = 1'b0;
  assign \A[1][131] [4] = 1'b0;
  assign \A[1][131] [3] = 1'b0;
  assign \A[1][131] [2] = 1'b0;
  assign \A[1][131] [1] = 1'b0;
  assign \A[1][132] [0] = 1'b0;
  assign \A[1][133] [4] = 1'b0;
  assign \A[1][133] [3] = 1'b0;
  assign \A[1][133] [2] = 1'b0;
  assign \A[1][133] [1] = 1'b0;
  assign \A[1][136] [4] = 1'b0;
  assign \A[1][136] [3] = 1'b0;
  assign \A[1][136] [2] = 1'b0;
  assign \A[1][136] [1] = 1'b0;
  assign \A[1][136] [0] = 1'b0;
  assign \A[1][138] [4] = 1'b0;
  assign \A[1][138] [3] = 1'b0;
  assign \A[1][138] [2] = 1'b0;
  assign \A[1][138] [1] = 1'b0;
  assign \A[1][139] [4] = 1'b0;
  assign \A[1][139] [3] = 1'b0;
  assign \A[1][139] [2] = 1'b0;
  assign \A[1][139] [1] = 1'b0;
  assign \A[1][139] [0] = 1'b0;
  assign \A[1][140] [4] = 1'b0;
  assign \A[1][140] [3] = 1'b0;
  assign \A[1][140] [2] = 1'b0;
  assign \A[1][140] [1] = 1'b0;
  assign \A[1][140] [0] = 1'b0;
  assign \A[1][141] [4] = 1'b0;
  assign \A[1][141] [3] = 1'b0;
  assign \A[1][141] [2] = 1'b0;
  assign \A[1][141] [0] = 1'b0;
  assign \A[1][142] [4] = 1'b0;
  assign \A[1][142] [3] = 1'b0;
  assign \A[1][142] [2] = 1'b0;
  assign \A[1][142] [1] = 1'b0;
  assign \A[1][142] [0] = 1'b0;
  assign \A[1][143] [4] = 1'b0;
  assign \A[1][143] [3] = 1'b0;
  assign \A[1][143] [2] = 1'b0;
  assign \A[1][144] [4] = 1'b0;
  assign \A[1][144] [3] = 1'b0;
  assign \A[1][144] [2] = 1'b0;
  assign \A[1][144] [1] = 1'b0;
  assign \A[1][144] [0] = 1'b0;
  assign \A[1][145] [4] = 1'b0;
  assign \A[1][145] [3] = 1'b0;
  assign \A[1][145] [2] = 1'b0;
  assign \A[1][145] [0] = 1'b0;
  assign \A[1][146] [4] = 1'b0;
  assign \A[1][146] [3] = 1'b0;
  assign \A[1][146] [2] = 1'b0;
  assign \A[1][147] [1] = 1'b0;
  assign \A[1][148] [1] = 1'b0;
  assign \A[1][150] [4] = 1'b0;
  assign \A[1][150] [3] = 1'b0;
  assign \A[1][150] [2] = 1'b0;
  assign \A[1][150] [1] = 1'b0;
  assign \A[1][150] [0] = 1'b0;
  assign \A[1][151] [4] = 1'b0;
  assign \A[1][151] [3] = 1'b0;
  assign \A[1][151] [2] = 1'b0;
  assign \A[1][152] [4] = 1'b0;
  assign \A[1][152] [3] = 1'b0;
  assign \A[1][152] [2] = 1'b0;
  assign \A[1][152] [1] = 1'b0;
  assign \A[1][153] [4] = 1'b0;
  assign \A[1][153] [3] = 1'b0;
  assign \A[1][153] [2] = 1'b0;
  assign \A[1][153] [1] = 1'b0;
  assign \A[1][153] [0] = 1'b0;
  assign \A[1][154] [4] = 1'b0;
  assign \A[1][154] [3] = 1'b0;
  assign \A[1][154] [2] = 1'b0;
  assign \A[1][154] [0] = 1'b0;
  assign \A[1][155] [0] = 1'b0;
  assign \A[1][157] [4] = 1'b0;
  assign \A[1][157] [3] = 1'b0;
  assign \A[1][157] [2] = 1'b0;
  assign \A[1][157] [1] = 1'b0;
  assign \A[1][158] [4] = 1'b0;
  assign \A[1][158] [3] = 1'b0;
  assign \A[1][158] [2] = 1'b0;
  assign \A[1][158] [1] = 1'b0;
  assign \A[1][159] [4] = 1'b0;
  assign \A[1][159] [3] = 1'b0;
  assign \A[1][159] [2] = 1'b0;
  assign \A[1][159] [1] = 1'b0;
  assign \A[1][159] [0] = 1'b0;
  assign \A[1][160] [4] = 1'b0;
  assign \A[1][160] [3] = 1'b0;
  assign \A[1][160] [2] = 1'b0;
  assign \A[1][160] [0] = 1'b0;
  assign \A[1][163] [4] = 1'b0;
  assign \A[1][163] [3] = 1'b0;
  assign \A[1][163] [2] = 1'b0;
  assign \A[1][163] [1] = 1'b0;
  assign \A[1][163] [0] = 1'b0;
  assign \A[1][165] [4] = 1'b0;
  assign \A[1][165] [3] = 1'b0;
  assign \A[1][165] [2] = 1'b0;
  assign \A[1][165] [1] = 1'b0;
  assign \A[1][165] [0] = 1'b0;
  assign \A[1][166] [4] = 1'b0;
  assign \A[1][166] [3] = 1'b0;
  assign \A[1][166] [2] = 1'b0;
  assign \A[1][166] [0] = 1'b0;
  assign \A[1][167] [0] = 1'b0;
  assign \A[1][168] [4] = 1'b0;
  assign \A[1][168] [3] = 1'b0;
  assign \A[1][168] [2] = 1'b0;
  assign \A[1][168] [1] = 1'b0;
  assign \A[1][168] [0] = 1'b0;
  assign \A[1][169] [0] = 1'b0;
  assign \A[1][170] [4] = 1'b0;
  assign \A[1][170] [3] = 1'b0;
  assign \A[1][170] [2] = 1'b0;
  assign \A[1][170] [1] = 1'b0;
  assign \A[1][171] [0] = 1'b0;
  assign \A[1][172] [4] = 1'b0;
  assign \A[1][172] [3] = 1'b0;
  assign \A[1][172] [2] = 1'b0;
  assign \A[1][172] [1] = 1'b0;
  assign \A[1][172] [0] = 1'b0;
  assign \A[1][173] [4] = 1'b0;
  assign \A[1][173] [3] = 1'b0;
  assign \A[1][173] [2] = 1'b0;
  assign \A[1][173] [1] = 1'b0;
  assign \A[1][174] [4] = 1'b0;
  assign \A[1][174] [3] = 1'b0;
  assign \A[1][174] [2] = 1'b0;
  assign \A[1][175] [4] = 1'b0;
  assign \A[1][175] [3] = 1'b0;
  assign \A[1][175] [2] = 1'b0;
  assign \A[1][175] [1] = 1'b0;
  assign \A[1][175] [0] = 1'b0;
  assign \A[1][176] [4] = 1'b0;
  assign \A[1][176] [3] = 1'b0;
  assign \A[1][176] [2] = 1'b0;
  assign \A[1][176] [1] = 1'b0;
  assign \A[1][180] [4] = 1'b0;
  assign \A[1][180] [3] = 1'b0;
  assign \A[1][180] [2] = 1'b0;
  assign \A[1][180] [1] = 1'b0;
  assign \A[1][180] [0] = 1'b0;
  assign \A[1][181] [4] = 1'b0;
  assign \A[1][181] [3] = 1'b0;
  assign \A[1][181] [2] = 1'b0;
  assign \A[1][181] [1] = 1'b0;
  assign \A[1][181] [0] = 1'b0;
  assign \A[1][182] [0] = 1'b0;
  assign \A[1][183] [4] = 1'b0;
  assign \A[1][183] [3] = 1'b0;
  assign \A[1][183] [2] = 1'b0;
  assign \A[1][183] [0] = 1'b0;
  assign \A[1][186] [1] = 1'b0;
  assign \A[1][187] [4] = 1'b0;
  assign \A[1][187] [3] = 1'b0;
  assign \A[1][187] [2] = 1'b0;
  assign \A[1][188] [4] = 1'b0;
  assign \A[1][188] [3] = 1'b0;
  assign \A[1][188] [2] = 1'b0;
  assign \A[1][188] [0] = 1'b0;
  assign \A[1][189] [1] = 1'b0;
  assign \A[1][190] [4] = 1'b0;
  assign \A[1][190] [3] = 1'b0;
  assign \A[1][190] [2] = 1'b0;
  assign \A[1][191] [4] = 1'b0;
  assign \A[1][191] [3] = 1'b0;
  assign \A[1][191] [2] = 1'b0;
  assign \A[1][191] [0] = 1'b0;
  assign \A[1][192] [4] = 1'b0;
  assign \A[1][192] [3] = 1'b0;
  assign \A[1][192] [2] = 1'b0;
  assign \A[1][195] [4] = 1'b0;
  assign \A[1][195] [3] = 1'b0;
  assign \A[1][195] [2] = 1'b0;
  assign \A[1][196] [4] = 1'b0;
  assign \A[1][196] [3] = 1'b0;
  assign \A[1][196] [2] = 1'b0;
  assign \A[1][197] [1] = 1'b0;
  assign \A[1][198] [4] = 1'b0;
  assign \A[1][198] [3] = 1'b0;
  assign \A[1][198] [2] = 1'b0;
  assign \A[1][198] [1] = 1'b0;
  assign \A[1][200] [4] = 1'b0;
  assign \A[1][200] [3] = 1'b0;
  assign \A[1][200] [2] = 1'b0;
  assign \A[1][200] [1] = 1'b0;
  assign \A[1][201] [4] = 1'b0;
  assign \A[1][201] [3] = 1'b0;
  assign \A[1][201] [2] = 1'b0;
  assign \A[1][201] [1] = 1'b0;
  assign \A[1][201] [0] = 1'b0;
  assign \A[1][202] [4] = 1'b0;
  assign \A[1][202] [3] = 1'b0;
  assign \A[1][202] [2] = 1'b0;
  assign \A[1][202] [1] = 1'b0;
  assign \A[1][203] [4] = 1'b0;
  assign \A[1][203] [3] = 1'b0;
  assign \A[1][203] [2] = 1'b0;
  assign \A[1][203] [1] = 1'b0;
  assign \A[1][203] [0] = 1'b0;
  assign \A[1][205] [4] = 1'b0;
  assign \A[1][205] [3] = 1'b0;
  assign \A[1][205] [2] = 1'b0;
  assign \A[1][205] [1] = 1'b0;
  assign \A[1][205] [0] = 1'b0;
  assign \A[1][206] [4] = 1'b0;
  assign \A[1][206] [3] = 1'b0;
  assign \A[1][206] [2] = 1'b0;
  assign \A[1][206] [1] = 1'b0;
  assign \A[1][206] [0] = 1'b0;
  assign \A[1][212] [4] = 1'b0;
  assign \A[1][212] [3] = 1'b0;
  assign \A[1][212] [2] = 1'b0;
  assign \A[1][212] [1] = 1'b0;
  assign \A[1][213] [4] = 1'b0;
  assign \A[1][213] [3] = 1'b0;
  assign \A[1][213] [2] = 1'b0;
  assign \A[1][213] [1] = 1'b0;
  assign \A[1][213] [0] = 1'b0;
  assign \A[1][214] [0] = 1'b0;
  assign \A[1][215] [4] = 1'b0;
  assign \A[1][215] [3] = 1'b0;
  assign \A[1][215] [2] = 1'b0;
  assign \A[1][215] [1] = 1'b0;
  assign \A[1][215] [0] = 1'b0;
  assign \A[1][217] [0] = 1'b0;
  assign \A[1][218] [4] = 1'b0;
  assign \A[1][218] [3] = 1'b0;
  assign \A[1][218] [2] = 1'b0;
  assign \A[1][218] [1] = 1'b0;
  assign \A[1][221] [4] = 1'b0;
  assign \A[1][221] [3] = 1'b0;
  assign \A[1][221] [2] = 1'b0;
  assign \A[1][221] [1] = 1'b0;
  assign \A[1][222] [4] = 1'b0;
  assign \A[1][222] [3] = 1'b0;
  assign \A[1][222] [2] = 1'b0;
  assign \A[1][222] [1] = 1'b0;
  assign \A[1][222] [0] = 1'b0;
  assign \A[1][223] [4] = 1'b0;
  assign \A[1][223] [3] = 1'b0;
  assign \A[1][223] [2] = 1'b0;
  assign \A[1][223] [1] = 1'b0;
  assign \A[1][224] [1] = 1'b0;
  assign \A[1][225] [0] = 1'b0;
  assign \A[1][226] [4] = 1'b0;
  assign \A[1][226] [3] = 1'b0;
  assign \A[1][226] [2] = 1'b0;
  assign \A[1][226] [1] = 1'b0;
  assign \A[1][226] [0] = 1'b0;
  assign \A[1][228] [4] = 1'b0;
  assign \A[1][228] [3] = 1'b0;
  assign \A[1][228] [1] = 1'b0;
  assign \A[1][228] [0] = 1'b0;
  assign \A[1][229] [4] = 1'b0;
  assign \A[1][229] [3] = 1'b0;
  assign \A[1][229] [2] = 1'b0;
  assign \A[1][229] [1] = 1'b0;
  assign \A[1][229] [0] = 1'b0;
  assign \A[1][230] [4] = 1'b0;
  assign \A[1][230] [3] = 1'b0;
  assign \A[1][230] [2] = 1'b0;
  assign \A[1][230] [1] = 1'b0;
  assign \A[1][231] [0] = 1'b0;
  assign \A[1][232] [4] = 1'b0;
  assign \A[1][232] [3] = 1'b0;
  assign \A[1][232] [2] = 1'b0;
  assign \A[1][232] [0] = 1'b0;
  assign \A[1][233] [4] = 1'b0;
  assign \A[1][233] [3] = 1'b0;
  assign \A[1][233] [2] = 1'b0;
  assign \A[1][233] [0] = 1'b0;
  assign \A[1][234] [4] = 1'b0;
  assign \A[1][234] [3] = 1'b0;
  assign \A[1][234] [2] = 1'b0;
  assign \A[1][234] [1] = 1'b0;
  assign \A[1][235] [4] = 1'b0;
  assign \A[1][235] [3] = 1'b0;
  assign \A[1][235] [2] = 1'b0;
  assign \A[1][235] [1] = 1'b0;
  assign \A[1][235] [0] = 1'b0;
  assign \A[1][236] [4] = 1'b0;
  assign \A[1][236] [3] = 1'b0;
  assign \A[1][236] [2] = 1'b0;
  assign \A[1][236] [1] = 1'b0;
  assign \A[1][238] [4] = 1'b0;
  assign \A[1][238] [3] = 1'b0;
  assign \A[1][238] [2] = 1'b0;
  assign \A[1][239] [0] = 1'b0;
  assign \A[1][241] [1] = 1'b0;
  assign \A[1][242] [0] = 1'b0;
  assign \A[1][243] [1] = 1'b0;
  assign \A[1][245] [4] = 1'b0;
  assign \A[1][245] [3] = 1'b0;
  assign \A[1][245] [2] = 1'b0;
  assign \A[1][245] [1] = 1'b0;
  assign \A[1][246] [4] = 1'b0;
  assign \A[1][246] [3] = 1'b0;
  assign \A[1][246] [2] = 1'b0;
  assign \A[1][246] [1] = 1'b0;
  assign \A[1][246] [0] = 1'b0;
  assign \A[1][249] [4] = 1'b0;
  assign \A[1][249] [3] = 1'b0;
  assign \A[1][249] [2] = 1'b0;
  assign \A[1][249] [1] = 1'b0;
  assign \A[1][249] [0] = 1'b0;
  assign \A[1][253] [4] = 1'b0;
  assign \A[1][253] [3] = 1'b0;
  assign \A[1][253] [2] = 1'b0;
  assign \A[1][253] [1] = 1'b0;
  assign \A[1][255] [0] = 1'b0;
  assign \A[2][0] [2] = 1'b0;
  assign \A[2][0] [0] = 1'b0;
  assign \A[2][1] [4] = 1'b0;
  assign \A[2][1] [3] = 1'b0;
  assign \A[2][1] [2] = 1'b0;
  assign \A[2][1] [1] = 1'b0;
  assign \A[2][1] [0] = 1'b0;
  assign \A[2][3] [4] = 1'b0;
  assign \A[2][3] [3] = 1'b0;
  assign \A[2][3] [2] = 1'b0;
  assign \A[2][3] [1] = 1'b0;
  assign \A[2][3] [0] = 1'b0;
  assign \A[2][5] [1] = 1'b0;
  assign \A[2][7] [1] = 1'b0;
  assign \A[2][8] [4] = 1'b0;
  assign \A[2][8] [3] = 1'b0;
  assign \A[2][8] [2] = 1'b0;
  assign \A[2][8] [1] = 1'b0;
  assign \A[2][9] [0] = 1'b0;
  assign \A[2][10] [0] = 1'b0;
  assign \A[2][11] [0] = 1'b0;
  assign \A[2][13] [2] = 1'b0;
  assign \A[2][18] [0] = 1'b0;
  assign \A[2][20] [1] = 1'b0;
  assign \A[2][21] [4] = 1'b0;
  assign \A[2][21] [3] = 1'b0;
  assign \A[2][21] [2] = 1'b0;
  assign \A[2][21] [0] = 1'b0;
  assign \A[2][22] [0] = 1'b0;
  assign \A[2][23] [4] = 1'b0;
  assign \A[2][23] [3] = 1'b0;
  assign \A[2][23] [2] = 1'b0;
  assign \A[2][23] [1] = 1'b0;
  assign \A[2][23] [0] = 1'b0;
  assign \A[2][24] [4] = 1'b0;
  assign \A[2][24] [3] = 1'b0;
  assign \A[2][24] [2] = 1'b0;
  assign \A[2][24] [1] = 1'b0;
  assign \A[2][24] [0] = 1'b0;
  assign \A[2][25] [0] = 1'b0;
  assign \A[2][26] [4] = 1'b0;
  assign \A[2][26] [3] = 1'b0;
  assign \A[2][26] [2] = 1'b0;
  assign \A[2][26] [1] = 1'b0;
  assign \A[2][26] [0] = 1'b0;
  assign \A[2][27] [0] = 1'b0;
  assign \A[2][28] [4] = 1'b0;
  assign \A[2][28] [3] = 1'b0;
  assign \A[2][28] [2] = 1'b0;
  assign \A[2][28] [1] = 1'b0;
  assign \A[2][28] [0] = 1'b0;
  assign \A[2][29] [4] = 1'b0;
  assign \A[2][29] [3] = 1'b0;
  assign \A[2][29] [2] = 1'b0;
  assign \A[2][29] [0] = 1'b0;
  assign \A[2][31] [0] = 1'b0;
  assign \A[2][32] [1] = 1'b0;
  assign \A[2][32] [0] = 1'b0;
  assign \A[2][36] [4] = 1'b0;
  assign \A[2][36] [3] = 1'b0;
  assign \A[2][36] [2] = 1'b0;
  assign \A[2][36] [1] = 1'b0;
  assign \A[2][36] [0] = 1'b0;
  assign \A[2][37] [0] = 1'b0;
  assign \A[2][38] [4] = 1'b0;
  assign \A[2][38] [3] = 1'b0;
  assign \A[2][38] [2] = 1'b0;
  assign \A[2][38] [1] = 1'b0;
  assign \A[2][38] [0] = 1'b0;
  assign \A[2][41] [4] = 1'b0;
  assign \A[2][41] [3] = 1'b0;
  assign \A[2][41] [2] = 1'b0;
  assign \A[2][41] [1] = 1'b0;
  assign \A[2][41] [0] = 1'b0;
  assign \A[2][42] [4] = 1'b0;
  assign \A[2][42] [3] = 1'b0;
  assign \A[2][42] [2] = 1'b0;
  assign \A[2][42] [1] = 1'b0;
  assign \A[2][44] [0] = 1'b0;
  assign \A[2][45] [1] = 1'b0;
  assign \A[2][47] [4] = 1'b0;
  assign \A[2][47] [3] = 1'b0;
  assign \A[2][47] [2] = 1'b0;
  assign \A[2][47] [1] = 1'b0;
  assign \A[2][47] [0] = 1'b0;
  assign \A[2][48] [4] = 1'b0;
  assign \A[2][48] [3] = 1'b0;
  assign \A[2][48] [2] = 1'b0;
  assign \A[2][48] [1] = 1'b0;
  assign \A[2][49] [4] = 1'b0;
  assign \A[2][49] [3] = 1'b0;
  assign \A[2][49] [2] = 1'b0;
  assign \A[2][49] [1] = 1'b0;
  assign \A[2][49] [0] = 1'b0;
  assign \A[2][50] [4] = 1'b0;
  assign \A[2][50] [3] = 1'b0;
  assign \A[2][50] [2] = 1'b0;
  assign \A[2][50] [1] = 1'b0;
  assign \A[2][53] [4] = 1'b0;
  assign \A[2][53] [3] = 1'b0;
  assign \A[2][53] [2] = 1'b0;
  assign \A[2][53] [1] = 1'b0;
  assign \A[2][53] [0] = 1'b0;
  assign \A[2][54] [4] = 1'b0;
  assign \A[2][54] [3] = 1'b0;
  assign \A[2][54] [2] = 1'b0;
  assign \A[2][54] [1] = 1'b0;
  assign \A[2][55] [4] = 1'b0;
  assign \A[2][55] [3] = 1'b0;
  assign \A[2][55] [2] = 1'b0;
  assign \A[2][55] [1] = 1'b0;
  assign \A[2][56] [4] = 1'b0;
  assign \A[2][56] [3] = 1'b0;
  assign \A[2][56] [2] = 1'b0;
  assign \A[2][56] [1] = 1'b0;
  assign \A[2][56] [0] = 1'b0;
  assign \A[2][57] [4] = 1'b0;
  assign \A[2][57] [3] = 1'b0;
  assign \A[2][57] [2] = 1'b0;
  assign \A[2][57] [1] = 1'b0;
  assign \A[2][59] [4] = 1'b0;
  assign \A[2][59] [3] = 1'b0;
  assign \A[2][59] [2] = 1'b0;
  assign \A[2][59] [0] = 1'b0;
  assign \A[2][60] [4] = 1'b0;
  assign \A[2][60] [3] = 1'b0;
  assign \A[2][60] [2] = 1'b0;
  assign \A[2][60] [1] = 1'b0;
  assign \A[2][63] [4] = 1'b0;
  assign \A[2][63] [3] = 1'b0;
  assign \A[2][63] [2] = 1'b0;
  assign \A[2][63] [1] = 1'b0;
  assign \A[2][65] [4] = 1'b0;
  assign \A[2][65] [3] = 1'b0;
  assign \A[2][65] [2] = 1'b0;
  assign \A[2][65] [1] = 1'b0;
  assign \A[2][65] [0] = 1'b0;
  assign \A[2][66] [4] = 1'b0;
  assign \A[2][66] [3] = 1'b0;
  assign \A[2][66] [2] = 1'b0;
  assign \A[2][66] [0] = 1'b0;
  assign \A[2][67] [4] = 1'b0;
  assign \A[2][67] [3] = 1'b0;
  assign \A[2][67] [2] = 1'b0;
  assign \A[2][67] [1] = 1'b0;
  assign \A[2][68] [4] = 1'b0;
  assign \A[2][68] [3] = 1'b0;
  assign \A[2][68] [2] = 1'b0;
  assign \A[2][68] [1] = 1'b0;
  assign \A[2][68] [0] = 1'b0;
  assign \A[2][71] [4] = 1'b0;
  assign \A[2][71] [3] = 1'b0;
  assign \A[2][71] [2] = 1'b0;
  assign \A[2][71] [0] = 1'b0;
  assign \A[2][72] [4] = 1'b0;
  assign \A[2][72] [3] = 1'b0;
  assign \A[2][72] [2] = 1'b0;
  assign \A[2][72] [1] = 1'b0;
  assign \A[2][73] [4] = 1'b0;
  assign \A[2][73] [3] = 1'b0;
  assign \A[2][73] [2] = 1'b0;
  assign \A[2][73] [1] = 1'b0;
  assign \A[2][75] [4] = 1'b0;
  assign \A[2][75] [3] = 1'b0;
  assign \A[2][75] [2] = 1'b0;
  assign \A[2][75] [1] = 1'b0;
  assign \A[2][75] [0] = 1'b0;
  assign \A[2][76] [4] = 1'b0;
  assign \A[2][76] [3] = 1'b0;
  assign \A[2][76] [2] = 1'b0;
  assign \A[2][76] [1] = 1'b0;
  assign \A[2][76] [0] = 1'b0;
  assign \A[2][77] [4] = 1'b0;
  assign \A[2][77] [3] = 1'b0;
  assign \A[2][77] [2] = 1'b0;
  assign \A[2][77] [1] = 1'b0;
  assign \A[2][77] [0] = 1'b0;
  assign \A[2][79] [1] = 1'b0;
  assign \A[2][81] [0] = 1'b0;
  assign \A[2][82] [4] = 1'b0;
  assign \A[2][82] [3] = 1'b0;
  assign \A[2][82] [2] = 1'b0;
  assign \A[2][82] [1] = 1'b0;
  assign \A[2][83] [1] = 1'b0;
  assign \A[2][83] [0] = 1'b0;
  assign \A[2][84] [4] = 1'b0;
  assign \A[2][84] [3] = 1'b0;
  assign \A[2][84] [2] = 1'b0;
  assign \A[2][84] [0] = 1'b0;
  assign \A[2][86] [4] = 1'b0;
  assign \A[2][86] [3] = 1'b0;
  assign \A[2][86] [2] = 1'b0;
  assign \A[2][86] [1] = 1'b0;
  assign \A[2][86] [0] = 1'b0;
  assign \A[2][87] [4] = 1'b0;
  assign \A[2][87] [3] = 1'b0;
  assign \A[2][87] [2] = 1'b0;
  assign \A[2][87] [1] = 1'b0;
  assign \A[2][87] [0] = 1'b0;
  assign \A[2][88] [4] = 1'b0;
  assign \A[2][88] [3] = 1'b0;
  assign \A[2][88] [2] = 1'b0;
  assign \A[2][89] [4] = 1'b0;
  assign \A[2][89] [3] = 1'b0;
  assign \A[2][89] [2] = 1'b0;
  assign \A[2][89] [1] = 1'b0;
  assign \A[2][89] [0] = 1'b0;
  assign \A[2][90] [4] = 1'b0;
  assign \A[2][90] [3] = 1'b0;
  assign \A[2][90] [2] = 1'b0;
  assign \A[2][91] [0] = 1'b0;
  assign \A[2][92] [4] = 1'b0;
  assign \A[2][92] [3] = 1'b0;
  assign \A[2][92] [2] = 1'b0;
  assign \A[2][92] [1] = 1'b0;
  assign \A[2][92] [0] = 1'b0;
  assign \A[2][93] [4] = 1'b0;
  assign \A[2][93] [3] = 1'b0;
  assign \A[2][93] [2] = 1'b0;
  assign \A[2][93] [1] = 1'b0;
  assign \A[2][94] [0] = 1'b0;
  assign \A[2][96] [0] = 1'b0;
  assign \A[2][97] [4] = 1'b0;
  assign \A[2][97] [3] = 1'b0;
  assign \A[2][97] [2] = 1'b0;
  assign \A[2][98] [0] = 1'b0;
  assign \A[2][99] [4] = 1'b0;
  assign \A[2][99] [3] = 1'b0;
  assign \A[2][99] [2] = 1'b0;
  assign \A[2][99] [1] = 1'b0;
  assign \A[2][100] [4] = 1'b0;
  assign \A[2][100] [3] = 1'b0;
  assign \A[2][100] [2] = 1'b0;
  assign \A[2][100] [1] = 1'b0;
  assign \A[2][101] [0] = 1'b0;
  assign \A[2][103] [4] = 1'b0;
  assign \A[2][103] [3] = 1'b0;
  assign \A[2][103] [2] = 1'b0;
  assign \A[2][103] [1] = 1'b0;
  assign \A[2][103] [0] = 1'b0;
  assign \A[2][104] [4] = 1'b0;
  assign \A[2][104] [3] = 1'b0;
  assign \A[2][104] [2] = 1'b0;
  assign \A[2][104] [0] = 1'b0;
  assign \A[2][106] [4] = 1'b0;
  assign \A[2][106] [3] = 1'b0;
  assign \A[2][106] [2] = 1'b0;
  assign \A[2][106] [1] = 1'b0;
  assign \A[2][107] [4] = 1'b0;
  assign \A[2][107] [3] = 1'b0;
  assign \A[2][107] [2] = 1'b0;
  assign \A[2][107] [1] = 1'b0;
  assign \A[2][107] [0] = 1'b0;
  assign \A[2][108] [4] = 1'b0;
  assign \A[2][108] [3] = 1'b0;
  assign \A[2][108] [2] = 1'b0;
  assign \A[2][108] [1] = 1'b0;
  assign \A[2][110] [4] = 1'b0;
  assign \A[2][110] [3] = 1'b0;
  assign \A[2][110] [2] = 1'b0;
  assign \A[2][111] [4] = 1'b0;
  assign \A[2][111] [3] = 1'b0;
  assign \A[2][111] [2] = 1'b0;
  assign \A[2][111] [1] = 1'b0;
  assign \A[2][111] [0] = 1'b0;
  assign \A[2][112] [4] = 1'b0;
  assign \A[2][112] [3] = 1'b0;
  assign \A[2][112] [2] = 1'b0;
  assign \A[2][113] [0] = 1'b0;
  assign \A[2][114] [4] = 1'b0;
  assign \A[2][114] [3] = 1'b0;
  assign \A[2][114] [2] = 1'b0;
  assign \A[2][114] [0] = 1'b0;
  assign \A[2][116] [4] = 1'b0;
  assign \A[2][116] [3] = 1'b0;
  assign \A[2][116] [2] = 1'b0;
  assign \A[2][116] [1] = 1'b0;
  assign \A[2][117] [4] = 1'b0;
  assign \A[2][117] [3] = 1'b0;
  assign \A[2][117] [2] = 1'b0;
  assign \A[2][117] [1] = 1'b0;
  assign \A[2][118] [0] = 1'b0;
  assign \A[2][119] [4] = 1'b0;
  assign \A[2][119] [3] = 1'b0;
  assign \A[2][119] [2] = 1'b0;
  assign \A[2][119] [0] = 1'b0;
  assign \A[2][120] [4] = 1'b0;
  assign \A[2][120] [3] = 1'b0;
  assign \A[2][120] [2] = 1'b0;
  assign \A[2][120] [1] = 1'b0;
  assign \A[2][120] [0] = 1'b0;
  assign \A[2][121] [4] = 1'b0;
  assign \A[2][121] [3] = 1'b0;
  assign \A[2][121] [2] = 1'b0;
  assign \A[2][121] [0] = 1'b0;
  assign \A[2][122] [4] = 1'b0;
  assign \A[2][122] [3] = 1'b0;
  assign \A[2][122] [2] = 1'b0;
  assign \A[2][122] [1] = 1'b0;
  assign \A[2][123] [4] = 1'b0;
  assign \A[2][123] [3] = 1'b0;
  assign \A[2][123] [2] = 1'b0;
  assign \A[2][123] [1] = 1'b0;
  assign \A[2][123] [0] = 1'b0;
  assign \A[2][124] [4] = 1'b0;
  assign \A[2][124] [3] = 1'b0;
  assign \A[2][124] [2] = 1'b0;
  assign \A[2][124] [1] = 1'b0;
  assign \A[2][125] [4] = 1'b0;
  assign \A[2][125] [3] = 1'b0;
  assign \A[2][125] [2] = 1'b0;
  assign \A[2][125] [1] = 1'b0;
  assign \A[2][126] [4] = 1'b0;
  assign \A[2][126] [3] = 1'b0;
  assign \A[2][126] [2] = 1'b0;
  assign \A[2][126] [1] = 1'b0;
  assign \A[2][126] [0] = 1'b0;
  assign \A[2][129] [4] = 1'b0;
  assign \A[2][129] [3] = 1'b0;
  assign \A[2][129] [2] = 1'b0;
  assign \A[2][130] [4] = 1'b0;
  assign \A[2][130] [3] = 1'b0;
  assign \A[2][130] [2] = 1'b0;
  assign \A[2][130] [1] = 1'b0;
  assign \A[2][131] [4] = 1'b0;
  assign \A[2][131] [3] = 1'b0;
  assign \A[2][131] [2] = 1'b0;
  assign \A[2][131] [0] = 1'b0;
  assign \A[2][132] [4] = 1'b0;
  assign \A[2][132] [3] = 1'b0;
  assign \A[2][132] [2] = 1'b0;
  assign \A[2][132] [1] = 1'b0;
  assign \A[2][133] [4] = 1'b0;
  assign \A[2][133] [3] = 1'b0;
  assign \A[2][133] [2] = 1'b0;
  assign \A[2][133] [1] = 1'b0;
  assign \A[2][133] [0] = 1'b0;
  assign \A[2][134] [0] = 1'b0;
  assign \A[2][135] [4] = 1'b0;
  assign \A[2][135] [3] = 1'b0;
  assign \A[2][135] [2] = 1'b0;
  assign \A[2][135] [1] = 1'b0;
  assign \A[2][135] [0] = 1'b0;
  assign \A[2][137] [4] = 1'b0;
  assign \A[2][137] [3] = 1'b0;
  assign \A[2][137] [1] = 1'b0;
  assign \A[2][137] [0] = 1'b0;
  assign \A[2][138] [4] = 1'b0;
  assign \A[2][138] [3] = 1'b0;
  assign \A[2][138] [2] = 1'b0;
  assign \A[2][138] [1] = 1'b0;
  assign \A[2][139] [4] = 1'b0;
  assign \A[2][139] [3] = 1'b0;
  assign \A[2][139] [2] = 1'b0;
  assign \A[2][139] [1] = 1'b0;
  assign \A[2][139] [0] = 1'b0;
  assign \A[2][140] [0] = 1'b0;
  assign \A[2][141] [4] = 1'b0;
  assign \A[2][141] [3] = 1'b0;
  assign \A[2][141] [2] = 1'b0;
  assign \A[2][141] [1] = 1'b0;
  assign \A[2][142] [4] = 1'b0;
  assign \A[2][142] [3] = 1'b0;
  assign \A[2][142] [2] = 1'b0;
  assign \A[2][142] [1] = 1'b0;
  assign \A[2][142] [0] = 1'b0;
  assign \A[2][144] [1] = 1'b0;
  assign \A[2][145] [4] = 1'b0;
  assign \A[2][145] [3] = 1'b0;
  assign \A[2][145] [2] = 1'b0;
  assign \A[2][146] [1] = 1'b0;
  assign \A[2][148] [4] = 1'b0;
  assign \A[2][148] [3] = 1'b0;
  assign \A[2][148] [2] = 1'b0;
  assign \A[2][148] [0] = 1'b0;
  assign \A[2][149] [4] = 1'b0;
  assign \A[2][149] [3] = 1'b0;
  assign \A[2][149] [2] = 1'b0;
  assign \A[2][149] [1] = 1'b0;
  assign \A[2][150] [4] = 1'b0;
  assign \A[2][150] [3] = 1'b0;
  assign \A[2][150] [2] = 1'b0;
  assign \A[2][150] [1] = 1'b0;
  assign \A[2][150] [0] = 1'b0;
  assign \A[2][151] [4] = 1'b0;
  assign \A[2][151] [3] = 1'b0;
  assign \A[2][151] [2] = 1'b0;
  assign \A[2][151] [1] = 1'b0;
  assign \A[2][151] [0] = 1'b0;
  assign \A[2][152] [4] = 1'b0;
  assign \A[2][152] [3] = 1'b0;
  assign \A[2][152] [2] = 1'b0;
  assign \A[2][152] [1] = 1'b0;
  assign \A[2][152] [0] = 1'b0;
  assign \A[2][154] [4] = 1'b0;
  assign \A[2][154] [3] = 1'b0;
  assign \A[2][154] [2] = 1'b0;
  assign \A[2][154] [1] = 1'b0;
  assign \A[2][155] [4] = 1'b0;
  assign \A[2][155] [3] = 1'b0;
  assign \A[2][155] [2] = 1'b0;
  assign \A[2][155] [0] = 1'b0;
  assign \A[2][156] [4] = 1'b0;
  assign \A[2][156] [3] = 1'b0;
  assign \A[2][156] [2] = 1'b0;
  assign \A[2][156] [1] = 1'b0;
  assign \A[2][157] [4] = 1'b0;
  assign \A[2][157] [3] = 1'b0;
  assign \A[2][157] [2] = 1'b0;
  assign \A[2][157] [1] = 1'b0;
  assign \A[2][157] [0] = 1'b0;
  assign \A[2][158] [4] = 1'b0;
  assign \A[2][158] [3] = 1'b0;
  assign \A[2][158] [2] = 1'b0;
  assign \A[2][158] [0] = 1'b0;
  assign \A[2][159] [1] = 1'b0;
  assign \A[2][160] [4] = 1'b0;
  assign \A[2][160] [3] = 1'b0;
  assign \A[2][160] [2] = 1'b0;
  assign \A[2][160] [1] = 1'b0;
  assign \A[2][160] [0] = 1'b0;
  assign \A[2][161] [4] = 1'b0;
  assign \A[2][161] [3] = 1'b0;
  assign \A[2][161] [1] = 1'b0;
  assign \A[2][161] [0] = 1'b0;
  assign \A[2][162] [4] = 1'b0;
  assign \A[2][162] [3] = 1'b0;
  assign \A[2][162] [2] = 1'b0;
  assign \A[2][162] [1] = 1'b0;
  assign \A[2][162] [0] = 1'b0;
  assign \A[2][163] [4] = 1'b0;
  assign \A[2][163] [3] = 1'b0;
  assign \A[2][163] [2] = 1'b0;
  assign \A[2][163] [1] = 1'b0;
  assign \A[2][165] [4] = 1'b0;
  assign \A[2][165] [3] = 1'b0;
  assign \A[2][165] [2] = 1'b0;
  assign \A[2][165] [1] = 1'b0;
  assign \A[2][166] [4] = 1'b0;
  assign \A[2][166] [3] = 1'b0;
  assign \A[2][166] [2] = 1'b0;
  assign \A[2][166] [1] = 1'b0;
  assign \A[2][167] [4] = 1'b0;
  assign \A[2][167] [3] = 1'b0;
  assign \A[2][167] [2] = 1'b0;
  assign \A[2][168] [4] = 1'b0;
  assign \A[2][168] [3] = 1'b0;
  assign \A[2][168] [2] = 1'b0;
  assign \A[2][168] [0] = 1'b0;
  assign \A[2][169] [4] = 1'b0;
  assign \A[2][169] [3] = 1'b0;
  assign \A[2][169] [2] = 1'b0;
  assign \A[2][170] [4] = 1'b0;
  assign \A[2][170] [3] = 1'b0;
  assign \A[2][170] [2] = 1'b0;
  assign \A[2][170] [1] = 1'b0;
  assign \A[2][170] [0] = 1'b0;
  assign \A[2][171] [4] = 1'b0;
  assign \A[2][171] [3] = 1'b0;
  assign \A[2][171] [2] = 1'b0;
  assign \A[2][171] [1] = 1'b0;
  assign \A[2][172] [4] = 1'b0;
  assign \A[2][172] [3] = 1'b0;
  assign \A[2][172] [2] = 1'b0;
  assign \A[2][172] [0] = 1'b0;
  assign \A[2][174] [0] = 1'b0;
  assign \A[2][175] [4] = 1'b0;
  assign \A[2][175] [3] = 1'b0;
  assign \A[2][175] [2] = 1'b0;
  assign \A[2][175] [1] = 1'b0;
  assign \A[2][177] [0] = 1'b0;
  assign \A[2][180] [0] = 1'b0;
  assign \A[2][181] [4] = 1'b0;
  assign \A[2][181] [3] = 1'b0;
  assign \A[2][181] [2] = 1'b0;
  assign \A[2][182] [4] = 1'b0;
  assign \A[2][182] [3] = 1'b0;
  assign \A[2][182] [2] = 1'b0;
  assign \A[2][182] [1] = 1'b0;
  assign \A[2][183] [4] = 1'b0;
  assign \A[2][183] [3] = 1'b0;
  assign \A[2][183] [2] = 1'b0;
  assign \A[2][183] [1] = 1'b0;
  assign \A[2][184] [4] = 1'b0;
  assign \A[2][184] [3] = 1'b0;
  assign \A[2][184] [2] = 1'b0;
  assign \A[2][184] [1] = 1'b0;
  assign \A[2][184] [0] = 1'b0;
  assign \A[2][185] [4] = 1'b0;
  assign \A[2][185] [3] = 1'b0;
  assign \A[2][185] [2] = 1'b0;
  assign \A[2][185] [1] = 1'b0;
  assign \A[2][185] [0] = 1'b0;
  assign \A[2][186] [4] = 1'b0;
  assign \A[2][186] [3] = 1'b0;
  assign \A[2][186] [2] = 1'b0;
  assign \A[2][186] [1] = 1'b0;
  assign \A[2][187] [4] = 1'b0;
  assign \A[2][187] [3] = 1'b0;
  assign \A[2][187] [2] = 1'b0;
  assign \A[2][187] [1] = 1'b0;
  assign \A[2][188] [4] = 1'b0;
  assign \A[2][188] [3] = 1'b0;
  assign \A[2][188] [2] = 1'b0;
  assign \A[2][188] [1] = 1'b0;
  assign \A[2][191] [4] = 1'b0;
  assign \A[2][191] [3] = 1'b0;
  assign \A[2][191] [2] = 1'b0;
  assign \A[2][191] [1] = 1'b0;
  assign \A[2][192] [4] = 1'b0;
  assign \A[2][192] [3] = 1'b0;
  assign \A[2][192] [2] = 1'b0;
  assign \A[2][192] [0] = 1'b0;
  assign \A[2][194] [4] = 1'b0;
  assign \A[2][194] [3] = 1'b0;
  assign \A[2][194] [2] = 1'b0;
  assign \A[2][194] [0] = 1'b0;
  assign \A[2][195] [4] = 1'b0;
  assign \A[2][195] [3] = 1'b0;
  assign \A[2][195] [2] = 1'b0;
  assign \A[2][195] [0] = 1'b0;
  assign \A[2][196] [4] = 1'b0;
  assign \A[2][196] [3] = 1'b0;
  assign \A[2][196] [2] = 1'b0;
  assign \A[2][196] [1] = 1'b0;
  assign \A[2][197] [4] = 1'b0;
  assign \A[2][197] [3] = 1'b0;
  assign \A[2][197] [2] = 1'b0;
  assign \A[2][197] [1] = 1'b0;
  assign \A[2][198] [4] = 1'b0;
  assign \A[2][198] [3] = 1'b0;
  assign \A[2][198] [2] = 1'b0;
  assign \A[2][198] [1] = 1'b0;
  assign \A[2][198] [0] = 1'b0;
  assign \A[2][199] [4] = 1'b0;
  assign \A[2][199] [3] = 1'b0;
  assign \A[2][199] [2] = 1'b0;
  assign \A[2][199] [1] = 1'b0;
  assign \A[2][199] [0] = 1'b0;
  assign \A[2][200] [0] = 1'b0;
  assign \A[2][201] [4] = 1'b0;
  assign \A[2][201] [3] = 1'b0;
  assign \A[2][201] [2] = 1'b0;
  assign \A[2][202] [4] = 1'b0;
  assign \A[2][202] [3] = 1'b0;
  assign \A[2][202] [2] = 1'b0;
  assign \A[2][202] [1] = 1'b0;
  assign \A[2][202] [0] = 1'b0;
  assign \A[2][203] [4] = 1'b0;
  assign \A[2][203] [3] = 1'b0;
  assign \A[2][203] [2] = 1'b0;
  assign \A[2][204] [4] = 1'b0;
  assign \A[2][204] [3] = 1'b0;
  assign \A[2][204] [2] = 1'b0;
  assign \A[2][204] [1] = 1'b0;
  assign \A[2][205] [4] = 1'b0;
  assign \A[2][205] [3] = 1'b0;
  assign \A[2][205] [2] = 1'b0;
  assign \A[2][205] [1] = 1'b0;
  assign \A[2][206] [4] = 1'b0;
  assign \A[2][206] [3] = 1'b0;
  assign \A[2][206] [2] = 1'b0;
  assign \A[2][206] [1] = 1'b0;
  assign \A[2][208] [4] = 1'b0;
  assign \A[2][208] [3] = 1'b0;
  assign \A[2][208] [2] = 1'b0;
  assign \A[2][208] [1] = 1'b0;
  assign \A[2][208] [0] = 1'b0;
  assign \A[2][209] [4] = 1'b0;
  assign \A[2][209] [3] = 1'b0;
  assign \A[2][209] [2] = 1'b0;
  assign \A[2][209] [1] = 1'b0;
  assign \A[2][210] [0] = 1'b0;
  assign \A[2][211] [4] = 1'b0;
  assign \A[2][211] [3] = 1'b0;
  assign \A[2][211] [2] = 1'b0;
  assign \A[2][211] [0] = 1'b0;
  assign \A[2][212] [4] = 1'b0;
  assign \A[2][212] [3] = 1'b0;
  assign \A[2][212] [2] = 1'b0;
  assign \A[2][212] [1] = 1'b0;
  assign \A[2][212] [0] = 1'b0;
  assign \A[2][214] [1] = 1'b0;
  assign \A[2][215] [0] = 1'b0;
  assign \A[2][217] [0] = 1'b0;
  assign \A[2][219] [0] = 1'b0;
  assign \A[2][220] [4] = 1'b0;
  assign \A[2][220] [3] = 1'b0;
  assign \A[2][220] [2] = 1'b0;
  assign \A[2][221] [4] = 1'b0;
  assign \A[2][221] [3] = 1'b0;
  assign \A[2][221] [2] = 1'b0;
  assign \A[2][221] [1] = 1'b0;
  assign \A[2][223] [4] = 1'b0;
  assign \A[2][223] [3] = 1'b0;
  assign \A[2][223] [2] = 1'b0;
  assign \A[2][223] [1] = 1'b0;
  assign \A[2][223] [0] = 1'b0;
  assign \A[2][226] [4] = 1'b0;
  assign \A[2][226] [3] = 1'b0;
  assign \A[2][226] [2] = 1'b0;
  assign \A[2][226] [1] = 1'b0;
  assign \A[2][228] [1] = 1'b0;
  assign \A[2][228] [0] = 1'b0;
  assign \A[2][229] [4] = 1'b0;
  assign \A[2][229] [3] = 1'b0;
  assign \A[2][229] [2] = 1'b0;
  assign \A[2][229] [1] = 1'b0;
  assign \A[2][229] [0] = 1'b0;
  assign \A[2][231] [0] = 1'b0;
  assign \A[2][233] [0] = 1'b0;
  assign \A[2][234] [1] = 1'b0;
  assign \A[2][234] [0] = 1'b0;
  assign \A[2][236] [1] = 1'b0;
  assign \A[2][236] [0] = 1'b0;
  assign \A[2][237] [4] = 1'b0;
  assign \A[2][237] [3] = 1'b0;
  assign \A[2][237] [2] = 1'b0;
  assign \A[2][237] [1] = 1'b0;
  assign \A[2][237] [0] = 1'b0;
  assign \A[2][239] [4] = 1'b0;
  assign \A[2][239] [3] = 1'b0;
  assign \A[2][239] [2] = 1'b0;
  assign \A[2][239] [1] = 1'b0;
  assign \A[2][241] [4] = 1'b0;
  assign \A[2][241] [3] = 1'b0;
  assign \A[2][241] [2] = 1'b0;
  assign \A[2][241] [1] = 1'b0;
  assign \A[2][241] [0] = 1'b0;
  assign \A[2][242] [0] = 1'b0;
  assign \A[2][243] [1] = 1'b0;
  assign \A[2][244] [1] = 1'b0;
  assign \A[2][244] [0] = 1'b0;
  assign \A[2][246] [4] = 1'b0;
  assign \A[2][246] [3] = 1'b0;
  assign \A[2][246] [2] = 1'b0;
  assign \A[2][246] [1] = 1'b0;
  assign \A[2][246] [0] = 1'b0;
  assign \A[2][247] [1] = 1'b0;
  assign \A[2][248] [4] = 1'b0;
  assign \A[2][248] [3] = 1'b0;
  assign \A[2][248] [2] = 1'b0;
  assign \A[2][248] [1] = 1'b0;
  assign \A[2][248] [0] = 1'b0;
  assign \A[2][249] [4] = 1'b0;
  assign \A[2][249] [3] = 1'b0;
  assign \A[2][249] [2] = 1'b0;
  assign \A[2][249] [1] = 1'b0;
  assign \A[2][249] [0] = 1'b0;
  assign \A[2][250] [4] = 1'b0;
  assign \A[2][250] [3] = 1'b0;
  assign \A[2][250] [2] = 1'b0;
  assign \A[2][250] [1] = 1'b0;
  assign \A[2][251] [4] = 1'b0;
  assign \A[2][251] [3] = 1'b0;
  assign \A[2][251] [2] = 1'b0;
  assign \A[2][251] [0] = 1'b0;
  assign \A[2][254] [0] = 1'b0;
  assign \A[2][255] [4] = 1'b0;
  assign \A[2][255] [3] = 1'b0;
  assign \A[2][255] [2] = 1'b0;
  assign \A[2][255] [1] = 1'b0;
  assign \A[2][255] [0] = 1'b0;
  assign \A[3][0] [4] = 1'b0;
  assign \A[3][0] [3] = 1'b0;
  assign \A[3][0] [2] = 1'b0;
  assign \A[3][0] [1] = 1'b0;
  assign \A[3][0] [0] = 1'b0;
  assign \A[3][1] [4] = 1'b0;
  assign \A[3][1] [3] = 1'b0;
  assign \A[3][1] [2] = 1'b0;
  assign \A[3][1] [1] = 1'b0;
  assign \A[3][3] [4] = 1'b0;
  assign \A[3][3] [3] = 1'b0;
  assign \A[3][3] [2] = 1'b0;
  assign \A[3][3] [1] = 1'b0;
  assign \A[3][3] [0] = 1'b0;
  assign \A[3][4] [4] = 1'b0;
  assign \A[3][4] [3] = 1'b0;
  assign \A[3][4] [2] = 1'b0;
  assign \A[3][4] [1] = 1'b0;
  assign \A[3][5] [0] = 1'b0;
  assign \A[3][6] [1] = 1'b0;
  assign \A[3][8] [4] = 1'b0;
  assign \A[3][8] [3] = 1'b0;
  assign \A[3][8] [2] = 1'b0;
  assign \A[3][8] [0] = 1'b0;
  assign \A[3][9] [0] = 1'b0;
  assign \A[3][12] [4] = 1'b0;
  assign \A[3][12] [3] = 1'b0;
  assign \A[3][12] [2] = 1'b0;
  assign \A[3][12] [1] = 1'b0;
  assign \A[3][12] [0] = 1'b0;
  assign \A[3][14] [4] = 1'b0;
  assign \A[3][14] [3] = 1'b0;
  assign \A[3][14] [2] = 1'b0;
  assign \A[3][14] [0] = 1'b0;
  assign \A[3][15] [4] = 1'b0;
  assign \A[3][15] [3] = 1'b0;
  assign \A[3][15] [2] = 1'b0;
  assign \A[3][17] [4] = 1'b0;
  assign \A[3][17] [3] = 1'b0;
  assign \A[3][17] [2] = 1'b0;
  assign \A[3][17] [1] = 1'b0;
  assign \A[3][17] [0] = 1'b0;
  assign \A[3][18] [0] = 1'b0;
  assign \A[3][19] [4] = 1'b0;
  assign \A[3][19] [3] = 1'b0;
  assign \A[3][19] [2] = 1'b0;
  assign \A[3][19] [1] = 1'b0;
  assign \A[3][19] [0] = 1'b0;
  assign \A[3][20] [0] = 1'b0;
  assign \A[3][21] [4] = 1'b0;
  assign \A[3][21] [3] = 1'b0;
  assign \A[3][21] [2] = 1'b0;
  assign \A[3][21] [1] = 1'b0;
  assign \A[3][21] [0] = 1'b0;
  assign \A[3][22] [4] = 1'b0;
  assign \A[3][22] [3] = 1'b0;
  assign \A[3][22] [2] = 1'b0;
  assign \A[3][22] [1] = 1'b0;
  assign \A[3][22] [0] = 1'b0;
  assign \A[3][23] [4] = 1'b0;
  assign \A[3][23] [3] = 1'b0;
  assign \A[3][23] [2] = 1'b0;
  assign \A[3][23] [1] = 1'b0;
  assign \A[3][23] [0] = 1'b0;
  assign \A[3][24] [4] = 1'b0;
  assign \A[3][24] [3] = 1'b0;
  assign \A[3][24] [2] = 1'b0;
  assign \A[3][24] [1] = 1'b0;
  assign \A[3][24] [0] = 1'b0;
  assign \A[3][25] [4] = 1'b0;
  assign \A[3][25] [3] = 1'b0;
  assign \A[3][25] [2] = 1'b0;
  assign \A[3][25] [1] = 1'b0;
  assign \A[3][26] [0] = 1'b0;
  assign \A[3][27] [4] = 1'b0;
  assign \A[3][27] [3] = 1'b0;
  assign \A[3][27] [2] = 1'b0;
  assign \A[3][27] [1] = 1'b0;
  assign \A[3][27] [0] = 1'b0;
  assign \A[3][28] [4] = 1'b0;
  assign \A[3][28] [3] = 1'b0;
  assign \A[3][28] [2] = 1'b0;
  assign \A[3][28] [0] = 1'b0;
  assign \A[3][29] [0] = 1'b0;
  assign \A[3][30] [4] = 1'b0;
  assign \A[3][30] [3] = 1'b0;
  assign \A[3][30] [2] = 1'b0;
  assign \A[3][30] [1] = 1'b0;
  assign \A[3][30] [0] = 1'b0;
  assign \A[3][31] [4] = 1'b0;
  assign \A[3][31] [3] = 1'b0;
  assign \A[3][31] [2] = 1'b0;
  assign \A[3][31] [1] = 1'b0;
  assign \A[3][32] [4] = 1'b0;
  assign \A[3][32] [3] = 1'b0;
  assign \A[3][32] [2] = 1'b0;
  assign \A[3][32] [1] = 1'b0;
  assign \A[3][32] [0] = 1'b0;
  assign \A[3][33] [0] = 1'b0;
  assign \A[3][38] [4] = 1'b0;
  assign \A[3][38] [3] = 1'b0;
  assign \A[3][38] [2] = 1'b0;
  assign \A[3][38] [1] = 1'b0;
  assign \A[3][39] [0] = 1'b0;
  assign \A[3][40] [4] = 1'b0;
  assign \A[3][40] [3] = 1'b0;
  assign \A[3][40] [2] = 1'b0;
  assign \A[3][40] [1] = 1'b0;
  assign \A[3][40] [0] = 1'b0;
  assign \A[3][42] [4] = 1'b0;
  assign \A[3][42] [3] = 1'b0;
  assign \A[3][42] [2] = 1'b0;
  assign \A[3][42] [1] = 1'b0;
  assign \A[3][42] [0] = 1'b0;
  assign \A[3][44] [4] = 1'b0;
  assign \A[3][44] [3] = 1'b0;
  assign \A[3][44] [2] = 1'b0;
  assign \A[3][44] [1] = 1'b0;
  assign \A[3][45] [4] = 1'b0;
  assign \A[3][45] [3] = 1'b0;
  assign \A[3][45] [2] = 1'b0;
  assign \A[3][45] [0] = 1'b0;
  assign \A[3][46] [4] = 1'b0;
  assign \A[3][46] [3] = 1'b0;
  assign \A[3][46] [2] = 1'b0;
  assign \A[3][46] [1] = 1'b0;
  assign \A[3][47] [0] = 1'b0;
  assign \A[3][51] [4] = 1'b0;
  assign \A[3][51] [3] = 1'b0;
  assign \A[3][51] [2] = 1'b0;
  assign \A[3][51] [1] = 1'b0;
  assign \A[3][51] [0] = 1'b0;
  assign \A[3][53] [4] = 1'b0;
  assign \A[3][53] [3] = 1'b0;
  assign \A[3][53] [2] = 1'b0;
  assign \A[3][53] [0] = 1'b0;
  assign \A[3][54] [1] = 1'b0;
  assign \A[3][56] [4] = 1'b0;
  assign \A[3][56] [3] = 1'b0;
  assign \A[3][56] [2] = 1'b0;
  assign \A[3][57] [4] = 1'b0;
  assign \A[3][57] [3] = 1'b0;
  assign \A[3][57] [2] = 1'b0;
  assign \A[3][57] [1] = 1'b0;
  assign \A[3][58] [4] = 1'b0;
  assign \A[3][58] [3] = 1'b0;
  assign \A[3][58] [2] = 1'b0;
  assign \A[3][58] [1] = 1'b0;
  assign \A[3][59] [4] = 1'b0;
  assign \A[3][59] [3] = 1'b0;
  assign \A[3][59] [2] = 1'b0;
  assign \A[3][59] [1] = 1'b0;
  assign \A[3][59] [0] = 1'b0;
  assign \A[3][60] [4] = 1'b0;
  assign \A[3][60] [3] = 1'b0;
  assign \A[3][60] [2] = 1'b0;
  assign \A[3][60] [1] = 1'b0;
  assign \A[3][60] [0] = 1'b0;
  assign \A[3][61] [4] = 1'b0;
  assign \A[3][61] [3] = 1'b0;
  assign \A[3][61] [2] = 1'b0;
  assign \A[3][61] [1] = 1'b0;
  assign \A[3][62] [4] = 1'b0;
  assign \A[3][62] [3] = 1'b0;
  assign \A[3][62] [2] = 1'b0;
  assign \A[3][62] [1] = 1'b0;
  assign \A[3][62] [0] = 1'b0;
  assign \A[3][63] [4] = 1'b0;
  assign \A[3][63] [3] = 1'b0;
  assign \A[3][63] [2] = 1'b0;
  assign \A[3][63] [1] = 1'b0;
  assign \A[3][63] [0] = 1'b0;
  assign \A[3][64] [4] = 1'b0;
  assign \A[3][64] [3] = 1'b0;
  assign \A[3][64] [2] = 1'b0;
  assign \A[3][64] [1] = 1'b0;
  assign \A[3][65] [4] = 1'b0;
  assign \A[3][65] [3] = 1'b0;
  assign \A[3][65] [2] = 1'b0;
  assign \A[3][65] [0] = 1'b0;
  assign \A[3][68] [4] = 1'b0;
  assign \A[3][68] [3] = 1'b0;
  assign \A[3][68] [2] = 1'b0;
  assign \A[3][68] [1] = 1'b0;
  assign \A[3][69] [4] = 1'b0;
  assign \A[3][69] [3] = 1'b0;
  assign \A[3][69] [2] = 1'b0;
  assign \A[3][69] [0] = 1'b0;
  assign \A[3][70] [4] = 1'b0;
  assign \A[3][70] [3] = 1'b0;
  assign \A[3][70] [2] = 1'b0;
  assign \A[3][71] [4] = 1'b0;
  assign \A[3][71] [3] = 1'b0;
  assign \A[3][71] [2] = 1'b0;
  assign \A[3][71] [1] = 1'b0;
  assign \A[3][71] [0] = 1'b0;
  assign \A[3][72] [4] = 1'b0;
  assign \A[3][72] [3] = 1'b0;
  assign \A[3][72] [2] = 1'b0;
  assign \A[3][73] [0] = 1'b0;
  assign \A[3][74] [1] = 1'b0;
  assign \A[3][74] [0] = 1'b0;
  assign \A[3][75] [4] = 1'b0;
  assign \A[3][75] [3] = 1'b0;
  assign \A[3][75] [2] = 1'b0;
  assign \A[3][75] [1] = 1'b0;
  assign \A[3][75] [0] = 1'b0;
  assign \A[3][76] [4] = 1'b0;
  assign \A[3][76] [3] = 1'b0;
  assign \A[3][76] [2] = 1'b0;
  assign \A[3][76] [0] = 1'b0;
  assign \A[3][77] [4] = 1'b0;
  assign \A[3][77] [3] = 1'b0;
  assign \A[3][77] [2] = 1'b0;
  assign \A[3][77] [1] = 1'b0;
  assign \A[3][78] [0] = 1'b0;
  assign \A[3][79] [4] = 1'b0;
  assign \A[3][79] [3] = 1'b0;
  assign \A[3][79] [2] = 1'b0;
  assign \A[3][79] [0] = 1'b0;
  assign \A[3][81] [4] = 1'b0;
  assign \A[3][81] [3] = 1'b0;
  assign \A[3][81] [2] = 1'b0;
  assign \A[3][81] [1] = 1'b0;
  assign \A[3][82] [4] = 1'b0;
  assign \A[3][82] [3] = 1'b0;
  assign \A[3][82] [2] = 1'b0;
  assign \A[3][82] [1] = 1'b0;
  assign \A[3][82] [0] = 1'b0;
  assign \A[3][85] [4] = 1'b0;
  assign \A[3][85] [3] = 1'b0;
  assign \A[3][85] [2] = 1'b0;
  assign \A[3][85] [0] = 1'b0;
  assign \A[3][86] [4] = 1'b0;
  assign \A[3][86] [3] = 1'b0;
  assign \A[3][86] [2] = 1'b0;
  assign \A[3][86] [1] = 1'b0;
  assign \A[3][87] [4] = 1'b0;
  assign \A[3][87] [3] = 1'b0;
  assign \A[3][87] [2] = 1'b0;
  assign \A[3][87] [1] = 1'b0;
  assign \A[3][88] [4] = 1'b0;
  assign \A[3][88] [3] = 1'b0;
  assign \A[3][88] [2] = 1'b0;
  assign \A[3][88] [1] = 1'b0;
  assign \A[3][88] [0] = 1'b0;
  assign \A[3][89] [0] = 1'b0;
  assign \A[3][90] [4] = 1'b0;
  assign \A[3][90] [3] = 1'b0;
  assign \A[3][90] [2] = 1'b0;
  assign \A[3][90] [1] = 1'b0;
  assign \A[3][91] [4] = 1'b0;
  assign \A[3][91] [3] = 1'b0;
  assign \A[3][91] [2] = 1'b0;
  assign \A[3][91] [0] = 1'b0;
  assign \A[3][94] [4] = 1'b0;
  assign \A[3][94] [3] = 1'b0;
  assign \A[3][94] [2] = 1'b0;
  assign \A[3][94] [1] = 1'b0;
  assign \A[3][94] [0] = 1'b0;
  assign \A[3][97] [4] = 1'b0;
  assign \A[3][97] [3] = 1'b0;
  assign \A[3][97] [2] = 1'b0;
  assign \A[3][97] [1] = 1'b0;
  assign \A[3][97] [0] = 1'b0;
  assign \A[3][100] [0] = 1'b0;
  assign \A[3][102] [4] = 1'b0;
  assign \A[3][102] [3] = 1'b0;
  assign \A[3][102] [2] = 1'b0;
  assign \A[3][102] [0] = 1'b0;
  assign \A[3][103] [4] = 1'b0;
  assign \A[3][103] [3] = 1'b0;
  assign \A[3][103] [2] = 1'b0;
  assign \A[3][103] [1] = 1'b0;
  assign \A[3][103] [0] = 1'b0;
  assign \A[3][104] [4] = 1'b0;
  assign \A[3][104] [3] = 1'b0;
  assign \A[3][104] [2] = 1'b0;
  assign \A[3][104] [1] = 1'b0;
  assign \A[3][106] [4] = 1'b0;
  assign \A[3][106] [3] = 1'b0;
  assign \A[3][106] [2] = 1'b0;
  assign \A[3][106] [0] = 1'b0;
  assign \A[3][107] [4] = 1'b0;
  assign \A[3][107] [3] = 1'b0;
  assign \A[3][107] [2] = 1'b0;
  assign \A[3][107] [1] = 1'b0;
  assign \A[3][107] [0] = 1'b0;
  assign \A[3][108] [4] = 1'b0;
  assign \A[3][108] [3] = 1'b0;
  assign \A[3][108] [1] = 1'b0;
  assign \A[3][108] [0] = 1'b0;
  assign \A[3][109] [4] = 1'b0;
  assign \A[3][109] [3] = 1'b0;
  assign \A[3][109] [2] = 1'b0;
  assign \A[3][110] [1] = 1'b0;
  assign \A[3][112] [4] = 1'b0;
  assign \A[3][112] [3] = 1'b0;
  assign \A[3][112] [2] = 1'b0;
  assign \A[3][112] [1] = 1'b0;
  assign \A[3][112] [0] = 1'b0;
  assign \A[3][113] [4] = 1'b0;
  assign \A[3][113] [3] = 1'b0;
  assign \A[3][113] [2] = 1'b0;
  assign \A[3][113] [1] = 1'b0;
  assign \A[3][114] [1] = 1'b0;
  assign \A[3][116] [4] = 1'b0;
  assign \A[3][116] [3] = 1'b0;
  assign \A[3][116] [2] = 1'b0;
  assign \A[3][116] [1] = 1'b0;
  assign \A[3][116] [0] = 1'b0;
  assign \A[3][118] [4] = 1'b0;
  assign \A[3][118] [3] = 1'b0;
  assign \A[3][118] [2] = 1'b0;
  assign \A[3][118] [1] = 1'b0;
  assign \A[3][118] [0] = 1'b0;
  assign \A[3][120] [0] = 1'b0;
  assign \A[3][121] [4] = 1'b0;
  assign \A[3][121] [3] = 1'b0;
  assign \A[3][121] [2] = 1'b0;
  assign \A[3][121] [1] = 1'b0;
  assign \A[3][122] [4] = 1'b0;
  assign \A[3][122] [3] = 1'b0;
  assign \A[3][122] [2] = 1'b0;
  assign \A[3][122] [1] = 1'b0;
  assign \A[3][122] [0] = 1'b0;
  assign \A[3][123] [4] = 1'b0;
  assign \A[3][123] [3] = 1'b0;
  assign \A[3][123] [2] = 1'b0;
  assign \A[3][123] [0] = 1'b0;
  assign \A[3][124] [4] = 1'b0;
  assign \A[3][124] [3] = 1'b0;
  assign \A[3][124] [2] = 1'b0;
  assign \A[3][124] [1] = 1'b0;
  assign \A[3][124] [0] = 1'b0;
  assign \A[3][125] [4] = 1'b0;
  assign \A[3][125] [3] = 1'b0;
  assign \A[3][125] [2] = 1'b0;
  assign \A[3][125] [1] = 1'b0;
  assign \A[3][125] [0] = 1'b0;
  assign \A[3][126] [4] = 1'b0;
  assign \A[3][126] [3] = 1'b0;
  assign \A[3][126] [2] = 1'b0;
  assign \A[3][126] [1] = 1'b0;
  assign \A[3][126] [0] = 1'b0;
  assign \A[3][127] [4] = 1'b0;
  assign \A[3][127] [3] = 1'b0;
  assign \A[3][127] [2] = 1'b0;
  assign \A[3][127] [1] = 1'b0;
  assign \A[3][129] [0] = 1'b0;
  assign \A[3][130] [0] = 1'b0;
  assign \A[3][131] [4] = 1'b0;
  assign \A[3][131] [3] = 1'b0;
  assign \A[3][131] [2] = 1'b0;
  assign \A[3][131] [1] = 1'b0;
  assign \A[3][131] [0] = 1'b0;
  assign \A[3][133] [4] = 1'b0;
  assign \A[3][133] [3] = 1'b0;
  assign \A[3][133] [2] = 1'b0;
  assign \A[3][133] [1] = 1'b0;
  assign \A[3][133] [0] = 1'b0;
  assign \A[3][134] [4] = 1'b0;
  assign \A[3][134] [3] = 1'b0;
  assign \A[3][134] [2] = 1'b0;
  assign \A[3][134] [1] = 1'b0;
  assign \A[3][134] [0] = 1'b0;
  assign \A[3][135] [0] = 1'b0;
  assign \A[3][136] [4] = 1'b0;
  assign \A[3][136] [3] = 1'b0;
  assign \A[3][136] [2] = 1'b0;
  assign \A[3][136] [0] = 1'b0;
  assign \A[3][137] [4] = 1'b0;
  assign \A[3][137] [3] = 1'b0;
  assign \A[3][137] [2] = 1'b0;
  assign \A[3][137] [1] = 1'b0;
  assign \A[3][138] [4] = 1'b0;
  assign \A[3][138] [3] = 1'b0;
  assign \A[3][138] [2] = 1'b0;
  assign \A[3][138] [1] = 1'b0;
  assign \A[3][138] [0] = 1'b0;
  assign \A[3][139] [4] = 1'b0;
  assign \A[3][139] [3] = 1'b0;
  assign \A[3][139] [2] = 1'b0;
  assign \A[3][139] [1] = 1'b0;
  assign \A[3][140] [0] = 1'b0;
  assign \A[3][141] [0] = 1'b0;
  assign \A[3][143] [4] = 1'b0;
  assign \A[3][143] [3] = 1'b0;
  assign \A[3][143] [2] = 1'b0;
  assign \A[3][143] [1] = 1'b0;
  assign \A[3][143] [0] = 1'b0;
  assign \A[3][144] [0] = 1'b0;
  assign \A[3][145] [4] = 1'b0;
  assign \A[3][145] [3] = 1'b0;
  assign \A[3][145] [2] = 1'b0;
  assign \A[3][145] [0] = 1'b0;
  assign \A[3][148] [4] = 1'b0;
  assign \A[3][148] [3] = 1'b0;
  assign \A[3][148] [2] = 1'b0;
  assign \A[3][148] [1] = 1'b0;
  assign \A[3][149] [4] = 1'b0;
  assign \A[3][149] [3] = 1'b0;
  assign \A[3][149] [2] = 1'b0;
  assign \A[3][150] [4] = 1'b0;
  assign \A[3][150] [3] = 1'b0;
  assign \A[3][150] [2] = 1'b0;
  assign \A[3][150] [0] = 1'b0;
  assign \A[3][152] [4] = 1'b0;
  assign \A[3][152] [3] = 1'b0;
  assign \A[3][152] [2] = 1'b0;
  assign \A[3][152] [1] = 1'b0;
  assign \A[3][153] [4] = 1'b0;
  assign \A[3][153] [3] = 1'b0;
  assign \A[3][153] [2] = 1'b0;
  assign \A[3][153] [1] = 1'b0;
  assign \A[3][153] [0] = 1'b0;
  assign \A[3][154] [4] = 1'b0;
  assign \A[3][154] [3] = 1'b0;
  assign \A[3][154] [2] = 1'b0;
  assign \A[3][154] [0] = 1'b0;
  assign \A[3][158] [0] = 1'b0;
  assign \A[3][159] [0] = 1'b0;
  assign \A[3][161] [1] = 1'b0;
  assign \A[3][162] [4] = 1'b0;
  assign \A[3][162] [3] = 1'b0;
  assign \A[3][162] [2] = 1'b0;
  assign \A[3][162] [1] = 1'b0;
  assign \A[3][163] [4] = 1'b0;
  assign \A[3][163] [3] = 1'b0;
  assign \A[3][163] [2] = 1'b0;
  assign \A[3][163] [1] = 1'b0;
  assign \A[3][163] [0] = 1'b0;
  assign \A[3][164] [4] = 1'b0;
  assign \A[3][164] [3] = 1'b0;
  assign \A[3][164] [2] = 1'b0;
  assign \A[3][164] [1] = 1'b0;
  assign \A[3][166] [4] = 1'b0;
  assign \A[3][166] [3] = 1'b0;
  assign \A[3][166] [2] = 1'b0;
  assign \A[3][166] [1] = 1'b0;
  assign \A[3][166] [0] = 1'b0;
  assign \A[3][167] [4] = 1'b0;
  assign \A[3][167] [3] = 1'b0;
  assign \A[3][167] [2] = 1'b0;
  assign \A[3][167] [1] = 1'b0;
  assign \A[3][167] [0] = 1'b0;
  assign \A[3][169] [4] = 1'b0;
  assign \A[3][169] [3] = 1'b0;
  assign \A[3][169] [2] = 1'b0;
  assign \A[3][169] [1] = 1'b0;
  assign \A[3][169] [0] = 1'b0;
  assign \A[3][170] [1] = 1'b0;
  assign \A[3][171] [4] = 1'b0;
  assign \A[3][171] [3] = 1'b0;
  assign \A[3][171] [2] = 1'b0;
  assign \A[3][171] [1] = 1'b0;
  assign \A[3][171] [0] = 1'b0;
  assign \A[3][172] [4] = 1'b0;
  assign \A[3][172] [3] = 1'b0;
  assign \A[3][172] [2] = 1'b0;
  assign \A[3][172] [1] = 1'b0;
  assign \A[3][173] [4] = 1'b0;
  assign \A[3][173] [3] = 1'b0;
  assign \A[3][173] [2] = 1'b0;
  assign \A[3][173] [1] = 1'b0;
  assign \A[3][173] [0] = 1'b0;
  assign \A[3][174] [0] = 1'b0;
  assign \A[3][175] [1] = 1'b0;
  assign \A[3][176] [4] = 1'b0;
  assign \A[3][176] [3] = 1'b0;
  assign \A[3][176] [2] = 1'b0;
  assign \A[3][176] [1] = 1'b0;
  assign \A[3][176] [0] = 1'b0;
  assign \A[3][177] [4] = 1'b0;
  assign \A[3][177] [3] = 1'b0;
  assign \A[3][177] [2] = 1'b0;
  assign \A[3][177] [1] = 1'b0;
  assign \A[3][177] [0] = 1'b0;
  assign \A[3][178] [4] = 1'b0;
  assign \A[3][178] [3] = 1'b0;
  assign \A[3][178] [2] = 1'b0;
  assign \A[3][178] [1] = 1'b0;
  assign \A[3][179] [4] = 1'b0;
  assign \A[3][179] [3] = 1'b0;
  assign \A[3][179] [2] = 1'b0;
  assign \A[3][179] [0] = 1'b0;
  assign \A[3][180] [4] = 1'b0;
  assign \A[3][180] [3] = 1'b0;
  assign \A[3][180] [2] = 1'b0;
  assign \A[3][180] [0] = 1'b0;
  assign \A[3][181] [4] = 1'b0;
  assign \A[3][181] [3] = 1'b0;
  assign \A[3][181] [2] = 1'b0;
  assign \A[3][181] [1] = 1'b0;
  assign \A[3][182] [4] = 1'b0;
  assign \A[3][182] [3] = 1'b0;
  assign \A[3][182] [2] = 1'b0;
  assign \A[3][182] [1] = 1'b0;
  assign \A[3][182] [0] = 1'b0;
  assign \A[3][184] [0] = 1'b0;
  assign \A[3][186] [4] = 1'b0;
  assign \A[3][186] [3] = 1'b0;
  assign \A[3][186] [2] = 1'b0;
  assign \A[3][186] [0] = 1'b0;
  assign \A[3][187] [4] = 1'b0;
  assign \A[3][187] [3] = 1'b0;
  assign \A[3][187] [2] = 1'b0;
  assign \A[3][187] [0] = 1'b0;
  assign \A[3][189] [4] = 1'b0;
  assign \A[3][189] [3] = 1'b0;
  assign \A[3][189] [2] = 1'b0;
  assign \A[3][189] [1] = 1'b0;
  assign \A[3][189] [0] = 1'b0;
  assign \A[3][190] [4] = 1'b0;
  assign \A[3][190] [3] = 1'b0;
  assign \A[3][190] [2] = 1'b0;
  assign \A[3][190] [1] = 1'b0;
  assign \A[3][190] [0] = 1'b0;
  assign \A[3][191] [0] = 1'b0;
  assign \A[3][192] [4] = 1'b0;
  assign \A[3][192] [3] = 1'b0;
  assign \A[3][192] [2] = 1'b0;
  assign \A[3][192] [1] = 1'b0;
  assign \A[3][193] [4] = 1'b0;
  assign \A[3][193] [3] = 1'b0;
  assign \A[3][193] [2] = 1'b0;
  assign \A[3][193] [1] = 1'b0;
  assign \A[3][193] [0] = 1'b0;
  assign \A[3][194] [0] = 1'b0;
  assign \A[3][195] [4] = 1'b0;
  assign \A[3][195] [3] = 1'b0;
  assign \A[3][195] [2] = 1'b0;
  assign \A[3][195] [0] = 1'b0;
  assign \A[3][196] [4] = 1'b0;
  assign \A[3][196] [3] = 1'b0;
  assign \A[3][196] [2] = 1'b0;
  assign \A[3][196] [1] = 1'b0;
  assign \A[3][196] [0] = 1'b0;
  assign \A[3][197] [4] = 1'b0;
  assign \A[3][197] [3] = 1'b0;
  assign \A[3][197] [2] = 1'b0;
  assign \A[3][197] [0] = 1'b0;
  assign \A[3][198] [1] = 1'b0;
  assign \A[3][199] [4] = 1'b0;
  assign \A[3][199] [3] = 1'b0;
  assign \A[3][199] [2] = 1'b0;
  assign \A[3][199] [1] = 1'b0;
  assign \A[3][199] [0] = 1'b0;
  assign \A[3][201] [4] = 1'b0;
  assign \A[3][201] [3] = 1'b0;
  assign \A[3][201] [2] = 1'b0;
  assign \A[3][201] [1] = 1'b0;
  assign \A[3][202] [4] = 1'b0;
  assign \A[3][202] [3] = 1'b0;
  assign \A[3][202] [2] = 1'b0;
  assign \A[3][202] [1] = 1'b0;
  assign \A[3][202] [0] = 1'b0;
  assign \A[3][203] [0] = 1'b0;
  assign \A[3][204] [4] = 1'b0;
  assign \A[3][204] [3] = 1'b0;
  assign \A[3][204] [2] = 1'b0;
  assign \A[3][204] [1] = 1'b0;
  assign \A[3][206] [0] = 1'b0;
  assign \A[3][207] [4] = 1'b0;
  assign \A[3][207] [3] = 1'b0;
  assign \A[3][207] [2] = 1'b0;
  assign \A[3][207] [1] = 1'b0;
  assign \A[3][207] [0] = 1'b0;
  assign \A[3][208] [4] = 1'b0;
  assign \A[3][208] [3] = 1'b0;
  assign \A[3][208] [2] = 1'b0;
  assign \A[3][208] [1] = 1'b0;
  assign \A[3][208] [0] = 1'b0;
  assign \A[3][211] [4] = 1'b0;
  assign \A[3][211] [3] = 1'b0;
  assign \A[3][211] [2] = 1'b0;
  assign \A[3][211] [0] = 1'b0;
  assign \A[3][213] [4] = 1'b0;
  assign \A[3][213] [3] = 1'b0;
  assign \A[3][213] [2] = 1'b0;
  assign \A[3][213] [1] = 1'b0;
  assign \A[3][213] [0] = 1'b0;
  assign \A[3][214] [0] = 1'b0;
  assign \A[3][216] [4] = 1'b0;
  assign \A[3][216] [3] = 1'b0;
  assign \A[3][216] [2] = 1'b0;
  assign \A[3][216] [0] = 1'b0;
  assign \A[3][217] [4] = 1'b0;
  assign \A[3][217] [3] = 1'b0;
  assign \A[3][217] [2] = 1'b0;
  assign \A[3][217] [1] = 1'b0;
  assign \A[3][217] [0] = 1'b0;
  assign \A[3][223] [4] = 1'b0;
  assign \A[3][223] [3] = 1'b0;
  assign \A[3][223] [2] = 1'b0;
  assign \A[3][223] [1] = 1'b0;
  assign \A[3][224] [4] = 1'b0;
  assign \A[3][224] [3] = 1'b0;
  assign \A[3][224] [2] = 1'b0;
  assign \A[3][224] [1] = 1'b0;
  assign \A[3][225] [4] = 1'b0;
  assign \A[3][225] [3] = 1'b0;
  assign \A[3][225] [2] = 1'b0;
  assign \A[3][225] [1] = 1'b0;
  assign \A[3][227] [4] = 1'b0;
  assign \A[3][227] [3] = 1'b0;
  assign \A[3][227] [2] = 1'b0;
  assign \A[3][227] [1] = 1'b0;
  assign \A[3][227] [0] = 1'b0;
  assign \A[3][228] [4] = 1'b0;
  assign \A[3][228] [3] = 1'b0;
  assign \A[3][228] [2] = 1'b0;
  assign \A[3][228] [1] = 1'b0;
  assign \A[3][228] [0] = 1'b0;
  assign \A[3][230] [0] = 1'b0;
  assign \A[3][231] [4] = 1'b0;
  assign \A[3][231] [3] = 1'b0;
  assign \A[3][231] [2] = 1'b0;
  assign \A[3][231] [1] = 1'b0;
  assign \A[3][231] [0] = 1'b0;
  assign \A[3][232] [4] = 1'b0;
  assign \A[3][232] [3] = 1'b0;
  assign \A[3][232] [2] = 1'b0;
  assign \A[3][232] [1] = 1'b0;
  assign \A[3][232] [0] = 1'b0;
  assign \A[3][233] [4] = 1'b0;
  assign \A[3][233] [3] = 1'b0;
  assign \A[3][233] [2] = 1'b0;
  assign \A[3][233] [1] = 1'b0;
  assign \A[3][234] [4] = 1'b0;
  assign \A[3][234] [3] = 1'b0;
  assign \A[3][234] [2] = 1'b0;
  assign \A[3][234] [1] = 1'b0;
  assign \A[3][234] [0] = 1'b0;
  assign \A[3][235] [4] = 1'b0;
  assign \A[3][235] [3] = 1'b0;
  assign \A[3][235] [2] = 1'b0;
  assign \A[3][235] [1] = 1'b0;
  assign \A[3][236] [4] = 1'b0;
  assign \A[3][236] [3] = 1'b0;
  assign \A[3][236] [2] = 1'b0;
  assign \A[3][236] [1] = 1'b0;
  assign \A[3][236] [0] = 1'b0;
  assign \A[3][237] [4] = 1'b0;
  assign \A[3][237] [3] = 1'b0;
  assign \A[3][237] [2] = 1'b0;
  assign \A[3][237] [1] = 1'b0;
  assign \A[3][237] [0] = 1'b0;
  assign \A[3][240] [4] = 1'b0;
  assign \A[3][240] [3] = 1'b0;
  assign \A[3][240] [2] = 1'b0;
  assign \A[3][240] [0] = 1'b0;
  assign \A[3][241] [4] = 1'b0;
  assign \A[3][241] [3] = 1'b0;
  assign \A[3][241] [2] = 1'b0;
  assign \A[3][241] [1] = 1'b0;
  assign \A[3][241] [0] = 1'b0;
  assign \A[3][242] [1] = 1'b0;
  assign \A[3][243] [4] = 1'b0;
  assign \A[3][243] [3] = 1'b0;
  assign \A[3][243] [2] = 1'b0;
  assign \A[3][243] [0] = 1'b0;
  assign \A[3][244] [4] = 1'b0;
  assign \A[3][244] [3] = 1'b0;
  assign \A[3][244] [2] = 1'b0;
  assign \A[3][244] [0] = 1'b0;
  assign \A[3][245] [4] = 1'b0;
  assign \A[3][245] [3] = 1'b0;
  assign \A[3][245] [2] = 1'b0;
  assign \A[3][245] [1] = 1'b0;
  assign \A[3][245] [0] = 1'b0;
  assign \A[3][247] [4] = 1'b0;
  assign \A[3][247] [3] = 1'b0;
  assign \A[3][247] [2] = 1'b0;
  assign \A[3][247] [1] = 1'b0;
  assign \A[3][249] [4] = 1'b0;
  assign \A[3][249] [3] = 1'b0;
  assign \A[3][249] [2] = 1'b0;
  assign \A[3][249] [1] = 1'b0;
  assign \A[3][250] [4] = 1'b0;
  assign \A[3][250] [3] = 1'b0;
  assign \A[3][250] [2] = 1'b0;
  assign \A[3][250] [1] = 1'b0;
  assign \A[3][250] [0] = 1'b0;
  assign \A[3][251] [0] = 1'b0;
  assign \A[3][252] [4] = 1'b0;
  assign \A[3][252] [3] = 1'b0;
  assign \A[3][252] [2] = 1'b0;
  assign \A[3][252] [1] = 1'b0;
  assign \A[3][252] [0] = 1'b0;
  assign \A[3][253] [4] = 1'b0;
  assign \A[3][253] [3] = 1'b0;
  assign \A[3][253] [2] = 1'b0;
  assign \A[3][253] [1] = 1'b0;
  assign \A[3][253] [0] = 1'b0;
  assign \A[3][254] [4] = 1'b0;
  assign \A[3][254] [3] = 1'b0;
  assign \A[3][254] [2] = 1'b0;
  assign \A[3][254] [1] = 1'b0;
  assign \A[3][254] [0] = 1'b0;
  assign \A[4][2] [4] = 1'b0;
  assign \A[4][2] [3] = 1'b0;
  assign \A[4][2] [2] = 1'b0;
  assign \A[4][2] [1] = 1'b0;
  assign \A[4][2] [0] = 1'b0;
  assign \A[4][3] [4] = 1'b0;
  assign \A[4][3] [3] = 1'b0;
  assign \A[4][3] [2] = 1'b0;
  assign \A[4][3] [1] = 1'b0;
  assign \A[4][4] [4] = 1'b0;
  assign \A[4][4] [3] = 1'b0;
  assign \A[4][4] [2] = 1'b0;
  assign \A[4][4] [1] = 1'b0;
  assign \A[4][4] [0] = 1'b0;
  assign \A[4][5] [0] = 1'b0;
  assign \A[4][6] [0] = 1'b0;
  assign \A[4][8] [4] = 1'b0;
  assign \A[4][8] [3] = 1'b0;
  assign \A[4][8] [2] = 1'b0;
  assign \A[4][8] [1] = 1'b0;
  assign \A[4][11] [1] = 1'b0;
  assign \A[4][12] [4] = 1'b0;
  assign \A[4][12] [3] = 1'b0;
  assign \A[4][12] [2] = 1'b0;
  assign \A[4][12] [1] = 1'b0;
  assign \A[4][12] [0] = 1'b0;
  assign \A[4][13] [4] = 1'b0;
  assign \A[4][13] [3] = 1'b0;
  assign \A[4][13] [2] = 1'b0;
  assign \A[4][13] [1] = 1'b0;
  assign \A[4][13] [0] = 1'b0;
  assign \A[4][14] [4] = 1'b0;
  assign \A[4][14] [3] = 1'b0;
  assign \A[4][14] [2] = 1'b0;
  assign \A[4][14] [1] = 1'b0;
  assign \A[4][15] [4] = 1'b0;
  assign \A[4][15] [3] = 1'b0;
  assign \A[4][15] [2] = 1'b0;
  assign \A[4][15] [1] = 1'b0;
  assign \A[4][17] [4] = 1'b0;
  assign \A[4][17] [3] = 1'b0;
  assign \A[4][17] [2] = 1'b0;
  assign \A[4][17] [1] = 1'b0;
  assign \A[4][17] [0] = 1'b0;
  assign \A[4][18] [4] = 1'b0;
  assign \A[4][18] [3] = 1'b0;
  assign \A[4][18] [2] = 1'b0;
  assign \A[4][18] [1] = 1'b0;
  assign \A[4][18] [0] = 1'b0;
  assign \A[4][21] [4] = 1'b0;
  assign \A[4][21] [3] = 1'b0;
  assign \A[4][21] [2] = 1'b0;
  assign \A[4][21] [1] = 1'b0;
  assign \A[4][22] [4] = 1'b0;
  assign \A[4][22] [3] = 1'b0;
  assign \A[4][22] [2] = 1'b0;
  assign \A[4][22] [1] = 1'b0;
  assign \A[4][22] [0] = 1'b0;
  assign \A[4][23] [0] = 1'b0;
  assign \A[4][24] [4] = 1'b0;
  assign \A[4][24] [3] = 1'b0;
  assign \A[4][24] [2] = 1'b0;
  assign \A[4][24] [1] = 1'b0;
  assign \A[4][26] [1] = 1'b0;
  assign \A[4][27] [4] = 1'b0;
  assign \A[4][27] [3] = 1'b0;
  assign \A[4][27] [2] = 1'b0;
  assign \A[4][27] [1] = 1'b0;
  assign \A[4][27] [0] = 1'b0;
  assign \A[4][29] [4] = 1'b0;
  assign \A[4][29] [3] = 1'b0;
  assign \A[4][29] [2] = 1'b0;
  assign \A[4][29] [0] = 1'b0;
  assign \A[4][30] [4] = 1'b0;
  assign \A[4][30] [3] = 1'b0;
  assign \A[4][30] [2] = 1'b0;
  assign \A[4][31] [1] = 1'b0;
  assign \A[4][32] [0] = 1'b0;
  assign \A[4][33] [0] = 1'b0;
  assign \A[4][34] [0] = 1'b0;
  assign \A[4][36] [4] = 1'b0;
  assign \A[4][36] [3] = 1'b0;
  assign \A[4][36] [2] = 1'b0;
  assign \A[4][36] [1] = 1'b0;
  assign \A[4][36] [0] = 1'b0;
  assign \A[4][37] [1] = 1'b0;
  assign \A[4][38] [4] = 1'b0;
  assign \A[4][38] [3] = 1'b0;
  assign \A[4][38] [2] = 1'b0;
  assign \A[4][38] [1] = 1'b0;
  assign \A[4][38] [0] = 1'b0;
  assign \A[4][40] [0] = 1'b0;
  assign \A[4][41] [4] = 1'b0;
  assign \A[4][41] [3] = 1'b0;
  assign \A[4][41] [2] = 1'b0;
  assign \A[4][41] [1] = 1'b0;
  assign \A[4][41] [0] = 1'b0;
  assign \A[4][42] [1] = 1'b0;
  assign \A[4][43] [0] = 1'b0;
  assign \A[4][44] [4] = 1'b0;
  assign \A[4][44] [3] = 1'b0;
  assign \A[4][44] [1] = 1'b0;
  assign \A[4][44] [0] = 1'b0;
  assign \A[4][45] [4] = 1'b0;
  assign \A[4][45] [3] = 1'b0;
  assign \A[4][45] [2] = 1'b0;
  assign \A[4][45] [1] = 1'b0;
  assign \A[4][45] [0] = 1'b0;
  assign \A[4][46] [4] = 1'b0;
  assign \A[4][46] [3] = 1'b0;
  assign \A[4][46] [2] = 1'b0;
  assign \A[4][46] [1] = 1'b0;
  assign \A[4][47] [4] = 1'b0;
  assign \A[4][47] [3] = 1'b0;
  assign \A[4][47] [2] = 1'b0;
  assign \A[4][47] [1] = 1'b0;
  assign \A[4][47] [0] = 1'b0;
  assign \A[4][49] [4] = 1'b0;
  assign \A[4][49] [3] = 1'b0;
  assign \A[4][49] [2] = 1'b0;
  assign \A[4][49] [0] = 1'b0;
  assign \A[4][50] [4] = 1'b0;
  assign \A[4][50] [3] = 1'b0;
  assign \A[4][50] [2] = 1'b0;
  assign \A[4][50] [1] = 1'b0;
  assign \A[4][50] [0] = 1'b0;
  assign \A[4][52] [0] = 1'b0;
  assign \A[4][55] [1] = 1'b0;
  assign \A[4][55] [0] = 1'b0;
  assign \A[4][56] [4] = 1'b0;
  assign \A[4][56] [3] = 1'b0;
  assign \A[4][56] [2] = 1'b0;
  assign \A[4][57] [4] = 1'b0;
  assign \A[4][57] [3] = 1'b0;
  assign \A[4][57] [2] = 1'b0;
  assign \A[4][57] [1] = 1'b0;
  assign \A[4][58] [4] = 1'b0;
  assign \A[4][58] [3] = 1'b0;
  assign \A[4][58] [2] = 1'b0;
  assign \A[4][58] [1] = 1'b0;
  assign \A[4][61] [4] = 1'b0;
  assign \A[4][61] [3] = 1'b0;
  assign \A[4][61] [2] = 1'b0;
  assign \A[4][61] [0] = 1'b0;
  assign \A[4][62] [4] = 1'b0;
  assign \A[4][62] [3] = 1'b0;
  assign \A[4][62] [2] = 1'b0;
  assign \A[4][62] [1] = 1'b0;
  assign \A[4][63] [4] = 1'b0;
  assign \A[4][63] [3] = 1'b0;
  assign \A[4][63] [2] = 1'b0;
  assign \A[4][63] [1] = 1'b0;
  assign \A[4][63] [0] = 1'b0;
  assign \A[4][64] [4] = 1'b0;
  assign \A[4][64] [3] = 1'b0;
  assign \A[4][64] [2] = 1'b0;
  assign \A[4][64] [0] = 1'b0;
  assign \A[4][65] [4] = 1'b0;
  assign \A[4][65] [3] = 1'b0;
  assign \A[4][65] [2] = 1'b0;
  assign \A[4][65] [1] = 1'b0;
  assign \A[4][66] [0] = 1'b0;
  assign \A[4][67] [0] = 1'b0;
  assign \A[4][70] [1] = 1'b0;
  assign \A[4][70] [0] = 1'b0;
  assign \A[4][71] [4] = 1'b0;
  assign \A[4][71] [3] = 1'b0;
  assign \A[4][71] [2] = 1'b0;
  assign \A[4][71] [0] = 1'b0;
  assign \A[4][72] [4] = 1'b0;
  assign \A[4][72] [3] = 1'b0;
  assign \A[4][72] [2] = 1'b0;
  assign \A[4][72] [1] = 1'b0;
  assign \A[4][72] [0] = 1'b0;
  assign \A[4][74] [4] = 1'b0;
  assign \A[4][74] [3] = 1'b0;
  assign \A[4][74] [2] = 1'b0;
  assign \A[4][74] [0] = 1'b0;
  assign \A[4][75] [4] = 1'b0;
  assign \A[4][75] [3] = 1'b0;
  assign \A[4][75] [2] = 1'b0;
  assign \A[4][75] [1] = 1'b0;
  assign \A[4][75] [0] = 1'b0;
  assign \A[4][76] [0] = 1'b0;
  assign \A[4][77] [4] = 1'b0;
  assign \A[4][77] [3] = 1'b0;
  assign \A[4][77] [2] = 1'b0;
  assign \A[4][77] [1] = 1'b0;
  assign \A[4][78] [2] = 1'b0;
  assign \A[4][80] [0] = 1'b0;
  assign \A[4][81] [4] = 1'b0;
  assign \A[4][81] [3] = 1'b0;
  assign \A[4][81] [2] = 1'b0;
  assign \A[4][81] [0] = 1'b0;
  assign \A[4][85] [4] = 1'b0;
  assign \A[4][85] [3] = 1'b0;
  assign \A[4][85] [2] = 1'b0;
  assign \A[4][85] [0] = 1'b0;
  assign \A[4][86] [4] = 1'b0;
  assign \A[4][86] [3] = 1'b0;
  assign \A[4][86] [2] = 1'b0;
  assign \A[4][87] [4] = 1'b0;
  assign \A[4][87] [3] = 1'b0;
  assign \A[4][87] [2] = 1'b0;
  assign \A[4][87] [1] = 1'b0;
  assign \A[4][88] [4] = 1'b0;
  assign \A[4][88] [3] = 1'b0;
  assign \A[4][88] [2] = 1'b0;
  assign \A[4][88] [1] = 1'b0;
  assign \A[4][88] [0] = 1'b0;
  assign \A[4][89] [4] = 1'b0;
  assign \A[4][89] [3] = 1'b0;
  assign \A[4][89] [2] = 1'b0;
  assign \A[4][89] [1] = 1'b0;
  assign \A[4][89] [0] = 1'b0;
  assign \A[4][90] [4] = 1'b0;
  assign \A[4][90] [3] = 1'b0;
  assign \A[4][90] [2] = 1'b0;
  assign \A[4][90] [1] = 1'b0;
  assign \A[4][90] [0] = 1'b0;
  assign \A[4][91] [0] = 1'b0;
  assign \A[4][92] [4] = 1'b0;
  assign \A[4][92] [3] = 1'b0;
  assign \A[4][92] [2] = 1'b0;
  assign \A[4][92] [1] = 1'b0;
  assign \A[4][93] [4] = 1'b0;
  assign \A[4][93] [3] = 1'b0;
  assign \A[4][93] [2] = 1'b0;
  assign \A[4][93] [1] = 1'b0;
  assign \A[4][93] [0] = 1'b0;
  assign \A[4][94] [0] = 1'b0;
  assign \A[4][96] [1] = 1'b0;
  assign \A[4][97] [4] = 1'b0;
  assign \A[4][97] [3] = 1'b0;
  assign \A[4][97] [2] = 1'b0;
  assign \A[4][97] [1] = 1'b0;
  assign \A[4][98] [4] = 1'b0;
  assign \A[4][98] [3] = 1'b0;
  assign \A[4][98] [2] = 1'b0;
  assign \A[4][98] [0] = 1'b0;
  assign \A[4][99] [4] = 1'b0;
  assign \A[4][99] [3] = 1'b0;
  assign \A[4][99] [2] = 1'b0;
  assign \A[4][99] [1] = 1'b0;
  assign \A[4][99] [0] = 1'b0;
  assign \A[4][100] [4] = 1'b0;
  assign \A[4][100] [3] = 1'b0;
  assign \A[4][100] [2] = 1'b0;
  assign \A[4][100] [1] = 1'b0;
  assign \A[4][100] [0] = 1'b0;
  assign \A[4][101] [4] = 1'b0;
  assign \A[4][101] [3] = 1'b0;
  assign \A[4][101] [2] = 1'b0;
  assign \A[4][101] [0] = 1'b0;
  assign \A[4][102] [4] = 1'b0;
  assign \A[4][102] [3] = 1'b0;
  assign \A[4][102] [2] = 1'b0;
  assign \A[4][102] [1] = 1'b0;
  assign \A[4][103] [0] = 1'b0;
  assign \A[4][104] [4] = 1'b0;
  assign \A[4][104] [3] = 1'b0;
  assign \A[4][104] [2] = 1'b0;
  assign \A[4][104] [1] = 1'b0;
  assign \A[4][105] [4] = 1'b0;
  assign \A[4][105] [3] = 1'b0;
  assign \A[4][105] [2] = 1'b0;
  assign \A[4][105] [1] = 1'b0;
  assign \A[4][105] [0] = 1'b0;
  assign \A[4][106] [0] = 1'b0;
  assign \A[4][107] [4] = 1'b0;
  assign \A[4][107] [3] = 1'b0;
  assign \A[4][107] [2] = 1'b0;
  assign \A[4][107] [1] = 1'b0;
  assign \A[4][107] [0] = 1'b0;
  assign \A[4][108] [4] = 1'b0;
  assign \A[4][108] [3] = 1'b0;
  assign \A[4][108] [2] = 1'b0;
  assign \A[4][108] [1] = 1'b0;
  assign \A[4][108] [0] = 1'b0;
  assign \A[4][109] [4] = 1'b0;
  assign \A[4][109] [3] = 1'b0;
  assign \A[4][109] [2] = 1'b0;
  assign \A[4][109] [1] = 1'b0;
  assign \A[4][109] [0] = 1'b0;
  assign \A[4][110] [1] = 1'b0;
  assign \A[4][114] [4] = 1'b0;
  assign \A[4][114] [3] = 1'b0;
  assign \A[4][114] [2] = 1'b0;
  assign \A[4][114] [0] = 1'b0;
  assign \A[4][115] [4] = 1'b0;
  assign \A[4][115] [3] = 1'b0;
  assign \A[4][115] [2] = 1'b0;
  assign \A[4][115] [1] = 1'b0;
  assign \A[4][115] [0] = 1'b0;
  assign \A[4][116] [4] = 1'b0;
  assign \A[4][116] [3] = 1'b0;
  assign \A[4][116] [2] = 1'b0;
  assign \A[4][117] [4] = 1'b0;
  assign \A[4][117] [3] = 1'b0;
  assign \A[4][117] [2] = 1'b0;
  assign \A[4][117] [1] = 1'b0;
  assign \A[4][120] [4] = 1'b0;
  assign \A[4][120] [3] = 1'b0;
  assign \A[4][120] [2] = 1'b0;
  assign \A[4][120] [1] = 1'b0;
  assign \A[4][120] [0] = 1'b0;
  assign \A[4][121] [4] = 1'b0;
  assign \A[4][121] [3] = 1'b0;
  assign \A[4][121] [2] = 1'b0;
  assign \A[4][121] [1] = 1'b0;
  assign \A[4][121] [0] = 1'b0;
  assign \A[4][122] [4] = 1'b0;
  assign \A[4][122] [3] = 1'b0;
  assign \A[4][122] [2] = 1'b0;
  assign \A[4][122] [1] = 1'b0;
  assign \A[4][122] [0] = 1'b0;
  assign \A[4][123] [4] = 1'b0;
  assign \A[4][123] [3] = 1'b0;
  assign \A[4][123] [2] = 1'b0;
  assign \A[4][123] [1] = 1'b0;
  assign \A[4][123] [0] = 1'b0;
  assign \A[4][124] [0] = 1'b0;
  assign \A[4][125] [0] = 1'b0;
  assign \A[4][126] [0] = 1'b0;
  assign \A[4][127] [1] = 1'b0;
  assign \A[4][128] [4] = 1'b0;
  assign \A[4][128] [3] = 1'b0;
  assign \A[4][128] [2] = 1'b0;
  assign \A[4][128] [1] = 1'b0;
  assign \A[4][128] [0] = 1'b0;
  assign \A[4][129] [0] = 1'b0;
  assign \A[4][130] [4] = 1'b0;
  assign \A[4][130] [3] = 1'b0;
  assign \A[4][130] [2] = 1'b0;
  assign \A[4][130] [1] = 1'b0;
  assign \A[4][130] [0] = 1'b0;
  assign \A[4][131] [4] = 1'b0;
  assign \A[4][131] [3] = 1'b0;
  assign \A[4][131] [1] = 1'b0;
  assign \A[4][131] [0] = 1'b0;
  assign \A[4][132] [4] = 1'b0;
  assign \A[4][132] [3] = 1'b0;
  assign \A[4][132] [2] = 1'b0;
  assign \A[4][134] [0] = 1'b0;
  assign \A[4][135] [4] = 1'b0;
  assign \A[4][135] [3] = 1'b0;
  assign \A[4][135] [2] = 1'b0;
  assign \A[4][135] [1] = 1'b0;
  assign \A[4][135] [0] = 1'b0;
  assign \A[4][136] [0] = 1'b0;
  assign \A[4][137] [4] = 1'b0;
  assign \A[4][137] [3] = 1'b0;
  assign \A[4][137] [2] = 1'b0;
  assign \A[4][137] [0] = 1'b0;
  assign \A[4][138] [4] = 1'b0;
  assign \A[4][138] [3] = 1'b0;
  assign \A[4][138] [2] = 1'b0;
  assign \A[4][138] [1] = 1'b0;
  assign \A[4][139] [4] = 1'b0;
  assign \A[4][139] [3] = 1'b0;
  assign \A[4][139] [2] = 1'b0;
  assign \A[4][139] [1] = 1'b0;
  assign \A[4][139] [0] = 1'b0;
  assign \A[4][140] [0] = 1'b0;
  assign \A[4][141] [4] = 1'b0;
  assign \A[4][141] [3] = 1'b0;
  assign \A[4][141] [2] = 1'b0;
  assign \A[4][141] [1] = 1'b0;
  assign \A[4][141] [0] = 1'b0;
  assign \A[4][142] [4] = 1'b0;
  assign \A[4][142] [3] = 1'b0;
  assign \A[4][142] [2] = 1'b0;
  assign \A[4][142] [1] = 1'b0;
  assign \A[4][143] [4] = 1'b0;
  assign \A[4][143] [3] = 1'b0;
  assign \A[4][143] [2] = 1'b0;
  assign \A[4][143] [1] = 1'b0;
  assign \A[4][146] [4] = 1'b0;
  assign \A[4][146] [3] = 1'b0;
  assign \A[4][146] [2] = 1'b0;
  assign \A[4][146] [1] = 1'b0;
  assign \A[4][147] [4] = 1'b0;
  assign \A[4][147] [3] = 1'b0;
  assign \A[4][147] [2] = 1'b0;
  assign \A[4][147] [1] = 1'b0;
  assign \A[4][147] [0] = 1'b0;
  assign \A[4][148] [0] = 1'b0;
  assign \A[4][151] [4] = 1'b0;
  assign \A[4][151] [3] = 1'b0;
  assign \A[4][151] [2] = 1'b0;
  assign \A[4][151] [1] = 1'b0;
  assign \A[4][151] [0] = 1'b0;
  assign \A[4][152] [4] = 1'b0;
  assign \A[4][152] [3] = 1'b0;
  assign \A[4][152] [2] = 1'b0;
  assign \A[4][152] [1] = 1'b0;
  assign \A[4][152] [0] = 1'b0;
  assign \A[4][153] [4] = 1'b0;
  assign \A[4][153] [3] = 1'b0;
  assign \A[4][153] [2] = 1'b0;
  assign \A[4][153] [1] = 1'b0;
  assign \A[4][153] [0] = 1'b0;
  assign \A[4][154] [4] = 1'b0;
  assign \A[4][154] [3] = 1'b0;
  assign \A[4][154] [2] = 1'b0;
  assign \A[4][154] [1] = 1'b0;
  assign \A[4][155] [0] = 1'b0;
  assign \A[4][156] [4] = 1'b0;
  assign \A[4][156] [3] = 1'b0;
  assign \A[4][156] [2] = 1'b0;
  assign \A[4][156] [1] = 1'b0;
  assign \A[4][156] [0] = 1'b0;
  assign \A[4][158] [0] = 1'b0;
  assign \A[4][159] [4] = 1'b0;
  assign \A[4][159] [3] = 1'b0;
  assign \A[4][159] [2] = 1'b0;
  assign \A[4][159] [1] = 1'b0;
  assign \A[4][160] [4] = 1'b0;
  assign \A[4][160] [3] = 1'b0;
  assign \A[4][160] [2] = 1'b0;
  assign \A[4][160] [0] = 1'b0;
  assign \A[4][161] [4] = 1'b0;
  assign \A[4][161] [3] = 1'b0;
  assign \A[4][161] [2] = 1'b0;
  assign \A[4][161] [1] = 1'b0;
  assign \A[4][162] [4] = 1'b0;
  assign \A[4][162] [3] = 1'b0;
  assign \A[4][162] [2] = 1'b0;
  assign \A[4][162] [0] = 1'b0;
  assign \A[4][163] [4] = 1'b0;
  assign \A[4][163] [3] = 1'b0;
  assign \A[4][163] [2] = 1'b0;
  assign \A[4][163] [0] = 1'b0;
  assign \A[4][164] [0] = 1'b0;
  assign \A[4][165] [4] = 1'b0;
  assign \A[4][165] [3] = 1'b0;
  assign \A[4][165] [2] = 1'b0;
  assign \A[4][165] [1] = 1'b0;
  assign \A[4][165] [0] = 1'b0;
  assign \A[4][167] [0] = 1'b0;
  assign \A[4][169] [0] = 1'b0;
  assign \A[4][170] [4] = 1'b0;
  assign \A[4][170] [3] = 1'b0;
  assign \A[4][170] [2] = 1'b0;
  assign \A[4][170] [1] = 1'b0;
  assign \A[4][170] [0] = 1'b0;
  assign \A[4][171] [4] = 1'b0;
  assign \A[4][171] [3] = 1'b0;
  assign \A[4][171] [2] = 1'b0;
  assign \A[4][171] [1] = 1'b0;
  assign \A[4][173] [4] = 1'b0;
  assign \A[4][173] [3] = 1'b0;
  assign \A[4][173] [2] = 1'b0;
  assign \A[4][173] [0] = 1'b0;
  assign \A[4][175] [4] = 1'b0;
  assign \A[4][175] [3] = 1'b0;
  assign \A[4][175] [2] = 1'b0;
  assign \A[4][175] [1] = 1'b0;
  assign \A[4][176] [4] = 1'b0;
  assign \A[4][176] [3] = 1'b0;
  assign \A[4][176] [2] = 1'b0;
  assign \A[4][176] [1] = 1'b0;
  assign \A[4][177] [4] = 1'b0;
  assign \A[4][177] [3] = 1'b0;
  assign \A[4][177] [2] = 1'b0;
  assign \A[4][179] [4] = 1'b0;
  assign \A[4][179] [3] = 1'b0;
  assign \A[4][179] [2] = 1'b0;
  assign \A[4][179] [1] = 1'b0;
  assign \A[4][181] [4] = 1'b0;
  assign \A[4][181] [3] = 1'b0;
  assign \A[4][181] [2] = 1'b0;
  assign \A[4][181] [1] = 1'b0;
  assign \A[4][181] [0] = 1'b0;
  assign \A[4][182] [1] = 1'b0;
  assign \A[4][184] [4] = 1'b0;
  assign \A[4][184] [3] = 1'b0;
  assign \A[4][184] [2] = 1'b0;
  assign \A[4][184] [1] = 1'b0;
  assign \A[4][184] [0] = 1'b0;
  assign \A[4][185] [4] = 1'b0;
  assign \A[4][185] [3] = 1'b0;
  assign \A[4][185] [2] = 1'b0;
  assign \A[4][185] [1] = 1'b0;
  assign \A[4][185] [0] = 1'b0;
  assign \A[4][186] [4] = 1'b0;
  assign \A[4][186] [3] = 1'b0;
  assign \A[4][186] [2] = 1'b0;
  assign \A[4][186] [1] = 1'b0;
  assign \A[4][187] [4] = 1'b0;
  assign \A[4][187] [3] = 1'b0;
  assign \A[4][187] [2] = 1'b0;
  assign \A[4][187] [1] = 1'b0;
  assign \A[4][188] [4] = 1'b0;
  assign \A[4][188] [3] = 1'b0;
  assign \A[4][188] [2] = 1'b0;
  assign \A[4][189] [4] = 1'b0;
  assign \A[4][189] [3] = 1'b0;
  assign \A[4][189] [2] = 1'b0;
  assign \A[4][189] [1] = 1'b0;
  assign \A[4][189] [0] = 1'b0;
  assign \A[4][190] [4] = 1'b0;
  assign \A[4][190] [3] = 1'b0;
  assign \A[4][190] [2] = 1'b0;
  assign \A[4][190] [0] = 1'b0;
  assign \A[4][191] [4] = 1'b0;
  assign \A[4][191] [3] = 1'b0;
  assign \A[4][191] [2] = 1'b0;
  assign \A[4][191] [1] = 1'b0;
  assign \A[4][192] [0] = 1'b0;
  assign \A[4][193] [4] = 1'b0;
  assign \A[4][193] [3] = 1'b0;
  assign \A[4][193] [2] = 1'b0;
  assign \A[4][193] [1] = 1'b0;
  assign \A[4][193] [0] = 1'b0;
  assign \A[4][194] [4] = 1'b0;
  assign \A[4][194] [3] = 1'b0;
  assign \A[4][194] [2] = 1'b0;
  assign \A[4][194] [1] = 1'b0;
  assign \A[4][195] [4] = 1'b0;
  assign \A[4][195] [3] = 1'b0;
  assign \A[4][195] [2] = 1'b0;
  assign \A[4][195] [1] = 1'b0;
  assign \A[4][196] [0] = 1'b0;
  assign \A[4][197] [1] = 1'b0;
  assign \A[4][198] [4] = 1'b0;
  assign \A[4][198] [3] = 1'b0;
  assign \A[4][198] [2] = 1'b0;
  assign \A[4][198] [1] = 1'b0;
  assign \A[4][198] [0] = 1'b0;
  assign \A[4][199] [4] = 1'b0;
  assign \A[4][199] [3] = 1'b0;
  assign \A[4][199] [2] = 1'b0;
  assign \A[4][199] [0] = 1'b0;
  assign \A[4][200] [4] = 1'b0;
  assign \A[4][200] [3] = 1'b0;
  assign \A[4][200] [2] = 1'b0;
  assign \A[4][200] [1] = 1'b0;
  assign \A[4][200] [0] = 1'b0;
  assign \A[4][201] [4] = 1'b0;
  assign \A[4][201] [3] = 1'b0;
  assign \A[4][201] [2] = 1'b0;
  assign \A[4][201] [1] = 1'b0;
  assign \A[4][201] [0] = 1'b0;
  assign \A[4][203] [4] = 1'b0;
  assign \A[4][203] [3] = 1'b0;
  assign \A[4][203] [2] = 1'b0;
  assign \A[4][203] [1] = 1'b0;
  assign \A[4][203] [0] = 1'b0;
  assign \A[4][205] [4] = 1'b0;
  assign \A[4][205] [3] = 1'b0;
  assign \A[4][205] [2] = 1'b0;
  assign \A[4][206] [4] = 1'b0;
  assign \A[4][206] [3] = 1'b0;
  assign \A[4][206] [2] = 1'b0;
  assign \A[4][206] [1] = 1'b0;
  assign \A[4][206] [0] = 1'b0;
  assign \A[4][207] [4] = 1'b0;
  assign \A[4][207] [3] = 1'b0;
  assign \A[4][207] [2] = 1'b0;
  assign \A[4][207] [0] = 1'b0;
  assign \A[4][208] [4] = 1'b0;
  assign \A[4][208] [3] = 1'b0;
  assign \A[4][208] [2] = 1'b0;
  assign \A[4][208] [1] = 1'b0;
  assign \A[4][209] [1] = 1'b0;
  assign \A[4][211] [4] = 1'b0;
  assign \A[4][211] [3] = 1'b0;
  assign \A[4][211] [2] = 1'b0;
  assign \A[4][211] [1] = 1'b0;
  assign \A[4][213] [4] = 1'b0;
  assign \A[4][213] [3] = 1'b0;
  assign \A[4][213] [2] = 1'b0;
  assign \A[4][213] [1] = 1'b0;
  assign \A[4][213] [0] = 1'b0;
  assign \A[4][216] [4] = 1'b0;
  assign \A[4][216] [3] = 1'b0;
  assign \A[4][216] [2] = 1'b0;
  assign \A[4][216] [1] = 1'b0;
  assign \A[4][216] [0] = 1'b0;
  assign \A[4][217] [4] = 1'b0;
  assign \A[4][217] [3] = 1'b0;
  assign \A[4][217] [2] = 1'b0;
  assign \A[4][219] [4] = 1'b0;
  assign \A[4][219] [3] = 1'b0;
  assign \A[4][219] [2] = 1'b0;
  assign \A[4][219] [0] = 1'b0;
  assign \A[4][220] [4] = 1'b0;
  assign \A[4][220] [3] = 1'b0;
  assign \A[4][220] [2] = 1'b0;
  assign \A[4][220] [0] = 1'b0;
  assign \A[4][222] [4] = 1'b0;
  assign \A[4][222] [3] = 1'b0;
  assign \A[4][222] [2] = 1'b0;
  assign \A[4][222] [1] = 1'b0;
  assign \A[4][222] [0] = 1'b0;
  assign \A[4][223] [4] = 1'b0;
  assign \A[4][223] [3] = 1'b0;
  assign \A[4][223] [2] = 1'b0;
  assign \A[4][223] [0] = 1'b0;
  assign \A[4][226] [4] = 1'b0;
  assign \A[4][226] [3] = 1'b0;
  assign \A[4][226] [2] = 1'b0;
  assign \A[4][226] [1] = 1'b0;
  assign \A[4][227] [4] = 1'b0;
  assign \A[4][227] [3] = 1'b0;
  assign \A[4][227] [2] = 1'b0;
  assign \A[4][227] [1] = 1'b0;
  assign \A[4][227] [0] = 1'b0;
  assign \A[4][228] [4] = 1'b0;
  assign \A[4][228] [3] = 1'b0;
  assign \A[4][228] [2] = 1'b0;
  assign \A[4][228] [0] = 1'b0;
  assign \A[4][231] [4] = 1'b0;
  assign \A[4][231] [3] = 1'b0;
  assign \A[4][231] [2] = 1'b0;
  assign \A[4][231] [1] = 1'b0;
  assign \A[4][231] [0] = 1'b0;
  assign \A[4][233] [0] = 1'b0;
  assign \A[4][235] [4] = 1'b0;
  assign \A[4][235] [3] = 1'b0;
  assign \A[4][235] [2] = 1'b0;
  assign \A[4][235] [1] = 1'b0;
  assign \A[4][236] [4] = 1'b0;
  assign \A[4][236] [3] = 1'b0;
  assign \A[4][236] [2] = 1'b0;
  assign \A[4][236] [1] = 1'b0;
  assign \A[4][236] [0] = 1'b0;
  assign \A[4][237] [4] = 1'b0;
  assign \A[4][237] [3] = 1'b0;
  assign \A[4][237] [2] = 1'b0;
  assign \A[4][237] [1] = 1'b0;
  assign \A[4][238] [0] = 1'b0;
  assign \A[4][239] [4] = 1'b0;
  assign \A[4][239] [3] = 1'b0;
  assign \A[4][239] [2] = 1'b0;
  assign \A[4][239] [0] = 1'b0;
  assign \A[4][240] [4] = 1'b0;
  assign \A[4][240] [3] = 1'b0;
  assign \A[4][240] [2] = 1'b0;
  assign \A[4][241] [4] = 1'b0;
  assign \A[4][241] [3] = 1'b0;
  assign \A[4][241] [2] = 1'b0;
  assign \A[4][241] [1] = 1'b0;
  assign \A[4][241] [0] = 1'b0;
  assign \A[4][242] [4] = 1'b0;
  assign \A[4][242] [3] = 1'b0;
  assign \A[4][242] [2] = 1'b0;
  assign \A[4][242] [1] = 1'b0;
  assign \A[4][245] [4] = 1'b0;
  assign \A[4][245] [3] = 1'b0;
  assign \A[4][245] [2] = 1'b0;
  assign \A[4][245] [1] = 1'b0;
  assign \A[4][246] [4] = 1'b0;
  assign \A[4][246] [3] = 1'b0;
  assign \A[4][246] [2] = 1'b0;
  assign \A[4][246] [1] = 1'b0;
  assign \A[4][247] [4] = 1'b0;
  assign \A[4][247] [3] = 1'b0;
  assign \A[4][247] [2] = 1'b0;
  assign \A[4][250] [4] = 1'b0;
  assign \A[4][250] [3] = 1'b0;
  assign \A[4][250] [2] = 1'b0;
  assign \A[4][250] [1] = 1'b0;
  assign \A[4][250] [0] = 1'b0;
  assign \A[4][251] [4] = 1'b0;
  assign \A[4][251] [3] = 1'b0;
  assign \A[4][251] [2] = 1'b0;
  assign \A[4][251] [1] = 1'b0;
  assign \A[4][252] [4] = 1'b0;
  assign \A[4][252] [3] = 1'b0;
  assign \A[4][252] [2] = 1'b0;
  assign \A[4][252] [1] = 1'b0;
  assign \A[4][253] [4] = 1'b0;
  assign \A[4][253] [3] = 1'b0;
  assign \A[4][253] [2] = 1'b0;
  assign \A[4][253] [1] = 1'b0;
  assign \A[4][255] [4] = 1'b0;
  assign \A[4][255] [3] = 1'b0;
  assign \A[4][255] [2] = 1'b0;
  assign \A[4][255] [1] = 1'b0;
  assign \A[5][0] [0] = 1'b0;
  assign \A[5][1] [4] = 1'b0;
  assign \A[5][1] [3] = 1'b0;
  assign \A[5][1] [2] = 1'b0;
  assign \A[5][1] [1] = 1'b0;
  assign \A[5][1] [0] = 1'b0;
  assign \A[5][4] [4] = 1'b0;
  assign \A[5][4] [3] = 1'b0;
  assign \A[5][4] [2] = 1'b0;
  assign \A[5][4] [1] = 1'b0;
  assign \A[5][4] [0] = 1'b0;
  assign \A[5][9] [4] = 1'b0;
  assign \A[5][9] [3] = 1'b0;
  assign \A[5][9] [2] = 1'b0;
  assign \A[5][9] [1] = 1'b0;
  assign \A[5][9] [0] = 1'b0;
  assign \A[5][12] [1] = 1'b0;
  assign \A[5][13] [1] = 1'b0;
  assign \A[5][15] [0] = 1'b0;
  assign \A[5][17] [4] = 1'b0;
  assign \A[5][17] [3] = 1'b0;
  assign \A[5][17] [2] = 1'b0;
  assign \A[5][17] [1] = 1'b0;
  assign \A[5][19] [4] = 1'b0;
  assign \A[5][19] [3] = 1'b0;
  assign \A[5][19] [2] = 1'b0;
  assign \A[5][19] [0] = 1'b0;
  assign \A[5][20] [4] = 1'b0;
  assign \A[5][20] [3] = 1'b0;
  assign \A[5][20] [2] = 1'b0;
  assign \A[5][20] [1] = 1'b0;
  assign \A[5][21] [4] = 1'b0;
  assign \A[5][21] [3] = 1'b0;
  assign \A[5][21] [2] = 1'b0;
  assign \A[5][21] [1] = 1'b0;
  assign \A[5][21] [0] = 1'b0;
  assign \A[5][22] [4] = 1'b0;
  assign \A[5][22] [3] = 1'b0;
  assign \A[5][22] [2] = 1'b0;
  assign \A[5][22] [0] = 1'b0;
  assign \A[5][24] [0] = 1'b0;
  assign \A[5][27] [4] = 1'b0;
  assign \A[5][27] [3] = 1'b0;
  assign \A[5][27] [2] = 1'b0;
  assign \A[5][27] [1] = 1'b0;
  assign \A[5][27] [0] = 1'b0;
  assign \A[5][28] [4] = 1'b0;
  assign \A[5][28] [3] = 1'b0;
  assign \A[5][28] [2] = 1'b0;
  assign \A[5][28] [1] = 1'b0;
  assign \A[5][28] [0] = 1'b0;
  assign \A[5][32] [4] = 1'b0;
  assign \A[5][32] [3] = 1'b0;
  assign \A[5][32] [2] = 1'b0;
  assign \A[5][32] [1] = 1'b0;
  assign \A[5][32] [0] = 1'b0;
  assign \A[5][33] [4] = 1'b0;
  assign \A[5][33] [3] = 1'b0;
  assign \A[5][33] [2] = 1'b0;
  assign \A[5][33] [1] = 1'b0;
  assign \A[5][33] [0] = 1'b0;
  assign \A[5][35] [4] = 1'b0;
  assign \A[5][35] [3] = 1'b0;
  assign \A[5][35] [2] = 1'b0;
  assign \A[5][35] [1] = 1'b0;
  assign \A[5][36] [4] = 1'b0;
  assign \A[5][36] [3] = 1'b0;
  assign \A[5][36] [2] = 1'b0;
  assign \A[5][36] [1] = 1'b0;
  assign \A[5][36] [0] = 1'b0;
  assign \A[5][37] [4] = 1'b0;
  assign \A[5][37] [3] = 1'b0;
  assign \A[5][37] [2] = 1'b0;
  assign \A[5][37] [1] = 1'b0;
  assign \A[5][38] [4] = 1'b0;
  assign \A[5][38] [3] = 1'b0;
  assign \A[5][38] [2] = 1'b0;
  assign \A[5][38] [0] = 1'b0;
  assign \A[5][39] [4] = 1'b0;
  assign \A[5][39] [3] = 1'b0;
  assign \A[5][39] [2] = 1'b0;
  assign \A[5][41] [0] = 1'b0;
  assign \A[5][42] [2] = 1'b0;
  assign \A[5][43] [0] = 1'b0;
  assign \A[5][44] [1] = 1'b0;
  assign \A[5][45] [0] = 1'b0;
  assign \A[5][46] [4] = 1'b0;
  assign \A[5][46] [3] = 1'b0;
  assign \A[5][46] [2] = 1'b0;
  assign \A[5][46] [1] = 1'b0;
  assign \A[5][46] [0] = 1'b0;
  assign \A[5][47] [4] = 1'b0;
  assign \A[5][47] [3] = 1'b0;
  assign \A[5][47] [2] = 1'b0;
  assign \A[5][47] [1] = 1'b0;
  assign \A[5][47] [0] = 1'b0;
  assign \A[5][48] [4] = 1'b0;
  assign \A[5][48] [3] = 1'b0;
  assign \A[5][48] [2] = 1'b0;
  assign \A[5][48] [1] = 1'b0;
  assign \A[5][48] [0] = 1'b0;
  assign \A[5][51] [4] = 1'b0;
  assign \A[5][51] [3] = 1'b0;
  assign \A[5][51] [2] = 1'b0;
  assign \A[5][51] [0] = 1'b0;
  assign \A[5][53] [4] = 1'b0;
  assign \A[5][53] [3] = 1'b0;
  assign \A[5][53] [2] = 1'b0;
  assign \A[5][53] [1] = 1'b0;
  assign \A[5][54] [4] = 1'b0;
  assign \A[5][54] [3] = 1'b0;
  assign \A[5][54] [2] = 1'b0;
  assign \A[5][54] [0] = 1'b0;
  assign \A[5][55] [4] = 1'b0;
  assign \A[5][55] [3] = 1'b0;
  assign \A[5][55] [2] = 1'b0;
  assign \A[5][55] [1] = 1'b0;
  assign \A[5][55] [0] = 1'b0;
  assign \A[5][56] [4] = 1'b0;
  assign \A[5][56] [3] = 1'b0;
  assign \A[5][56] [2] = 1'b0;
  assign \A[5][56] [1] = 1'b0;
  assign \A[5][56] [0] = 1'b0;
  assign \A[5][57] [4] = 1'b0;
  assign \A[5][57] [3] = 1'b0;
  assign \A[5][57] [2] = 1'b0;
  assign \A[5][57] [1] = 1'b0;
  assign \A[5][57] [0] = 1'b0;
  assign \A[5][60] [0] = 1'b0;
  assign \A[5][61] [4] = 1'b0;
  assign \A[5][61] [3] = 1'b0;
  assign \A[5][61] [2] = 1'b0;
  assign \A[5][61] [1] = 1'b0;
  assign \A[5][61] [0] = 1'b0;
  assign \A[5][62] [4] = 1'b0;
  assign \A[5][62] [3] = 1'b0;
  assign \A[5][62] [2] = 1'b0;
  assign \A[5][62] [1] = 1'b0;
  assign \A[5][63] [4] = 1'b0;
  assign \A[5][63] [3] = 1'b0;
  assign \A[5][63] [2] = 1'b0;
  assign \A[5][63] [0] = 1'b0;
  assign \A[5][64] [4] = 1'b0;
  assign \A[5][64] [3] = 1'b0;
  assign \A[5][64] [2] = 1'b0;
  assign \A[5][64] [0] = 1'b0;
  assign \A[5][66] [4] = 1'b0;
  assign \A[5][66] [3] = 1'b0;
  assign \A[5][66] [2] = 1'b0;
  assign \A[5][66] [1] = 1'b0;
  assign \A[5][66] [0] = 1'b0;
  assign \A[5][67] [4] = 1'b0;
  assign \A[5][67] [3] = 1'b0;
  assign \A[5][67] [2] = 1'b0;
  assign \A[5][67] [1] = 1'b0;
  assign \A[5][68] [4] = 1'b0;
  assign \A[5][68] [3] = 1'b0;
  assign \A[5][68] [2] = 1'b0;
  assign \A[5][68] [1] = 1'b0;
  assign \A[5][69] [4] = 1'b0;
  assign \A[5][69] [3] = 1'b0;
  assign \A[5][69] [2] = 1'b0;
  assign \A[5][69] [1] = 1'b0;
  assign \A[5][70] [4] = 1'b0;
  assign \A[5][70] [3] = 1'b0;
  assign \A[5][70] [2] = 1'b0;
  assign \A[5][71] [0] = 1'b0;
  assign \A[5][73] [0] = 1'b0;
  assign \A[5][74] [4] = 1'b0;
  assign \A[5][74] [3] = 1'b0;
  assign \A[5][74] [2] = 1'b0;
  assign \A[5][77] [4] = 1'b0;
  assign \A[5][77] [3] = 1'b0;
  assign \A[5][77] [2] = 1'b0;
  assign \A[5][77] [1] = 1'b0;
  assign \A[5][77] [0] = 1'b0;
  assign \A[5][79] [4] = 1'b0;
  assign \A[5][79] [3] = 1'b0;
  assign \A[5][79] [2] = 1'b0;
  assign \A[5][79] [1] = 1'b0;
  assign \A[5][79] [0] = 1'b0;
  assign \A[5][80] [4] = 1'b0;
  assign \A[5][80] [3] = 1'b0;
  assign \A[5][80] [2] = 1'b0;
  assign \A[5][80] [1] = 1'b0;
  assign \A[5][80] [0] = 1'b0;
  assign \A[5][81] [4] = 1'b0;
  assign \A[5][81] [3] = 1'b0;
  assign \A[5][81] [2] = 1'b0;
  assign \A[5][81] [1] = 1'b0;
  assign \A[5][81] [0] = 1'b0;
  assign \A[5][82] [0] = 1'b0;
  assign \A[5][84] [4] = 1'b0;
  assign \A[5][84] [3] = 1'b0;
  assign \A[5][84] [2] = 1'b0;
  assign \A[5][84] [0] = 1'b0;
  assign \A[5][85] [4] = 1'b0;
  assign \A[5][85] [3] = 1'b0;
  assign \A[5][85] [2] = 1'b0;
  assign \A[5][85] [1] = 1'b0;
  assign \A[5][86] [4] = 1'b0;
  assign \A[5][86] [3] = 1'b0;
  assign \A[5][86] [2] = 1'b0;
  assign \A[5][86] [1] = 1'b0;
  assign \A[5][87] [4] = 1'b0;
  assign \A[5][87] [3] = 1'b0;
  assign \A[5][87] [2] = 1'b0;
  assign \A[5][87] [1] = 1'b0;
  assign \A[5][88] [4] = 1'b0;
  assign \A[5][88] [3] = 1'b0;
  assign \A[5][88] [2] = 1'b0;
  assign \A[5][88] [1] = 1'b0;
  assign \A[5][89] [0] = 1'b0;
  assign \A[5][90] [0] = 1'b0;
  assign \A[5][91] [0] = 1'b0;
  assign \A[5][92] [4] = 1'b0;
  assign \A[5][92] [3] = 1'b0;
  assign \A[5][92] [2] = 1'b0;
  assign \A[5][92] [1] = 1'b0;
  assign \A[5][93] [4] = 1'b0;
  assign \A[5][93] [3] = 1'b0;
  assign \A[5][93] [2] = 1'b0;
  assign \A[5][93] [1] = 1'b0;
  assign \A[5][93] [0] = 1'b0;
  assign \A[5][94] [4] = 1'b0;
  assign \A[5][94] [3] = 1'b0;
  assign \A[5][94] [2] = 1'b0;
  assign \A[5][94] [1] = 1'b0;
  assign \A[5][94] [0] = 1'b0;
  assign \A[5][96] [4] = 1'b0;
  assign \A[5][96] [3] = 1'b0;
  assign \A[5][96] [2] = 1'b0;
  assign \A[5][96] [1] = 1'b0;
  assign \A[5][97] [4] = 1'b0;
  assign \A[5][97] [3] = 1'b0;
  assign \A[5][97] [2] = 1'b0;
  assign \A[5][97] [1] = 1'b0;
  assign \A[5][97] [0] = 1'b0;
  assign \A[5][99] [4] = 1'b0;
  assign \A[5][99] [3] = 1'b0;
  assign \A[5][99] [2] = 1'b0;
  assign \A[5][100] [4] = 1'b0;
  assign \A[5][100] [3] = 1'b0;
  assign \A[5][100] [2] = 1'b0;
  assign \A[5][100] [1] = 1'b0;
  assign \A[5][102] [4] = 1'b0;
  assign \A[5][102] [3] = 1'b0;
  assign \A[5][102] [2] = 1'b0;
  assign \A[5][102] [1] = 1'b0;
  assign \A[5][103] [4] = 1'b0;
  assign \A[5][103] [3] = 1'b0;
  assign \A[5][103] [2] = 1'b0;
  assign \A[5][103] [0] = 1'b0;
  assign \A[5][104] [4] = 1'b0;
  assign \A[5][104] [3] = 1'b0;
  assign \A[5][104] [2] = 1'b0;
  assign \A[5][104] [1] = 1'b0;
  assign \A[5][104] [0] = 1'b0;
  assign \A[5][105] [4] = 1'b0;
  assign \A[5][105] [3] = 1'b0;
  assign \A[5][105] [2] = 1'b0;
  assign \A[5][105] [1] = 1'b0;
  assign \A[5][105] [0] = 1'b0;
  assign \A[5][106] [4] = 1'b0;
  assign \A[5][106] [3] = 1'b0;
  assign \A[5][106] [2] = 1'b0;
  assign \A[5][106] [1] = 1'b0;
  assign \A[5][106] [0] = 1'b0;
  assign \A[5][107] [0] = 1'b0;
  assign \A[5][108] [1] = 1'b0;
  assign \A[5][109] [4] = 1'b0;
  assign \A[5][109] [3] = 1'b0;
  assign \A[5][109] [2] = 1'b0;
  assign \A[5][109] [1] = 1'b0;
  assign \A[5][109] [0] = 1'b0;
  assign \A[5][110] [4] = 1'b0;
  assign \A[5][110] [3] = 1'b0;
  assign \A[5][110] [2] = 1'b0;
  assign \A[5][111] [4] = 1'b0;
  assign \A[5][111] [3] = 1'b0;
  assign \A[5][111] [2] = 1'b0;
  assign \A[5][111] [1] = 1'b0;
  assign \A[5][112] [4] = 1'b0;
  assign \A[5][112] [3] = 1'b0;
  assign \A[5][112] [2] = 1'b0;
  assign \A[5][112] [1] = 1'b0;
  assign \A[5][112] [0] = 1'b0;
  assign \A[5][114] [4] = 1'b0;
  assign \A[5][114] [3] = 1'b0;
  assign \A[5][114] [2] = 1'b0;
  assign \A[5][114] [0] = 1'b0;
  assign \A[5][115] [4] = 1'b0;
  assign \A[5][115] [3] = 1'b0;
  assign \A[5][115] [2] = 1'b0;
  assign \A[5][115] [1] = 1'b0;
  assign \A[5][115] [0] = 1'b0;
  assign \A[5][116] [4] = 1'b0;
  assign \A[5][116] [3] = 1'b0;
  assign \A[5][116] [2] = 1'b0;
  assign \A[5][116] [1] = 1'b0;
  assign \A[5][116] [0] = 1'b0;
  assign \A[5][117] [4] = 1'b0;
  assign \A[5][117] [3] = 1'b0;
  assign \A[5][117] [2] = 1'b0;
  assign \A[5][117] [1] = 1'b0;
  assign \A[5][117] [0] = 1'b0;
  assign \A[5][118] [4] = 1'b0;
  assign \A[5][118] [3] = 1'b0;
  assign \A[5][118] [2] = 1'b0;
  assign \A[5][119] [4] = 1'b0;
  assign \A[5][119] [3] = 1'b0;
  assign \A[5][119] [2] = 1'b0;
  assign \A[5][119] [1] = 1'b0;
  assign \A[5][119] [0] = 1'b0;
  assign \A[5][121] [1] = 1'b0;
  assign \A[5][122] [4] = 1'b0;
  assign \A[5][122] [3] = 1'b0;
  assign \A[5][122] [2] = 1'b0;
  assign \A[5][122] [1] = 1'b0;
  assign \A[5][122] [0] = 1'b0;
  assign \A[5][123] [4] = 1'b0;
  assign \A[5][123] [3] = 1'b0;
  assign \A[5][123] [2] = 1'b0;
  assign \A[5][123] [1] = 1'b0;
  assign \A[5][123] [0] = 1'b0;
  assign \A[5][124] [0] = 1'b0;
  assign \A[5][128] [4] = 1'b0;
  assign \A[5][128] [3] = 1'b0;
  assign \A[5][128] [2] = 1'b0;
  assign \A[5][128] [1] = 1'b0;
  assign \A[5][130] [4] = 1'b0;
  assign \A[5][130] [3] = 1'b0;
  assign \A[5][130] [2] = 1'b0;
  assign \A[5][130] [0] = 1'b0;
  assign \A[5][131] [4] = 1'b0;
  assign \A[5][131] [3] = 1'b0;
  assign \A[5][131] [2] = 1'b0;
  assign \A[5][131] [1] = 1'b0;
  assign \A[5][131] [0] = 1'b0;
  assign \A[5][132] [4] = 1'b0;
  assign \A[5][132] [3] = 1'b0;
  assign \A[5][132] [2] = 1'b0;
  assign \A[5][132] [1] = 1'b0;
  assign \A[5][134] [4] = 1'b0;
  assign \A[5][134] [3] = 1'b0;
  assign \A[5][134] [2] = 1'b0;
  assign \A[5][134] [1] = 1'b0;
  assign \A[5][135] [4] = 1'b0;
  assign \A[5][135] [3] = 1'b0;
  assign \A[5][135] [2] = 1'b0;
  assign \A[5][135] [1] = 1'b0;
  assign \A[5][135] [0] = 1'b0;
  assign \A[5][136] [4] = 1'b0;
  assign \A[5][136] [3] = 1'b0;
  assign \A[5][136] [2] = 1'b0;
  assign \A[5][136] [1] = 1'b0;
  assign \A[5][136] [0] = 1'b0;
  assign \A[5][137] [0] = 1'b0;
  assign \A[5][138] [4] = 1'b0;
  assign \A[5][138] [3] = 1'b0;
  assign \A[5][138] [2] = 1'b0;
  assign \A[5][138] [1] = 1'b0;
  assign \A[5][138] [0] = 1'b0;
  assign \A[5][139] [0] = 1'b0;
  assign \A[5][140] [1] = 1'b0;
  assign \A[5][141] [0] = 1'b0;
  assign \A[5][142] [0] = 1'b0;
  assign \A[5][143] [4] = 1'b0;
  assign \A[5][143] [3] = 1'b0;
  assign \A[5][143] [2] = 1'b0;
  assign \A[5][143] [1] = 1'b0;
  assign \A[5][144] [1] = 1'b0;
  assign \A[5][144] [0] = 1'b0;
  assign \A[5][145] [4] = 1'b0;
  assign \A[5][145] [3] = 1'b0;
  assign \A[5][145] [2] = 1'b0;
  assign \A[5][145] [1] = 1'b0;
  assign \A[5][145] [0] = 1'b0;
  assign \A[5][146] [1] = 1'b0;
  assign \A[5][148] [4] = 1'b0;
  assign \A[5][148] [3] = 1'b0;
  assign \A[5][148] [2] = 1'b0;
  assign \A[5][148] [1] = 1'b0;
  assign \A[5][148] [0] = 1'b0;
  assign \A[5][149] [4] = 1'b0;
  assign \A[5][149] [3] = 1'b0;
  assign \A[5][149] [2] = 1'b0;
  assign \A[5][149] [0] = 1'b0;
  assign \A[5][150] [4] = 1'b0;
  assign \A[5][150] [3] = 1'b0;
  assign \A[5][150] [2] = 1'b0;
  assign \A[5][150] [1] = 1'b0;
  assign \A[5][150] [0] = 1'b0;
  assign \A[5][151] [4] = 1'b0;
  assign \A[5][151] [3] = 1'b0;
  assign \A[5][151] [2] = 1'b0;
  assign \A[5][151] [1] = 1'b0;
  assign \A[5][152] [1] = 1'b0;
  assign \A[5][153] [4] = 1'b0;
  assign \A[5][153] [3] = 1'b0;
  assign \A[5][153] [2] = 1'b0;
  assign \A[5][153] [1] = 1'b0;
  assign \A[5][154] [1] = 1'b0;
  assign \A[5][155] [0] = 1'b0;
  assign \A[5][158] [4] = 1'b0;
  assign \A[5][158] [3] = 1'b0;
  assign \A[5][158] [2] = 1'b0;
  assign \A[5][158] [1] = 1'b0;
  assign \A[5][158] [0] = 1'b0;
  assign \A[5][160] [0] = 1'b0;
  assign \A[5][162] [0] = 1'b0;
  assign \A[5][164] [4] = 1'b0;
  assign \A[5][164] [3] = 1'b0;
  assign \A[5][164] [2] = 1'b0;
  assign \A[5][164] [1] = 1'b0;
  assign \A[5][164] [0] = 1'b0;
  assign \A[5][165] [4] = 1'b0;
  assign \A[5][165] [3] = 1'b0;
  assign \A[5][165] [2] = 1'b0;
  assign \A[5][165] [1] = 1'b0;
  assign \A[5][166] [4] = 1'b0;
  assign \A[5][166] [3] = 1'b0;
  assign \A[5][166] [2] = 1'b0;
  assign \A[5][166] [0] = 1'b0;
  assign \A[5][167] [0] = 1'b0;
  assign \A[5][168] [4] = 1'b0;
  assign \A[5][168] [3] = 1'b0;
  assign \A[5][168] [2] = 1'b0;
  assign \A[5][168] [1] = 1'b0;
  assign \A[5][168] [0] = 1'b0;
  assign \A[5][169] [4] = 1'b0;
  assign \A[5][169] [3] = 1'b0;
  assign \A[5][169] [2] = 1'b0;
  assign \A[5][172] [4] = 1'b0;
  assign \A[5][172] [3] = 1'b0;
  assign \A[5][172] [2] = 1'b0;
  assign \A[5][172] [1] = 1'b0;
  assign \A[5][172] [0] = 1'b0;
  assign \A[5][173] [4] = 1'b0;
  assign \A[5][173] [3] = 1'b0;
  assign \A[5][173] [2] = 1'b0;
  assign \A[5][173] [1] = 1'b0;
  assign \A[5][175] [1] = 1'b0;
  assign \A[5][177] [0] = 1'b0;
  assign \A[5][178] [4] = 1'b0;
  assign \A[5][178] [3] = 1'b0;
  assign \A[5][178] [2] = 1'b0;
  assign \A[5][178] [1] = 1'b0;
  assign \A[5][179] [4] = 1'b0;
  assign \A[5][179] [3] = 1'b0;
  assign \A[5][179] [2] = 1'b0;
  assign \A[5][179] [1] = 1'b0;
  assign \A[5][180] [0] = 1'b0;
  assign \A[5][181] [4] = 1'b0;
  assign \A[5][181] [3] = 1'b0;
  assign \A[5][181] [2] = 1'b0;
  assign \A[5][181] [0] = 1'b0;
  assign \A[5][182] [4] = 1'b0;
  assign \A[5][182] [3] = 1'b0;
  assign \A[5][182] [2] = 1'b0;
  assign \A[5][182] [0] = 1'b0;
  assign \A[5][183] [4] = 1'b0;
  assign \A[5][183] [3] = 1'b0;
  assign \A[5][183] [2] = 1'b0;
  assign \A[5][183] [1] = 1'b0;
  assign \A[5][185] [4] = 1'b0;
  assign \A[5][185] [3] = 1'b0;
  assign \A[5][185] [2] = 1'b0;
  assign \A[5][185] [1] = 1'b0;
  assign \A[5][186] [4] = 1'b0;
  assign \A[5][186] [3] = 1'b0;
  assign \A[5][186] [2] = 1'b0;
  assign \A[5][186] [1] = 1'b0;
  assign \A[5][186] [0] = 1'b0;
  assign \A[5][187] [4] = 1'b0;
  assign \A[5][187] [3] = 1'b0;
  assign \A[5][187] [2] = 1'b0;
  assign \A[5][187] [0] = 1'b0;
  assign \A[5][188] [4] = 1'b0;
  assign \A[5][188] [3] = 1'b0;
  assign \A[5][188] [2] = 1'b0;
  assign \A[5][188] [1] = 1'b0;
  assign \A[5][189] [4] = 1'b0;
  assign \A[5][189] [3] = 1'b0;
  assign \A[5][189] [2] = 1'b0;
  assign \A[5][189] [0] = 1'b0;
  assign \A[5][190] [4] = 1'b0;
  assign \A[5][190] [3] = 1'b0;
  assign \A[5][190] [2] = 1'b0;
  assign \A[5][190] [1] = 1'b0;
  assign \A[5][191] [1] = 1'b0;
  assign \A[5][192] [1] = 1'b0;
  assign \A[5][192] [0] = 1'b0;
  assign \A[5][193] [4] = 1'b0;
  assign \A[5][193] [3] = 1'b0;
  assign \A[5][193] [2] = 1'b0;
  assign \A[5][193] [1] = 1'b0;
  assign \A[5][194] [4] = 1'b0;
  assign \A[5][194] [3] = 1'b0;
  assign \A[5][194] [2] = 1'b0;
  assign \A[5][194] [1] = 1'b0;
  assign \A[5][194] [0] = 1'b0;
  assign \A[5][195] [4] = 1'b0;
  assign \A[5][195] [3] = 1'b0;
  assign \A[5][195] [2] = 1'b0;
  assign \A[5][195] [1] = 1'b0;
  assign \A[5][195] [0] = 1'b0;
  assign \A[5][196] [4] = 1'b0;
  assign \A[5][196] [3] = 1'b0;
  assign \A[5][196] [2] = 1'b0;
  assign \A[5][197] [4] = 1'b0;
  assign \A[5][197] [3] = 1'b0;
  assign \A[5][197] [2] = 1'b0;
  assign \A[5][197] [1] = 1'b0;
  assign \A[5][198] [4] = 1'b0;
  assign \A[5][198] [3] = 1'b0;
  assign \A[5][198] [2] = 1'b0;
  assign \A[5][198] [1] = 1'b0;
  assign \A[5][199] [4] = 1'b0;
  assign \A[5][199] [3] = 1'b0;
  assign \A[5][199] [2] = 1'b0;
  assign \A[5][199] [1] = 1'b0;
  assign \A[5][199] [0] = 1'b0;
  assign \A[5][200] [4] = 1'b0;
  assign \A[5][200] [3] = 1'b0;
  assign \A[5][200] [2] = 1'b0;
  assign \A[5][200] [1] = 1'b0;
  assign \A[5][201] [4] = 1'b0;
  assign \A[5][201] [3] = 1'b0;
  assign \A[5][201] [2] = 1'b0;
  assign \A[5][201] [1] = 1'b0;
  assign \A[5][202] [0] = 1'b0;
  assign \A[5][203] [4] = 1'b0;
  assign \A[5][203] [3] = 1'b0;
  assign \A[5][203] [2] = 1'b0;
  assign \A[5][203] [1] = 1'b0;
  assign \A[5][204] [4] = 1'b0;
  assign \A[5][204] [3] = 1'b0;
  assign \A[5][204] [2] = 1'b0;
  assign \A[5][204] [1] = 1'b0;
  assign \A[5][204] [0] = 1'b0;
  assign \A[5][206] [0] = 1'b0;
  assign \A[5][207] [4] = 1'b0;
  assign \A[5][207] [3] = 1'b0;
  assign \A[5][207] [2] = 1'b0;
  assign \A[5][207] [1] = 1'b0;
  assign \A[5][207] [0] = 1'b0;
  assign \A[5][209] [0] = 1'b0;
  assign \A[5][210] [0] = 1'b0;
  assign \A[5][211] [4] = 1'b0;
  assign \A[5][211] [3] = 1'b0;
  assign \A[5][211] [2] = 1'b0;
  assign \A[5][211] [1] = 1'b0;
  assign \A[5][211] [0] = 1'b0;
  assign \A[5][212] [4] = 1'b0;
  assign \A[5][212] [3] = 1'b0;
  assign \A[5][212] [1] = 1'b0;
  assign \A[5][212] [0] = 1'b0;
  assign \A[5][213] [4] = 1'b0;
  assign \A[5][213] [3] = 1'b0;
  assign \A[5][213] [2] = 1'b0;
  assign \A[5][213] [1] = 1'b0;
  assign \A[5][213] [0] = 1'b0;
  assign \A[5][215] [4] = 1'b0;
  assign \A[5][215] [3] = 1'b0;
  assign \A[5][215] [2] = 1'b0;
  assign \A[5][215] [1] = 1'b0;
  assign \A[5][216] [0] = 1'b0;
  assign \A[5][217] [4] = 1'b0;
  assign \A[5][217] [3] = 1'b0;
  assign \A[5][217] [2] = 1'b0;
  assign \A[5][217] [1] = 1'b0;
  assign \A[5][218] [4] = 1'b0;
  assign \A[5][218] [3] = 1'b0;
  assign \A[5][218] [2] = 1'b0;
  assign \A[5][218] [1] = 1'b0;
  assign \A[5][218] [0] = 1'b0;
  assign \A[5][219] [4] = 1'b0;
  assign \A[5][219] [3] = 1'b0;
  assign \A[5][219] [2] = 1'b0;
  assign \A[5][219] [0] = 1'b0;
  assign \A[5][220] [4] = 1'b0;
  assign \A[5][220] [3] = 1'b0;
  assign \A[5][220] [2] = 1'b0;
  assign \A[5][220] [1] = 1'b0;
  assign \A[5][220] [0] = 1'b0;
  assign \A[5][221] [0] = 1'b0;
  assign \A[5][222] [4] = 1'b0;
  assign \A[5][222] [3] = 1'b0;
  assign \A[5][222] [2] = 1'b0;
  assign \A[5][222] [1] = 1'b0;
  assign \A[5][223] [0] = 1'b0;
  assign \A[5][224] [4] = 1'b0;
  assign \A[5][224] [3] = 1'b0;
  assign \A[5][224] [2] = 1'b0;
  assign \A[5][224] [1] = 1'b0;
  assign \A[5][225] [4] = 1'b0;
  assign \A[5][225] [3] = 1'b0;
  assign \A[5][225] [2] = 1'b0;
  assign \A[5][225] [1] = 1'b0;
  assign \A[5][229] [4] = 1'b0;
  assign \A[5][229] [3] = 1'b0;
  assign \A[5][229] [2] = 1'b0;
  assign \A[5][229] [1] = 1'b0;
  assign \A[5][229] [0] = 1'b0;
  assign \A[5][232] [4] = 1'b0;
  assign \A[5][232] [3] = 1'b0;
  assign \A[5][232] [2] = 1'b0;
  assign \A[5][232] [1] = 1'b0;
  assign \A[5][233] [4] = 1'b0;
  assign \A[5][233] [3] = 1'b0;
  assign \A[5][233] [2] = 1'b0;
  assign \A[5][234] [4] = 1'b0;
  assign \A[5][234] [3] = 1'b0;
  assign \A[5][234] [2] = 1'b0;
  assign \A[5][234] [0] = 1'b0;
  assign \A[5][235] [0] = 1'b0;
  assign \A[5][236] [0] = 1'b0;
  assign \A[5][237] [1] = 1'b0;
  assign \A[5][239] [4] = 1'b0;
  assign \A[5][239] [3] = 1'b0;
  assign \A[5][239] [2] = 1'b0;
  assign \A[5][239] [1] = 1'b0;
  assign \A[5][239] [0] = 1'b0;
  assign \A[5][240] [1] = 1'b0;
  assign \A[5][241] [0] = 1'b0;
  assign \A[5][242] [0] = 1'b0;
  assign \A[5][243] [0] = 1'b0;
  assign \A[5][244] [4] = 1'b0;
  assign \A[5][244] [3] = 1'b0;
  assign \A[5][244] [2] = 1'b0;
  assign \A[5][244] [1] = 1'b0;
  assign \A[5][246] [4] = 1'b0;
  assign \A[5][246] [3] = 1'b0;
  assign \A[5][246] [2] = 1'b0;
  assign \A[5][246] [1] = 1'b0;
  assign \A[5][247] [4] = 1'b0;
  assign \A[5][247] [3] = 1'b0;
  assign \A[5][247] [2] = 1'b0;
  assign \A[5][247] [1] = 1'b0;
  assign \A[5][247] [0] = 1'b0;
  assign \A[5][249] [4] = 1'b0;
  assign \A[5][249] [3] = 1'b0;
  assign \A[5][249] [2] = 1'b0;
  assign \A[5][249] [1] = 1'b0;
  assign \A[5][249] [0] = 1'b0;
  assign \A[5][250] [4] = 1'b0;
  assign \A[5][250] [3] = 1'b0;
  assign \A[5][250] [2] = 1'b0;
  assign \A[5][250] [1] = 1'b0;
  assign \A[5][251] [4] = 1'b0;
  assign \A[5][251] [3] = 1'b0;
  assign \A[5][251] [2] = 1'b0;
  assign \A[5][251] [1] = 1'b0;
  assign \A[5][252] [4] = 1'b0;
  assign \A[5][252] [3] = 1'b0;
  assign \A[5][252] [2] = 1'b0;
  assign \A[5][252] [1] = 1'b0;
  assign \A[5][253] [4] = 1'b0;
  assign \A[5][253] [3] = 1'b0;
  assign \A[5][253] [2] = 1'b0;
  assign \A[5][253] [1] = 1'b0;
  assign \A[5][253] [0] = 1'b0;
  assign \A[6][0] [4] = 1'b0;
  assign \A[6][0] [3] = 1'b0;
  assign \A[6][0] [2] = 1'b0;
  assign \A[6][0] [0] = 1'b0;
  assign \A[6][1] [4] = 1'b0;
  assign \A[6][1] [3] = 1'b0;
  assign \A[6][1] [2] = 1'b0;
  assign \A[6][1] [1] = 1'b0;
  assign \A[6][3] [4] = 1'b0;
  assign \A[6][3] [3] = 1'b0;
  assign \A[6][3] [2] = 1'b0;
  assign \A[6][3] [1] = 1'b0;
  assign \A[6][3] [0] = 1'b0;
  assign \A[6][4] [4] = 1'b0;
  assign \A[6][4] [3] = 1'b0;
  assign \A[6][4] [2] = 1'b0;
  assign \A[6][4] [1] = 1'b0;
  assign \A[6][4] [0] = 1'b0;
  assign \A[6][5] [4] = 1'b0;
  assign \A[6][5] [3] = 1'b0;
  assign \A[6][5] [2] = 1'b0;
  assign \A[6][5] [1] = 1'b0;
  assign \A[6][5] [0] = 1'b0;
  assign \A[6][6] [4] = 1'b0;
  assign \A[6][6] [3] = 1'b0;
  assign \A[6][6] [2] = 1'b0;
  assign \A[6][6] [1] = 1'b0;
  assign \A[6][6] [0] = 1'b0;
  assign \A[6][7] [1] = 1'b0;
  assign \A[6][8] [4] = 1'b0;
  assign \A[6][8] [3] = 1'b0;
  assign \A[6][8] [2] = 1'b0;
  assign \A[6][9] [4] = 1'b0;
  assign \A[6][9] [3] = 1'b0;
  assign \A[6][9] [2] = 1'b0;
  assign \A[6][9] [1] = 1'b0;
  assign \A[6][10] [4] = 1'b0;
  assign \A[6][10] [3] = 1'b0;
  assign \A[6][10] [2] = 1'b0;
  assign \A[6][11] [4] = 1'b0;
  assign \A[6][11] [3] = 1'b0;
  assign \A[6][11] [2] = 1'b0;
  assign \A[6][12] [4] = 1'b0;
  assign \A[6][12] [3] = 1'b0;
  assign \A[6][12] [2] = 1'b0;
  assign \A[6][12] [0] = 1'b0;
  assign \A[6][13] [0] = 1'b0;
  assign \A[6][14] [0] = 1'b0;
  assign \A[6][15] [0] = 1'b0;
  assign \A[6][17] [4] = 1'b0;
  assign \A[6][17] [3] = 1'b0;
  assign \A[6][17] [2] = 1'b0;
  assign \A[6][17] [1] = 1'b0;
  assign \A[6][18] [4] = 1'b0;
  assign \A[6][18] [3] = 1'b0;
  assign \A[6][18] [2] = 1'b0;
  assign \A[6][18] [1] = 1'b0;
  assign \A[6][18] [0] = 1'b0;
  assign \A[6][19] [4] = 1'b0;
  assign \A[6][19] [3] = 1'b0;
  assign \A[6][19] [2] = 1'b0;
  assign \A[6][19] [1] = 1'b0;
  assign \A[6][19] [0] = 1'b0;
  assign \A[6][20] [4] = 1'b0;
  assign \A[6][20] [3] = 1'b0;
  assign \A[6][20] [2] = 1'b0;
  assign \A[6][20] [1] = 1'b0;
  assign \A[6][20] [0] = 1'b0;
  assign \A[6][21] [4] = 1'b0;
  assign \A[6][21] [3] = 1'b0;
  assign \A[6][21] [2] = 1'b0;
  assign \A[6][21] [1] = 1'b0;
  assign \A[6][22] [4] = 1'b0;
  assign \A[6][22] [3] = 1'b0;
  assign \A[6][22] [2] = 1'b0;
  assign \A[6][22] [1] = 1'b0;
  assign \A[6][22] [0] = 1'b0;
  assign \A[6][23] [4] = 1'b0;
  assign \A[6][23] [3] = 1'b0;
  assign \A[6][23] [2] = 1'b0;
  assign \A[6][23] [0] = 1'b0;
  assign \A[6][24] [4] = 1'b0;
  assign \A[6][24] [3] = 1'b0;
  assign \A[6][24] [2] = 1'b0;
  assign \A[6][24] [1] = 1'b0;
  assign \A[6][25] [0] = 1'b0;
  assign \A[6][26] [4] = 1'b0;
  assign \A[6][26] [3] = 1'b0;
  assign \A[6][26] [1] = 1'b0;
  assign \A[6][26] [0] = 1'b0;
  assign \A[6][27] [4] = 1'b0;
  assign \A[6][27] [3] = 1'b0;
  assign \A[6][27] [2] = 1'b0;
  assign \A[6][27] [1] = 1'b0;
  assign \A[6][27] [0] = 1'b0;
  assign \A[6][28] [1] = 1'b0;
  assign \A[6][29] [4] = 1'b0;
  assign \A[6][29] [3] = 1'b0;
  assign \A[6][29] [2] = 1'b0;
  assign \A[6][29] [1] = 1'b0;
  assign \A[6][29] [0] = 1'b0;
  assign \A[6][31] [4] = 1'b0;
  assign \A[6][31] [3] = 1'b0;
  assign \A[6][31] [2] = 1'b0;
  assign \A[6][31] [1] = 1'b0;
  assign \A[6][33] [4] = 1'b0;
  assign \A[6][33] [3] = 1'b0;
  assign \A[6][33] [2] = 1'b0;
  assign \A[6][33] [0] = 1'b0;
  assign \A[6][34] [4] = 1'b0;
  assign \A[6][34] [3] = 1'b0;
  assign \A[6][34] [2] = 1'b0;
  assign \A[6][34] [1] = 1'b0;
  assign \A[6][35] [4] = 1'b0;
  assign \A[6][35] [3] = 1'b0;
  assign \A[6][35] [2] = 1'b0;
  assign \A[6][35] [1] = 1'b0;
  assign \A[6][36] [4] = 1'b0;
  assign \A[6][36] [3] = 1'b0;
  assign \A[6][36] [2] = 1'b0;
  assign \A[6][36] [1] = 1'b0;
  assign \A[6][36] [0] = 1'b0;
  assign \A[6][37] [4] = 1'b0;
  assign \A[6][37] [3] = 1'b0;
  assign \A[6][37] [2] = 1'b0;
  assign \A[6][37] [1] = 1'b0;
  assign \A[6][38] [4] = 1'b0;
  assign \A[6][38] [3] = 1'b0;
  assign \A[6][38] [2] = 1'b0;
  assign \A[6][38] [1] = 1'b0;
  assign \A[6][38] [0] = 1'b0;
  assign \A[6][39] [4] = 1'b0;
  assign \A[6][39] [3] = 1'b0;
  assign \A[6][39] [2] = 1'b0;
  assign \A[6][39] [1] = 1'b0;
  assign \A[6][39] [0] = 1'b0;
  assign \A[6][40] [4] = 1'b0;
  assign \A[6][40] [3] = 1'b0;
  assign \A[6][40] [2] = 1'b0;
  assign \A[6][40] [1] = 1'b0;
  assign \A[6][41] [1] = 1'b0;
  assign \A[6][42] [4] = 1'b0;
  assign \A[6][42] [3] = 1'b0;
  assign \A[6][42] [2] = 1'b0;
  assign \A[6][42] [1] = 1'b0;
  assign \A[6][42] [0] = 1'b0;
  assign \A[6][43] [4] = 1'b0;
  assign \A[6][43] [3] = 1'b0;
  assign \A[6][43] [2] = 1'b0;
  assign \A[6][43] [1] = 1'b0;
  assign \A[6][44] [4] = 1'b0;
  assign \A[6][44] [3] = 1'b0;
  assign \A[6][44] [2] = 1'b0;
  assign \A[6][44] [1] = 1'b0;
  assign \A[6][44] [0] = 1'b0;
  assign \A[6][46] [4] = 1'b0;
  assign \A[6][46] [3] = 1'b0;
  assign \A[6][46] [2] = 1'b0;
  assign \A[6][49] [4] = 1'b0;
  assign \A[6][49] [3] = 1'b0;
  assign \A[6][49] [2] = 1'b0;
  assign \A[6][50] [4] = 1'b0;
  assign \A[6][50] [3] = 1'b0;
  assign \A[6][50] [2] = 1'b0;
  assign \A[6][50] [1] = 1'b0;
  assign \A[6][50] [0] = 1'b0;
  assign \A[6][51] [4] = 1'b0;
  assign \A[6][51] [3] = 1'b0;
  assign \A[6][51] [2] = 1'b0;
  assign \A[6][51] [0] = 1'b0;
  assign \A[6][52] [4] = 1'b0;
  assign \A[6][52] [3] = 1'b0;
  assign \A[6][52] [2] = 1'b0;
  assign \A[6][52] [1] = 1'b0;
  assign \A[6][53] [4] = 1'b0;
  assign \A[6][53] [3] = 1'b0;
  assign \A[6][53] [2] = 1'b0;
  assign \A[6][53] [1] = 1'b0;
  assign \A[6][54] [4] = 1'b0;
  assign \A[6][54] [3] = 1'b0;
  assign \A[6][54] [2] = 1'b0;
  assign \A[6][54] [1] = 1'b0;
  assign \A[6][54] [0] = 1'b0;
  assign \A[6][55] [4] = 1'b0;
  assign \A[6][55] [3] = 1'b0;
  assign \A[6][55] [2] = 1'b0;
  assign \A[6][55] [1] = 1'b0;
  assign \A[6][55] [0] = 1'b0;
  assign \A[6][56] [4] = 1'b0;
  assign \A[6][56] [3] = 1'b0;
  assign \A[6][56] [2] = 1'b0;
  assign \A[6][56] [1] = 1'b0;
  assign \A[6][60] [4] = 1'b0;
  assign \A[6][60] [3] = 1'b0;
  assign \A[6][60] [2] = 1'b0;
  assign \A[6][61] [4] = 1'b0;
  assign \A[6][61] [3] = 1'b0;
  assign \A[6][61] [2] = 1'b0;
  assign \A[6][61] [1] = 1'b0;
  assign \A[6][62] [4] = 1'b0;
  assign \A[6][62] [3] = 1'b0;
  assign \A[6][62] [2] = 1'b0;
  assign \A[6][62] [1] = 1'b0;
  assign \A[6][62] [0] = 1'b0;
  assign \A[6][63] [4] = 1'b0;
  assign \A[6][63] [3] = 1'b0;
  assign \A[6][63] [2] = 1'b0;
  assign \A[6][63] [0] = 1'b0;
  assign \A[6][64] [4] = 1'b0;
  assign \A[6][64] [3] = 1'b0;
  assign \A[6][64] [2] = 1'b0;
  assign \A[6][64] [1] = 1'b0;
  assign \A[6][65] [4] = 1'b0;
  assign \A[6][65] [3] = 1'b0;
  assign \A[6][65] [2] = 1'b0;
  assign \A[6][66] [4] = 1'b0;
  assign \A[6][66] [3] = 1'b0;
  assign \A[6][66] [2] = 1'b0;
  assign \A[6][67] [4] = 1'b0;
  assign \A[6][67] [3] = 1'b0;
  assign \A[6][67] [2] = 1'b0;
  assign \A[6][67] [1] = 1'b0;
  assign \A[6][68] [4] = 1'b0;
  assign \A[6][68] [3] = 1'b0;
  assign \A[6][68] [2] = 1'b0;
  assign \A[6][68] [1] = 1'b0;
  assign \A[6][68] [0] = 1'b0;
  assign \A[6][69] [4] = 1'b0;
  assign \A[6][69] [3] = 1'b0;
  assign \A[6][69] [2] = 1'b0;
  assign \A[6][69] [1] = 1'b0;
  assign \A[6][70] [4] = 1'b0;
  assign \A[6][70] [3] = 1'b0;
  assign \A[6][70] [2] = 1'b0;
  assign \A[6][70] [1] = 1'b0;
  assign \A[6][70] [0] = 1'b0;
  assign \A[6][71] [4] = 1'b0;
  assign \A[6][71] [3] = 1'b0;
  assign \A[6][71] [2] = 1'b0;
  assign \A[6][72] [4] = 1'b0;
  assign \A[6][72] [3] = 1'b0;
  assign \A[6][72] [2] = 1'b0;
  assign \A[6][72] [1] = 1'b0;
  assign \A[6][72] [0] = 1'b0;
  assign \A[6][74] [4] = 1'b0;
  assign \A[6][74] [3] = 1'b0;
  assign \A[6][74] [2] = 1'b0;
  assign \A[6][74] [1] = 1'b0;
  assign \A[6][74] [0] = 1'b0;
  assign \A[6][75] [4] = 1'b0;
  assign \A[6][75] [3] = 1'b0;
  assign \A[6][75] [2] = 1'b0;
  assign \A[6][75] [1] = 1'b0;
  assign \A[6][76] [4] = 1'b0;
  assign \A[6][76] [3] = 1'b0;
  assign \A[6][76] [2] = 1'b0;
  assign \A[6][76] [1] = 1'b0;
  assign \A[6][77] [4] = 1'b0;
  assign \A[6][77] [3] = 1'b0;
  assign \A[6][77] [2] = 1'b0;
  assign \A[6][77] [1] = 1'b0;
  assign \A[6][78] [4] = 1'b0;
  assign \A[6][78] [3] = 1'b0;
  assign \A[6][78] [2] = 1'b0;
  assign \A[6][78] [1] = 1'b0;
  assign \A[6][78] [0] = 1'b0;
  assign \A[6][79] [4] = 1'b0;
  assign \A[6][79] [3] = 1'b0;
  assign \A[6][79] [1] = 1'b0;
  assign \A[6][79] [0] = 1'b0;
  assign \A[6][80] [4] = 1'b0;
  assign \A[6][80] [3] = 1'b0;
  assign \A[6][80] [2] = 1'b0;
  assign \A[6][80] [1] = 1'b0;
  assign \A[6][80] [0] = 1'b0;
  assign \A[6][81] [4] = 1'b0;
  assign \A[6][81] [3] = 1'b0;
  assign \A[6][81] [2] = 1'b0;
  assign \A[6][82] [4] = 1'b0;
  assign \A[6][82] [3] = 1'b0;
  assign \A[6][82] [2] = 1'b0;
  assign \A[6][82] [0] = 1'b0;
  assign \A[6][83] [4] = 1'b0;
  assign \A[6][83] [3] = 1'b0;
  assign \A[6][83] [2] = 1'b0;
  assign \A[6][83] [1] = 1'b0;
  assign \A[6][84] [4] = 1'b0;
  assign \A[6][84] [3] = 1'b0;
  assign \A[6][84] [2] = 1'b0;
  assign \A[6][84] [0] = 1'b0;
  assign \A[6][85] [4] = 1'b0;
  assign \A[6][85] [3] = 1'b0;
  assign \A[6][85] [2] = 1'b0;
  assign \A[6][86] [4] = 1'b0;
  assign \A[6][86] [3] = 1'b0;
  assign \A[6][86] [2] = 1'b0;
  assign \A[6][87] [0] = 1'b0;
  assign \A[6][88] [4] = 1'b0;
  assign \A[6][88] [3] = 1'b0;
  assign \A[6][88] [2] = 1'b0;
  assign \A[6][88] [1] = 1'b0;
  assign \A[6][88] [0] = 1'b0;
  assign \A[6][89] [4] = 1'b0;
  assign \A[6][89] [3] = 1'b0;
  assign \A[6][89] [2] = 1'b0;
  assign \A[6][89] [1] = 1'b0;
  assign \A[6][89] [0] = 1'b0;
  assign \A[6][90] [0] = 1'b0;
  assign \A[6][91] [1] = 1'b0;
  assign \A[6][92] [4] = 1'b0;
  assign \A[6][92] [3] = 1'b0;
  assign \A[6][92] [2] = 1'b0;
  assign \A[6][92] [1] = 1'b0;
  assign \A[6][93] [4] = 1'b0;
  assign \A[6][93] [3] = 1'b0;
  assign \A[6][93] [2] = 1'b0;
  assign \A[6][93] [0] = 1'b0;
  assign \A[6][95] [4] = 1'b0;
  assign \A[6][95] [3] = 1'b0;
  assign \A[6][95] [2] = 1'b0;
  assign \A[6][95] [1] = 1'b0;
  assign \A[6][95] [0] = 1'b0;
  assign \A[6][96] [4] = 1'b0;
  assign \A[6][96] [3] = 1'b0;
  assign \A[6][96] [2] = 1'b0;
  assign \A[6][96] [0] = 1'b0;
  assign \A[6][97] [4] = 1'b0;
  assign \A[6][97] [3] = 1'b0;
  assign \A[6][97] [2] = 1'b0;
  assign \A[6][97] [1] = 1'b0;
  assign \A[6][98] [4] = 1'b0;
  assign \A[6][98] [3] = 1'b0;
  assign \A[6][98] [2] = 1'b0;
  assign \A[6][98] [0] = 1'b0;
  assign \A[6][100] [4] = 1'b0;
  assign \A[6][100] [3] = 1'b0;
  assign \A[6][100] [2] = 1'b0;
  assign \A[6][100] [0] = 1'b0;
  assign \A[6][101] [4] = 1'b0;
  assign \A[6][101] [3] = 1'b0;
  assign \A[6][101] [2] = 1'b0;
  assign \A[6][101] [1] = 1'b0;
  assign \A[6][102] [4] = 1'b0;
  assign \A[6][102] [3] = 1'b0;
  assign \A[6][102] [2] = 1'b0;
  assign \A[6][102] [1] = 1'b0;
  assign \A[6][103] [4] = 1'b0;
  assign \A[6][103] [3] = 1'b0;
  assign \A[6][103] [2] = 1'b0;
  assign \A[6][103] [1] = 1'b0;
  assign \A[6][103] [0] = 1'b0;
  assign \A[6][104] [4] = 1'b0;
  assign \A[6][104] [3] = 1'b0;
  assign \A[6][104] [2] = 1'b0;
  assign \A[6][104] [1] = 1'b0;
  assign \A[6][104] [0] = 1'b0;
  assign \A[6][105] [4] = 1'b0;
  assign \A[6][105] [3] = 1'b0;
  assign \A[6][105] [2] = 1'b0;
  assign \A[6][106] [4] = 1'b0;
  assign \A[6][106] [3] = 1'b0;
  assign \A[6][106] [2] = 1'b0;
  assign \A[6][106] [1] = 1'b0;
  assign \A[6][107] [4] = 1'b0;
  assign \A[6][107] [3] = 1'b0;
  assign \A[6][107] [2] = 1'b0;
  assign \A[6][107] [0] = 1'b0;
  assign \A[6][108] [4] = 1'b0;
  assign \A[6][108] [3] = 1'b0;
  assign \A[6][108] [2] = 1'b0;
  assign \A[6][108] [1] = 1'b0;
  assign \A[6][108] [0] = 1'b0;
  assign \A[6][109] [4] = 1'b0;
  assign \A[6][109] [3] = 1'b0;
  assign \A[6][109] [2] = 1'b0;
  assign \A[6][109] [0] = 1'b0;
  assign \A[6][110] [4] = 1'b0;
  assign \A[6][110] [3] = 1'b0;
  assign \A[6][110] [2] = 1'b0;
  assign \A[6][110] [0] = 1'b0;
  assign \A[6][111] [4] = 1'b0;
  assign \A[6][111] [3] = 1'b0;
  assign \A[6][111] [2] = 1'b0;
  assign \A[6][111] [1] = 1'b0;
  assign \A[6][112] [4] = 1'b0;
  assign \A[6][112] [3] = 1'b0;
  assign \A[6][112] [2] = 1'b0;
  assign \A[6][112] [1] = 1'b0;
  assign \A[6][113] [4] = 1'b0;
  assign \A[6][113] [3] = 1'b0;
  assign \A[6][113] [2] = 1'b0;
  assign \A[6][113] [0] = 1'b0;
  assign \A[6][114] [4] = 1'b0;
  assign \A[6][114] [3] = 1'b0;
  assign \A[6][114] [2] = 1'b0;
  assign \A[6][115] [4] = 1'b0;
  assign \A[6][115] [3] = 1'b0;
  assign \A[6][115] [2] = 1'b0;
  assign \A[6][115] [1] = 1'b0;
  assign \A[6][116] [4] = 1'b0;
  assign \A[6][116] [3] = 1'b0;
  assign \A[6][116] [2] = 1'b0;
  assign \A[6][116] [1] = 1'b0;
  assign \A[6][116] [0] = 1'b0;
  assign \A[6][117] [4] = 1'b0;
  assign \A[6][117] [3] = 1'b0;
  assign \A[6][117] [2] = 1'b0;
  assign \A[6][117] [0] = 1'b0;
  assign \A[6][119] [4] = 1'b0;
  assign \A[6][119] [3] = 1'b0;
  assign \A[6][119] [2] = 1'b0;
  assign \A[6][119] [1] = 1'b0;
  assign \A[6][121] [4] = 1'b0;
  assign \A[6][121] [3] = 1'b0;
  assign \A[6][121] [2] = 1'b0;
  assign \A[6][122] [0] = 1'b0;
  assign \A[6][123] [4] = 1'b0;
  assign \A[6][123] [3] = 1'b0;
  assign \A[6][123] [2] = 1'b0;
  assign \A[6][123] [1] = 1'b0;
  assign \A[6][123] [0] = 1'b0;
  assign \A[6][124] [4] = 1'b0;
  assign \A[6][124] [3] = 1'b0;
  assign \A[6][124] [2] = 1'b0;
  assign \A[6][124] [1] = 1'b0;
  assign \A[6][124] [0] = 1'b0;
  assign \A[6][127] [4] = 1'b0;
  assign \A[6][127] [3] = 1'b0;
  assign \A[6][127] [2] = 1'b0;
  assign \A[6][127] [0] = 1'b0;
  assign \A[6][129] [4] = 1'b0;
  assign \A[6][129] [3] = 1'b0;
  assign \A[6][129] [2] = 1'b0;
  assign \A[6][129] [0] = 1'b0;
  assign \A[6][130] [4] = 1'b0;
  assign \A[6][130] [3] = 1'b0;
  assign \A[6][130] [2] = 1'b0;
  assign \A[6][130] [1] = 1'b0;
  assign \A[6][130] [0] = 1'b0;
  assign \A[6][131] [4] = 1'b0;
  assign \A[6][131] [3] = 1'b0;
  assign \A[6][131] [2] = 1'b0;
  assign \A[6][131] [1] = 1'b0;
  assign \A[6][132] [4] = 1'b0;
  assign \A[6][132] [3] = 1'b0;
  assign \A[6][132] [2] = 1'b0;
  assign \A[6][132] [0] = 1'b0;
  assign \A[6][134] [4] = 1'b0;
  assign \A[6][134] [3] = 1'b0;
  assign \A[6][134] [2] = 1'b0;
  assign \A[6][134] [1] = 1'b0;
  assign \A[6][134] [0] = 1'b0;
  assign \A[6][135] [0] = 1'b0;
  assign \A[6][136] [4] = 1'b0;
  assign \A[6][136] [3] = 1'b0;
  assign \A[6][136] [2] = 1'b0;
  assign \A[6][136] [1] = 1'b0;
  assign \A[6][137] [4] = 1'b0;
  assign \A[6][137] [3] = 1'b0;
  assign \A[6][137] [2] = 1'b0;
  assign \A[6][137] [1] = 1'b0;
  assign \A[6][137] [0] = 1'b0;
  assign \A[6][138] [0] = 1'b0;
  assign \A[6][139] [4] = 1'b0;
  assign \A[6][139] [3] = 1'b0;
  assign \A[6][139] [2] = 1'b0;
  assign \A[6][139] [0] = 1'b0;
  assign \A[6][140] [0] = 1'b0;
  assign \A[6][141] [4] = 1'b0;
  assign \A[6][141] [3] = 1'b0;
  assign \A[6][141] [2] = 1'b0;
  assign \A[6][141] [1] = 1'b0;
  assign \A[6][141] [0] = 1'b0;
  assign \A[6][142] [4] = 1'b0;
  assign \A[6][142] [3] = 1'b0;
  assign \A[6][142] [2] = 1'b0;
  assign \A[6][142] [1] = 1'b0;
  assign \A[6][143] [4] = 1'b0;
  assign \A[6][143] [3] = 1'b0;
  assign \A[6][143] [2] = 1'b0;
  assign \A[6][143] [0] = 1'b0;
  assign \A[6][144] [4] = 1'b0;
  assign \A[6][144] [3] = 1'b0;
  assign \A[6][144] [2] = 1'b0;
  assign \A[6][146] [4] = 1'b0;
  assign \A[6][146] [3] = 1'b0;
  assign \A[6][146] [2] = 1'b0;
  assign \A[6][146] [1] = 1'b0;
  assign \A[6][147] [4] = 1'b0;
  assign \A[6][147] [3] = 1'b0;
  assign \A[6][147] [2] = 1'b0;
  assign \A[6][147] [1] = 1'b0;
  assign \A[6][147] [0] = 1'b0;
  assign \A[6][149] [4] = 1'b0;
  assign \A[6][149] [3] = 1'b0;
  assign \A[6][149] [2] = 1'b0;
  assign \A[6][149] [1] = 1'b0;
  assign \A[6][149] [0] = 1'b0;
  assign \A[6][152] [4] = 1'b0;
  assign \A[6][152] [3] = 1'b0;
  assign \A[6][152] [2] = 1'b0;
  assign \A[6][152] [1] = 1'b0;
  assign \A[6][152] [0] = 1'b0;
  assign \A[6][153] [0] = 1'b0;
  assign \A[6][154] [4] = 1'b0;
  assign \A[6][154] [3] = 1'b0;
  assign \A[6][154] [2] = 1'b0;
  assign \A[6][154] [1] = 1'b0;
  assign \A[6][155] [4] = 1'b0;
  assign \A[6][155] [3] = 1'b0;
  assign \A[6][155] [2] = 1'b0;
  assign \A[6][155] [0] = 1'b0;
  assign \A[6][156] [4] = 1'b0;
  assign \A[6][156] [3] = 1'b0;
  assign \A[6][156] [2] = 1'b0;
  assign \A[6][156] [1] = 1'b0;
  assign \A[6][157] [0] = 1'b0;
  assign \A[6][159] [4] = 1'b0;
  assign \A[6][159] [3] = 1'b0;
  assign \A[6][159] [2] = 1'b0;
  assign \A[6][159] [1] = 1'b0;
  assign \A[6][160] [4] = 1'b0;
  assign \A[6][160] [3] = 1'b0;
  assign \A[6][160] [2] = 1'b0;
  assign \A[6][160] [1] = 1'b0;
  assign \A[6][162] [4] = 1'b0;
  assign \A[6][162] [3] = 1'b0;
  assign \A[6][162] [2] = 1'b0;
  assign \A[6][162] [1] = 1'b0;
  assign \A[6][162] [0] = 1'b0;
  assign \A[6][164] [0] = 1'b0;
  assign \A[6][165] [4] = 1'b0;
  assign \A[6][165] [3] = 1'b0;
  assign \A[6][165] [2] = 1'b0;
  assign \A[6][165] [1] = 1'b0;
  assign \A[6][166] [4] = 1'b0;
  assign \A[6][166] [3] = 1'b0;
  assign \A[6][166] [2] = 1'b0;
  assign \A[6][166] [1] = 1'b0;
  assign \A[6][166] [0] = 1'b0;
  assign \A[6][167] [4] = 1'b0;
  assign \A[6][167] [3] = 1'b0;
  assign \A[6][167] [2] = 1'b0;
  assign \A[6][167] [1] = 1'b0;
  assign \A[6][168] [4] = 1'b0;
  assign \A[6][168] [3] = 1'b0;
  assign \A[6][168] [2] = 1'b0;
  assign \A[6][168] [1] = 1'b0;
  assign \A[6][169] [4] = 1'b0;
  assign \A[6][169] [3] = 1'b0;
  assign \A[6][169] [2] = 1'b0;
  assign \A[6][169] [1] = 1'b0;
  assign \A[6][169] [0] = 1'b0;
  assign \A[6][170] [1] = 1'b0;
  assign \A[6][171] [4] = 1'b0;
  assign \A[6][171] [3] = 1'b0;
  assign \A[6][171] [2] = 1'b0;
  assign \A[6][172] [4] = 1'b0;
  assign \A[6][172] [3] = 1'b0;
  assign \A[6][172] [2] = 1'b0;
  assign \A[6][173] [4] = 1'b0;
  assign \A[6][173] [3] = 1'b0;
  assign \A[6][173] [2] = 1'b0;
  assign \A[6][173] [0] = 1'b0;
  assign \A[6][174] [4] = 1'b0;
  assign \A[6][174] [3] = 1'b0;
  assign \A[6][174] [2] = 1'b0;
  assign \A[6][174] [1] = 1'b0;
  assign \A[6][174] [0] = 1'b0;
  assign \A[6][176] [4] = 1'b0;
  assign \A[6][176] [3] = 1'b0;
  assign \A[6][176] [2] = 1'b0;
  assign \A[6][176] [1] = 1'b0;
  assign \A[6][176] [0] = 1'b0;
  assign \A[6][179] [1] = 1'b0;
  assign \A[6][179] [0] = 1'b0;
  assign \A[6][180] [1] = 1'b0;
  assign \A[6][180] [0] = 1'b0;
  assign \A[6][181] [4] = 1'b0;
  assign \A[6][181] [3] = 1'b0;
  assign \A[6][181] [2] = 1'b0;
  assign \A[6][181] [1] = 1'b0;
  assign \A[6][181] [0] = 1'b0;
  assign \A[6][182] [0] = 1'b0;
  assign \A[6][183] [1] = 1'b0;
  assign \A[6][183] [0] = 1'b0;
  assign \A[6][184] [4] = 1'b0;
  assign \A[6][184] [3] = 1'b0;
  assign \A[6][184] [2] = 1'b0;
  assign \A[6][184] [1] = 1'b0;
  assign \A[6][185] [4] = 1'b0;
  assign \A[6][185] [3] = 1'b0;
  assign \A[6][185] [2] = 1'b0;
  assign \A[6][185] [0] = 1'b0;
  assign \A[6][186] [4] = 1'b0;
  assign \A[6][186] [3] = 1'b0;
  assign \A[6][186] [2] = 1'b0;
  assign \A[6][186] [1] = 1'b0;
  assign \A[6][186] [0] = 1'b0;
  assign \A[6][187] [0] = 1'b0;
  assign \A[6][188] [0] = 1'b0;
  assign \A[6][189] [4] = 1'b0;
  assign \A[6][189] [3] = 1'b0;
  assign \A[6][189] [2] = 1'b0;
  assign \A[6][189] [1] = 1'b0;
  assign \A[6][191] [4] = 1'b0;
  assign \A[6][191] [3] = 1'b0;
  assign \A[6][191] [2] = 1'b0;
  assign \A[6][191] [1] = 1'b0;
  assign \A[6][192] [4] = 1'b0;
  assign \A[6][192] [3] = 1'b0;
  assign \A[6][192] [2] = 1'b0;
  assign \A[6][192] [1] = 1'b0;
  assign \A[6][192] [0] = 1'b0;
  assign \A[6][194] [1] = 1'b0;
  assign \A[6][195] [4] = 1'b0;
  assign \A[6][195] [3] = 1'b0;
  assign \A[6][195] [2] = 1'b0;
  assign \A[6][195] [1] = 1'b0;
  assign \A[6][196] [0] = 1'b0;
  assign \A[6][197] [0] = 1'b0;
  assign \A[6][198] [0] = 1'b0;
  assign \A[6][199] [4] = 1'b0;
  assign \A[6][199] [3] = 1'b0;
  assign \A[6][199] [2] = 1'b0;
  assign \A[6][199] [1] = 1'b0;
  assign \A[6][199] [0] = 1'b0;
  assign \A[6][200] [4] = 1'b0;
  assign \A[6][200] [3] = 1'b0;
  assign \A[6][200] [2] = 1'b0;
  assign \A[6][200] [1] = 1'b0;
  assign \A[6][202] [4] = 1'b0;
  assign \A[6][202] [3] = 1'b0;
  assign \A[6][202] [2] = 1'b0;
  assign \A[6][202] [1] = 1'b0;
  assign \A[6][202] [0] = 1'b0;
  assign \A[6][205] [0] = 1'b0;
  assign \A[6][206] [4] = 1'b0;
  assign \A[6][206] [3] = 1'b0;
  assign \A[6][206] [2] = 1'b0;
  assign \A[6][206] [1] = 1'b0;
  assign \A[6][207] [4] = 1'b0;
  assign \A[6][207] [3] = 1'b0;
  assign \A[6][207] [2] = 1'b0;
  assign \A[6][207] [0] = 1'b0;
  assign \A[6][208] [4] = 1'b0;
  assign \A[6][208] [3] = 1'b0;
  assign \A[6][208] [2] = 1'b0;
  assign \A[6][208] [1] = 1'b0;
  assign \A[6][209] [4] = 1'b0;
  assign \A[6][209] [3] = 1'b0;
  assign \A[6][209] [2] = 1'b0;
  assign \A[6][209] [1] = 1'b0;
  assign \A[6][211] [4] = 1'b0;
  assign \A[6][211] [3] = 1'b0;
  assign \A[6][211] [2] = 1'b0;
  assign \A[6][211] [0] = 1'b0;
  assign \A[6][212] [4] = 1'b0;
  assign \A[6][212] [3] = 1'b0;
  assign \A[6][212] [2] = 1'b0;
  assign \A[6][212] [1] = 1'b0;
  assign \A[6][212] [0] = 1'b0;
  assign \A[6][213] [4] = 1'b0;
  assign \A[6][213] [3] = 1'b0;
  assign \A[6][213] [2] = 1'b0;
  assign \A[6][213] [0] = 1'b0;
  assign \A[6][214] [4] = 1'b0;
  assign \A[6][214] [3] = 1'b0;
  assign \A[6][214] [2] = 1'b0;
  assign \A[6][214] [1] = 1'b0;
  assign \A[6][214] [0] = 1'b0;
  assign \A[6][215] [0] = 1'b0;
  assign \A[6][216] [4] = 1'b0;
  assign \A[6][216] [3] = 1'b0;
  assign \A[6][216] [2] = 1'b0;
  assign \A[6][216] [1] = 1'b0;
  assign \A[6][216] [0] = 1'b0;
  assign \A[6][219] [4] = 1'b0;
  assign \A[6][219] [3] = 1'b0;
  assign \A[6][219] [2] = 1'b0;
  assign \A[6][219] [1] = 1'b0;
  assign \A[6][219] [0] = 1'b0;
  assign \A[6][220] [4] = 1'b0;
  assign \A[6][220] [3] = 1'b0;
  assign \A[6][220] [2] = 1'b0;
  assign \A[6][220] [1] = 1'b0;
  assign \A[6][221] [0] = 1'b0;
  assign \A[6][222] [1] = 1'b0;
  assign \A[6][224] [4] = 1'b0;
  assign \A[6][224] [3] = 1'b0;
  assign \A[6][224] [2] = 1'b0;
  assign \A[6][224] [1] = 1'b0;
  assign \A[6][224] [0] = 1'b0;
  assign \A[6][225] [4] = 1'b0;
  assign \A[6][225] [3] = 1'b0;
  assign \A[6][225] [2] = 1'b0;
  assign \A[6][225] [1] = 1'b0;
  assign \A[6][229] [1] = 1'b0;
  assign \A[6][230] [4] = 1'b0;
  assign \A[6][230] [3] = 1'b0;
  assign \A[6][230] [2] = 1'b0;
  assign \A[6][230] [1] = 1'b0;
  assign \A[6][231] [1] = 1'b0;
  assign \A[6][232] [4] = 1'b0;
  assign \A[6][232] [3] = 1'b0;
  assign \A[6][232] [2] = 1'b0;
  assign \A[6][232] [1] = 1'b0;
  assign \A[6][232] [0] = 1'b0;
  assign \A[6][234] [1] = 1'b0;
  assign \A[6][235] [4] = 1'b0;
  assign \A[6][235] [3] = 1'b0;
  assign \A[6][235] [2] = 1'b0;
  assign \A[6][235] [1] = 1'b0;
  assign \A[6][235] [0] = 1'b0;
  assign \A[6][236] [4] = 1'b0;
  assign \A[6][236] [3] = 1'b0;
  assign \A[6][236] [2] = 1'b0;
  assign \A[6][236] [1] = 1'b0;
  assign \A[6][236] [0] = 1'b0;
  assign \A[6][237] [0] = 1'b0;
  assign \A[6][238] [1] = 1'b0;
  assign \A[6][239] [0] = 1'b0;
  assign \A[6][240] [4] = 1'b0;
  assign \A[6][240] [3] = 1'b0;
  assign \A[6][240] [2] = 1'b0;
  assign \A[6][240] [1] = 1'b0;
  assign \A[6][241] [4] = 1'b0;
  assign \A[6][241] [3] = 1'b0;
  assign \A[6][241] [2] = 1'b0;
  assign \A[6][241] [1] = 1'b0;
  assign \A[6][242] [4] = 1'b0;
  assign \A[6][242] [3] = 1'b0;
  assign \A[6][242] [2] = 1'b0;
  assign \A[6][242] [1] = 1'b0;
  assign \A[6][243] [4] = 1'b0;
  assign \A[6][243] [3] = 1'b0;
  assign \A[6][243] [2] = 1'b0;
  assign \A[6][243] [1] = 1'b0;
  assign \A[6][245] [4] = 1'b0;
  assign \A[6][245] [3] = 1'b0;
  assign \A[6][245] [2] = 1'b0;
  assign \A[6][245] [1] = 1'b0;
  assign \A[6][245] [0] = 1'b0;
  assign \A[6][246] [4] = 1'b0;
  assign \A[6][246] [3] = 1'b0;
  assign \A[6][246] [2] = 1'b0;
  assign \A[6][248] [4] = 1'b0;
  assign \A[6][248] [3] = 1'b0;
  assign \A[6][248] [2] = 1'b0;
  assign \A[6][248] [1] = 1'b0;
  assign \A[6][248] [0] = 1'b0;
  assign \A[6][249] [4] = 1'b0;
  assign \A[6][249] [3] = 1'b0;
  assign \A[6][249] [2] = 1'b0;
  assign \A[6][249] [1] = 1'b0;
  assign \A[6][249] [0] = 1'b0;
  assign \A[6][250] [4] = 1'b0;
  assign \A[6][250] [3] = 1'b0;
  assign \A[6][250] [2] = 1'b0;
  assign \A[6][250] [1] = 1'b0;
  assign \A[6][251] [4] = 1'b0;
  assign \A[6][251] [3] = 1'b0;
  assign \A[6][251] [2] = 1'b0;
  assign \A[6][251] [0] = 1'b0;
  assign \A[6][252] [0] = 1'b0;
  assign \A[6][253] [4] = 1'b0;
  assign \A[6][253] [3] = 1'b0;
  assign \A[6][253] [2] = 1'b0;
  assign \A[6][253] [0] = 1'b0;
  assign \A[6][255] [1] = 1'b0;
  assign \A[7][2] [4] = 1'b0;
  assign \A[7][2] [3] = 1'b0;
  assign \A[7][2] [2] = 1'b0;
  assign \A[7][2] [1] = 1'b0;
  assign \A[7][2] [0] = 1'b0;
  assign \A[7][3] [4] = 1'b0;
  assign \A[7][3] [3] = 1'b0;
  assign \A[7][3] [2] = 1'b0;
  assign \A[7][3] [1] = 1'b0;
  assign \A[7][3] [0] = 1'b0;
  assign \A[7][4] [0] = 1'b0;
  assign \A[7][5] [4] = 1'b0;
  assign \A[7][5] [3] = 1'b0;
  assign \A[7][5] [2] = 1'b0;
  assign \A[7][5] [1] = 1'b0;
  assign \A[7][5] [0] = 1'b0;
  assign \A[7][6] [4] = 1'b0;
  assign \A[7][6] [3] = 1'b0;
  assign \A[7][6] [2] = 1'b0;
  assign \A[7][6] [0] = 1'b0;
  assign \A[7][7] [4] = 1'b0;
  assign \A[7][7] [3] = 1'b0;
  assign \A[7][7] [2] = 1'b0;
  assign \A[7][7] [1] = 1'b0;
  assign \A[7][8] [0] = 1'b0;
  assign \A[7][10] [4] = 1'b0;
  assign \A[7][10] [3] = 1'b0;
  assign \A[7][10] [2] = 1'b0;
  assign \A[7][10] [1] = 1'b0;
  assign \A[7][12] [4] = 1'b0;
  assign \A[7][12] [3] = 1'b0;
  assign \A[7][12] [2] = 1'b0;
  assign \A[7][12] [0] = 1'b0;
  assign \A[7][15] [4] = 1'b0;
  assign \A[7][15] [3] = 1'b0;
  assign \A[7][15] [2] = 1'b0;
  assign \A[7][15] [0] = 1'b0;
  assign \A[7][16] [4] = 1'b0;
  assign \A[7][16] [3] = 1'b0;
  assign \A[7][16] [2] = 1'b0;
  assign \A[7][16] [1] = 1'b0;
  assign \A[7][17] [4] = 1'b0;
  assign \A[7][17] [3] = 1'b0;
  assign \A[7][17] [2] = 1'b0;
  assign \A[7][17] [1] = 1'b0;
  assign \A[7][18] [0] = 1'b0;
  assign \A[7][19] [4] = 1'b0;
  assign \A[7][19] [3] = 1'b0;
  assign \A[7][19] [2] = 1'b0;
  assign \A[7][19] [1] = 1'b0;
  assign \A[7][19] [0] = 1'b0;
  assign \A[7][20] [4] = 1'b0;
  assign \A[7][20] [3] = 1'b0;
  assign \A[7][20] [2] = 1'b0;
  assign \A[7][20] [1] = 1'b0;
  assign \A[7][20] [0] = 1'b0;
  assign \A[7][21] [0] = 1'b0;
  assign \A[7][23] [4] = 1'b0;
  assign \A[7][23] [3] = 1'b0;
  assign \A[7][23] [2] = 1'b0;
  assign \A[7][23] [1] = 1'b0;
  assign \A[7][24] [4] = 1'b0;
  assign \A[7][24] [3] = 1'b0;
  assign \A[7][24] [2] = 1'b0;
  assign \A[7][24] [1] = 1'b0;
  assign \A[7][25] [4] = 1'b0;
  assign \A[7][25] [3] = 1'b0;
  assign \A[7][25] [1] = 1'b0;
  assign \A[7][25] [0] = 1'b0;
  assign \A[7][26] [1] = 1'b0;
  assign \A[7][27] [4] = 1'b0;
  assign \A[7][27] [3] = 1'b0;
  assign \A[7][27] [2] = 1'b0;
  assign \A[7][27] [1] = 1'b0;
  assign \A[7][27] [0] = 1'b0;
  assign \A[7][28] [4] = 1'b0;
  assign \A[7][28] [3] = 1'b0;
  assign \A[7][28] [2] = 1'b0;
  assign \A[7][28] [1] = 1'b0;
  assign \A[7][29] [1] = 1'b0;
  assign \A[7][30] [4] = 1'b0;
  assign \A[7][30] [3] = 1'b0;
  assign \A[7][30] [2] = 1'b0;
  assign \A[7][30] [1] = 1'b0;
  assign \A[7][30] [0] = 1'b0;
  assign \A[7][31] [4] = 1'b0;
  assign \A[7][31] [3] = 1'b0;
  assign \A[7][31] [2] = 1'b0;
  assign \A[7][31] [0] = 1'b0;
  assign \A[7][32] [4] = 1'b0;
  assign \A[7][32] [3] = 1'b0;
  assign \A[7][32] [2] = 1'b0;
  assign \A[7][32] [1] = 1'b0;
  assign \A[7][32] [0] = 1'b0;
  assign \A[7][33] [4] = 1'b0;
  assign \A[7][33] [3] = 1'b0;
  assign \A[7][33] [2] = 1'b0;
  assign \A[7][33] [1] = 1'b0;
  assign \A[7][33] [0] = 1'b0;
  assign \A[7][34] [4] = 1'b0;
  assign \A[7][34] [3] = 1'b0;
  assign \A[7][34] [2] = 1'b0;
  assign \A[7][34] [1] = 1'b0;
  assign \A[7][34] [0] = 1'b0;
  assign \A[7][35] [4] = 1'b0;
  assign \A[7][35] [3] = 1'b0;
  assign \A[7][35] [2] = 1'b0;
  assign \A[7][35] [1] = 1'b0;
  assign \A[7][36] [4] = 1'b0;
  assign \A[7][36] [3] = 1'b0;
  assign \A[7][36] [2] = 1'b0;
  assign \A[7][36] [1] = 1'b0;
  assign \A[7][36] [0] = 1'b0;
  assign \A[7][37] [4] = 1'b0;
  assign \A[7][37] [3] = 1'b0;
  assign \A[7][37] [2] = 1'b0;
  assign \A[7][37] [1] = 1'b0;
  assign \A[7][37] [0] = 1'b0;
  assign \A[7][38] [0] = 1'b0;
  assign \A[7][39] [1] = 1'b0;
  assign \A[7][41] [0] = 1'b0;
  assign \A[7][42] [0] = 1'b0;
  assign \A[7][44] [4] = 1'b0;
  assign \A[7][44] [3] = 1'b0;
  assign \A[7][44] [2] = 1'b0;
  assign \A[7][44] [1] = 1'b0;
  assign \A[7][45] [4] = 1'b0;
  assign \A[7][45] [3] = 1'b0;
  assign \A[7][45] [2] = 1'b0;
  assign \A[7][45] [1] = 1'b0;
  assign \A[7][47] [4] = 1'b0;
  assign \A[7][47] [3] = 1'b0;
  assign \A[7][47] [2] = 1'b0;
  assign \A[7][47] [1] = 1'b0;
  assign \A[7][48] [4] = 1'b0;
  assign \A[7][48] [3] = 1'b0;
  assign \A[7][48] [2] = 1'b0;
  assign \A[7][48] [1] = 1'b0;
  assign \A[7][49] [0] = 1'b0;
  assign \A[7][50] [4] = 1'b0;
  assign \A[7][50] [3] = 1'b0;
  assign \A[7][50] [2] = 1'b0;
  assign \A[7][50] [0] = 1'b0;
  assign \A[7][51] [1] = 1'b0;
  assign \A[7][52] [4] = 1'b0;
  assign \A[7][52] [3] = 1'b0;
  assign \A[7][52] [2] = 1'b0;
  assign \A[7][52] [1] = 1'b0;
  assign \A[7][53] [4] = 1'b0;
  assign \A[7][53] [3] = 1'b0;
  assign \A[7][53] [2] = 1'b0;
  assign \A[7][53] [1] = 1'b0;
  assign \A[7][53] [0] = 1'b0;
  assign \A[7][54] [4] = 1'b0;
  assign \A[7][54] [3] = 1'b0;
  assign \A[7][54] [2] = 1'b0;
  assign \A[7][54] [1] = 1'b0;
  assign \A[7][54] [0] = 1'b0;
  assign \A[7][55] [4] = 1'b0;
  assign \A[7][55] [3] = 1'b0;
  assign \A[7][55] [2] = 1'b0;
  assign \A[7][55] [1] = 1'b0;
  assign \A[7][57] [1] = 1'b0;
  assign \A[7][57] [0] = 1'b0;
  assign \A[7][58] [2] = 1'b0;
  assign \A[7][59] [0] = 1'b0;
  assign \A[7][60] [4] = 1'b0;
  assign \A[7][60] [3] = 1'b0;
  assign \A[7][60] [2] = 1'b0;
  assign \A[7][60] [1] = 1'b0;
  assign \A[7][60] [0] = 1'b0;
  assign \A[7][61] [4] = 1'b0;
  assign \A[7][61] [3] = 1'b0;
  assign \A[7][61] [2] = 1'b0;
  assign \A[7][61] [1] = 1'b0;
  assign \A[7][61] [0] = 1'b0;
  assign \A[7][62] [1] = 1'b0;
  assign \A[7][63] [0] = 1'b0;
  assign \A[7][64] [0] = 1'b0;
  assign \A[7][65] [4] = 1'b0;
  assign \A[7][65] [3] = 1'b0;
  assign \A[7][65] [2] = 1'b0;
  assign \A[7][65] [0] = 1'b0;
  assign \A[7][66] [4] = 1'b0;
  assign \A[7][66] [3] = 1'b0;
  assign \A[7][66] [2] = 1'b0;
  assign \A[7][66] [1] = 1'b0;
  assign \A[7][68] [4] = 1'b0;
  assign \A[7][68] [3] = 1'b0;
  assign \A[7][68] [2] = 1'b0;
  assign \A[7][68] [1] = 1'b0;
  assign \A[7][70] [0] = 1'b0;
  assign \A[7][71] [4] = 1'b0;
  assign \A[7][71] [3] = 1'b0;
  assign \A[7][71] [2] = 1'b0;
  assign \A[7][71] [1] = 1'b0;
  assign \A[7][72] [4] = 1'b0;
  assign \A[7][72] [3] = 1'b0;
  assign \A[7][72] [2] = 1'b0;
  assign \A[7][72] [1] = 1'b0;
  assign \A[7][73] [1] = 1'b0;
  assign \A[7][74] [2] = 1'b0;
  assign \A[7][75] [1] = 1'b0;
  assign \A[7][76] [0] = 1'b0;
  assign \A[7][77] [1] = 1'b0;
  assign \A[7][78] [0] = 1'b0;
  assign \A[7][79] [4] = 1'b0;
  assign \A[7][79] [3] = 1'b0;
  assign \A[7][79] [2] = 1'b0;
  assign \A[7][79] [1] = 1'b0;
  assign \A[7][79] [0] = 1'b0;
  assign \A[7][81] [0] = 1'b0;
  assign \A[7][83] [0] = 1'b0;
  assign \A[7][84] [0] = 1'b0;
  assign \A[7][85] [4] = 1'b0;
  assign \A[7][85] [3] = 1'b0;
  assign \A[7][85] [2] = 1'b0;
  assign \A[7][85] [1] = 1'b0;
  assign \A[7][86] [4] = 1'b0;
  assign \A[7][86] [3] = 1'b0;
  assign \A[7][86] [1] = 1'b0;
  assign \A[7][87] [4] = 1'b0;
  assign \A[7][87] [3] = 1'b0;
  assign \A[7][87] [2] = 1'b0;
  assign \A[7][87] [1] = 1'b0;
  assign \A[7][88] [4] = 1'b0;
  assign \A[7][88] [3] = 1'b0;
  assign \A[7][88] [2] = 1'b0;
  assign \A[7][88] [1] = 1'b0;
  assign \A[7][89] [4] = 1'b0;
  assign \A[7][89] [3] = 1'b0;
  assign \A[7][89] [2] = 1'b0;
  assign \A[7][89] [1] = 1'b0;
  assign \A[7][89] [0] = 1'b0;
  assign \A[7][90] [4] = 1'b0;
  assign \A[7][90] [3] = 1'b0;
  assign \A[7][90] [2] = 1'b0;
  assign \A[7][90] [1] = 1'b0;
  assign \A[7][90] [0] = 1'b0;
  assign \A[7][91] [4] = 1'b0;
  assign \A[7][91] [3] = 1'b0;
  assign \A[7][91] [2] = 1'b0;
  assign \A[7][91] [1] = 1'b0;
  assign \A[7][91] [0] = 1'b0;
  assign \A[7][93] [0] = 1'b0;
  assign \A[7][94] [1] = 1'b0;
  assign \A[7][94] [0] = 1'b0;
  assign \A[7][95] [1] = 1'b0;
  assign \A[7][96] [4] = 1'b0;
  assign \A[7][96] [3] = 1'b0;
  assign \A[7][96] [2] = 1'b0;
  assign \A[7][96] [1] = 1'b0;
  assign \A[7][96] [0] = 1'b0;
  assign \A[7][98] [0] = 1'b0;
  assign \A[7][100] [4] = 1'b0;
  assign \A[7][100] [3] = 1'b0;
  assign \A[7][100] [2] = 1'b0;
  assign \A[7][100] [1] = 1'b0;
  assign \A[7][101] [4] = 1'b0;
  assign \A[7][101] [3] = 1'b0;
  assign \A[7][101] [2] = 1'b0;
  assign \A[7][101] [1] = 1'b0;
  assign \A[7][102] [4] = 1'b0;
  assign \A[7][102] [3] = 1'b0;
  assign \A[7][102] [1] = 1'b0;
  assign \A[7][104] [4] = 1'b0;
  assign \A[7][104] [3] = 1'b0;
  assign \A[7][104] [2] = 1'b0;
  assign \A[7][104] [1] = 1'b0;
  assign \A[7][105] [4] = 1'b0;
  assign \A[7][105] [3] = 1'b0;
  assign \A[7][105] [2] = 1'b0;
  assign \A[7][105] [1] = 1'b0;
  assign \A[7][105] [0] = 1'b0;
  assign \A[7][106] [4] = 1'b0;
  assign \A[7][106] [3] = 1'b0;
  assign \A[7][106] [2] = 1'b0;
  assign \A[7][106] [1] = 1'b0;
  assign \A[7][106] [0] = 1'b0;
  assign \A[7][107] [4] = 1'b0;
  assign \A[7][107] [3] = 1'b0;
  assign \A[7][107] [2] = 1'b0;
  assign \A[7][107] [0] = 1'b0;
  assign \A[7][108] [4] = 1'b0;
  assign \A[7][108] [3] = 1'b0;
  assign \A[7][108] [2] = 1'b0;
  assign \A[7][108] [1] = 1'b0;
  assign \A[7][108] [0] = 1'b0;
  assign \A[7][109] [0] = 1'b0;
  assign \A[7][110] [4] = 1'b0;
  assign \A[7][110] [3] = 1'b0;
  assign \A[7][110] [2] = 1'b0;
  assign \A[7][110] [1] = 1'b0;
  assign \A[7][110] [0] = 1'b0;
  assign \A[7][111] [2] = 1'b0;
  assign \A[7][112] [4] = 1'b0;
  assign \A[7][112] [3] = 1'b0;
  assign \A[7][112] [2] = 1'b0;
  assign \A[7][112] [1] = 1'b0;
  assign \A[7][112] [0] = 1'b0;
  assign \A[7][114] [4] = 1'b0;
  assign \A[7][114] [3] = 1'b0;
  assign \A[7][114] [2] = 1'b0;
  assign \A[7][114] [1] = 1'b0;
  assign \A[7][115] [4] = 1'b0;
  assign \A[7][115] [3] = 1'b0;
  assign \A[7][115] [2] = 1'b0;
  assign \A[7][115] [1] = 1'b0;
  assign \A[7][115] [0] = 1'b0;
  assign \A[7][116] [4] = 1'b0;
  assign \A[7][116] [3] = 1'b0;
  assign \A[7][116] [2] = 1'b0;
  assign \A[7][116] [1] = 1'b0;
  assign \A[7][116] [0] = 1'b0;
  assign \A[7][117] [4] = 1'b0;
  assign \A[7][117] [3] = 1'b0;
  assign \A[7][117] [2] = 1'b0;
  assign \A[7][117] [1] = 1'b0;
  assign \A[7][118] [4] = 1'b0;
  assign \A[7][118] [3] = 1'b0;
  assign \A[7][118] [2] = 1'b0;
  assign \A[7][118] [1] = 1'b0;
  assign \A[7][119] [4] = 1'b0;
  assign \A[7][119] [3] = 1'b0;
  assign \A[7][119] [2] = 1'b0;
  assign \A[7][119] [1] = 1'b0;
  assign \A[7][119] [0] = 1'b0;
  assign \A[7][120] [4] = 1'b0;
  assign \A[7][120] [3] = 1'b0;
  assign \A[7][120] [2] = 1'b0;
  assign \A[7][120] [1] = 1'b0;
  assign \A[7][122] [4] = 1'b0;
  assign \A[7][122] [3] = 1'b0;
  assign \A[7][122] [2] = 1'b0;
  assign \A[7][122] [1] = 1'b0;
  assign \A[7][122] [0] = 1'b0;
  assign \A[7][123] [4] = 1'b0;
  assign \A[7][123] [3] = 1'b0;
  assign \A[7][123] [2] = 1'b0;
  assign \A[7][123] [1] = 1'b0;
  assign \A[7][123] [0] = 1'b0;
  assign \A[7][124] [4] = 1'b0;
  assign \A[7][124] [3] = 1'b0;
  assign \A[7][124] [1] = 1'b0;
  assign \A[7][124] [0] = 1'b0;
  assign \A[7][125] [4] = 1'b0;
  assign \A[7][125] [3] = 1'b0;
  assign \A[7][125] [2] = 1'b0;
  assign \A[7][125] [1] = 1'b0;
  assign \A[7][125] [0] = 1'b0;
  assign \A[7][126] [0] = 1'b0;
  assign \A[7][128] [4] = 1'b0;
  assign \A[7][128] [3] = 1'b0;
  assign \A[7][128] [2] = 1'b0;
  assign \A[7][128] [0] = 1'b0;
  assign \A[7][129] [0] = 1'b0;
  assign \A[7][130] [4] = 1'b0;
  assign \A[7][130] [3] = 1'b0;
  assign \A[7][130] [2] = 1'b0;
  assign \A[7][131] [4] = 1'b0;
  assign \A[7][131] [3] = 1'b0;
  assign \A[7][131] [2] = 1'b0;
  assign \A[7][131] [1] = 1'b0;
  assign \A[7][131] [0] = 1'b0;
  assign \A[7][132] [4] = 1'b0;
  assign \A[7][132] [3] = 1'b0;
  assign \A[7][132] [2] = 1'b0;
  assign \A[7][132] [1] = 1'b0;
  assign \A[7][132] [0] = 1'b0;
  assign \A[7][133] [4] = 1'b0;
  assign \A[7][133] [3] = 1'b0;
  assign \A[7][133] [2] = 1'b0;
  assign \A[7][133] [1] = 1'b0;
  assign \A[7][134] [4] = 1'b0;
  assign \A[7][134] [3] = 1'b0;
  assign \A[7][134] [2] = 1'b0;
  assign \A[7][134] [1] = 1'b0;
  assign \A[7][135] [4] = 1'b0;
  assign \A[7][135] [3] = 1'b0;
  assign \A[7][135] [2] = 1'b0;
  assign \A[7][136] [4] = 1'b0;
  assign \A[7][136] [3] = 1'b0;
  assign \A[7][136] [2] = 1'b0;
  assign \A[7][136] [1] = 1'b0;
  assign \A[7][137] [4] = 1'b0;
  assign \A[7][137] [3] = 1'b0;
  assign \A[7][137] [2] = 1'b0;
  assign \A[7][137] [1] = 1'b0;
  assign \A[7][137] [0] = 1'b0;
  assign \A[7][138] [4] = 1'b0;
  assign \A[7][138] [3] = 1'b0;
  assign \A[7][138] [2] = 1'b0;
  assign \A[7][138] [0] = 1'b0;
  assign \A[7][139] [4] = 1'b0;
  assign \A[7][139] [3] = 1'b0;
  assign \A[7][139] [2] = 1'b0;
  assign \A[7][139] [1] = 1'b0;
  assign \A[7][139] [0] = 1'b0;
  assign \A[7][140] [4] = 1'b0;
  assign \A[7][140] [3] = 1'b0;
  assign \A[7][140] [2] = 1'b0;
  assign \A[7][140] [1] = 1'b0;
  assign \A[7][140] [0] = 1'b0;
  assign \A[7][141] [4] = 1'b0;
  assign \A[7][141] [3] = 1'b0;
  assign \A[7][141] [2] = 1'b0;
  assign \A[7][141] [1] = 1'b0;
  assign \A[7][141] [0] = 1'b0;
  assign \A[7][144] [4] = 1'b0;
  assign \A[7][144] [3] = 1'b0;
  assign \A[7][144] [2] = 1'b0;
  assign \A[7][144] [1] = 1'b0;
  assign \A[7][145] [4] = 1'b0;
  assign \A[7][145] [3] = 1'b0;
  assign \A[7][145] [2] = 1'b0;
  assign \A[7][145] [0] = 1'b0;
  assign \A[7][146] [1] = 1'b0;
  assign \A[7][147] [4] = 1'b0;
  assign \A[7][147] [3] = 1'b0;
  assign \A[7][147] [2] = 1'b0;
  assign \A[7][147] [1] = 1'b0;
  assign \A[7][147] [0] = 1'b0;
  assign \A[7][148] [4] = 1'b0;
  assign \A[7][148] [3] = 1'b0;
  assign \A[7][148] [2] = 1'b0;
  assign \A[7][148] [1] = 1'b0;
  assign \A[7][148] [0] = 1'b0;
  assign \A[7][149] [4] = 1'b0;
  assign \A[7][149] [3] = 1'b0;
  assign \A[7][149] [2] = 1'b0;
  assign \A[7][149] [1] = 1'b0;
  assign \A[7][150] [4] = 1'b0;
  assign \A[7][150] [3] = 1'b0;
  assign \A[7][150] [2] = 1'b0;
  assign \A[7][150] [1] = 1'b0;
  assign \A[7][151] [4] = 1'b0;
  assign \A[7][151] [3] = 1'b0;
  assign \A[7][151] [2] = 1'b0;
  assign \A[7][151] [1] = 1'b0;
  assign \A[7][152] [4] = 1'b0;
  assign \A[7][152] [3] = 1'b0;
  assign \A[7][152] [2] = 1'b0;
  assign \A[7][152] [1] = 1'b0;
  assign \A[7][153] [4] = 1'b0;
  assign \A[7][153] [3] = 1'b0;
  assign \A[7][153] [2] = 1'b0;
  assign \A[7][153] [1] = 1'b0;
  assign \A[7][154] [4] = 1'b0;
  assign \A[7][154] [3] = 1'b0;
  assign \A[7][154] [2] = 1'b0;
  assign \A[7][154] [0] = 1'b0;
  assign \A[7][155] [4] = 1'b0;
  assign \A[7][155] [3] = 1'b0;
  assign \A[7][155] [2] = 1'b0;
  assign \A[7][155] [1] = 1'b0;
  assign \A[7][155] [0] = 1'b0;
  assign \A[7][156] [4] = 1'b0;
  assign \A[7][156] [3] = 1'b0;
  assign \A[7][156] [2] = 1'b0;
  assign \A[7][156] [1] = 1'b0;
  assign \A[7][157] [4] = 1'b0;
  assign \A[7][157] [3] = 1'b0;
  assign \A[7][157] [2] = 1'b0;
  assign \A[7][157] [1] = 1'b0;
  assign \A[7][159] [4] = 1'b0;
  assign \A[7][159] [3] = 1'b0;
  assign \A[7][159] [2] = 1'b0;
  assign \A[7][159] [1] = 1'b0;
  assign \A[7][160] [4] = 1'b0;
  assign \A[7][160] [3] = 1'b0;
  assign \A[7][160] [2] = 1'b0;
  assign \A[7][160] [1] = 1'b0;
  assign \A[7][160] [0] = 1'b0;
  assign \A[7][161] [4] = 1'b0;
  assign \A[7][161] [3] = 1'b0;
  assign \A[7][161] [2] = 1'b0;
  assign \A[7][161] [1] = 1'b0;
  assign \A[7][162] [4] = 1'b0;
  assign \A[7][162] [3] = 1'b0;
  assign \A[7][162] [2] = 1'b0;
  assign \A[7][162] [1] = 1'b0;
  assign \A[7][163] [4] = 1'b0;
  assign \A[7][163] [3] = 1'b0;
  assign \A[7][163] [2] = 1'b0;
  assign \A[7][163] [0] = 1'b0;
  assign \A[7][164] [4] = 1'b0;
  assign \A[7][164] [3] = 1'b0;
  assign \A[7][164] [2] = 1'b0;
  assign \A[7][164] [1] = 1'b0;
  assign \A[7][164] [0] = 1'b0;
  assign \A[7][165] [4] = 1'b0;
  assign \A[7][165] [3] = 1'b0;
  assign \A[7][165] [2] = 1'b0;
  assign \A[7][165] [0] = 1'b0;
  assign \A[7][166] [4] = 1'b0;
  assign \A[7][166] [3] = 1'b0;
  assign \A[7][166] [2] = 1'b0;
  assign \A[7][166] [0] = 1'b0;
  assign \A[7][168] [4] = 1'b0;
  assign \A[7][168] [3] = 1'b0;
  assign \A[7][168] [2] = 1'b0;
  assign \A[7][168] [0] = 1'b0;
  assign \A[7][169] [4] = 1'b0;
  assign \A[7][169] [3] = 1'b0;
  assign \A[7][169] [2] = 1'b0;
  assign \A[7][169] [0] = 1'b0;
  assign \A[7][171] [4] = 1'b0;
  assign \A[7][171] [3] = 1'b0;
  assign \A[7][171] [2] = 1'b0;
  assign \A[7][171] [1] = 1'b0;
  assign \A[7][172] [4] = 1'b0;
  assign \A[7][172] [3] = 1'b0;
  assign \A[7][172] [2] = 1'b0;
  assign \A[7][172] [1] = 1'b0;
  assign \A[7][172] [0] = 1'b0;
  assign \A[7][173] [4] = 1'b0;
  assign \A[7][173] [3] = 1'b0;
  assign \A[7][173] [2] = 1'b0;
  assign \A[7][174] [4] = 1'b0;
  assign \A[7][174] [3] = 1'b0;
  assign \A[7][174] [2] = 1'b0;
  assign \A[7][174] [1] = 1'b0;
  assign \A[7][175] [4] = 1'b0;
  assign \A[7][175] [3] = 1'b0;
  assign \A[7][175] [2] = 1'b0;
  assign \A[7][175] [1] = 1'b0;
  assign \A[7][175] [0] = 1'b0;
  assign \A[7][176] [4] = 1'b0;
  assign \A[7][176] [3] = 1'b0;
  assign \A[7][176] [2] = 1'b0;
  assign \A[7][176] [1] = 1'b0;
  assign \A[7][177] [4] = 1'b0;
  assign \A[7][177] [3] = 1'b0;
  assign \A[7][177] [1] = 1'b0;
  assign \A[7][178] [4] = 1'b0;
  assign \A[7][178] [3] = 1'b0;
  assign \A[7][178] [2] = 1'b0;
  assign \A[7][178] [1] = 1'b0;
  assign \A[7][179] [4] = 1'b0;
  assign \A[7][179] [3] = 1'b0;
  assign \A[7][179] [2] = 1'b0;
  assign \A[7][179] [1] = 1'b0;
  assign \A[7][182] [4] = 1'b0;
  assign \A[7][182] [3] = 1'b0;
  assign \A[7][182] [2] = 1'b0;
  assign \A[7][182] [1] = 1'b0;
  assign \A[7][182] [0] = 1'b0;
  assign \A[7][183] [4] = 1'b0;
  assign \A[7][183] [3] = 1'b0;
  assign \A[7][183] [2] = 1'b0;
  assign \A[7][183] [1] = 1'b0;
  assign \A[7][184] [4] = 1'b0;
  assign \A[7][184] [3] = 1'b0;
  assign \A[7][184] [2] = 1'b0;
  assign \A[7][184] [1] = 1'b0;
  assign \A[7][185] [4] = 1'b0;
  assign \A[7][185] [3] = 1'b0;
  assign \A[7][185] [2] = 1'b0;
  assign \A[7][185] [1] = 1'b0;
  assign \A[7][186] [4] = 1'b0;
  assign \A[7][186] [3] = 1'b0;
  assign \A[7][186] [2] = 1'b0;
  assign \A[7][186] [1] = 1'b0;
  assign \A[7][187] [4] = 1'b0;
  assign \A[7][187] [3] = 1'b0;
  assign \A[7][187] [2] = 1'b0;
  assign \A[7][187] [1] = 1'b0;
  assign \A[7][187] [0] = 1'b0;
  assign \A[7][188] [4] = 1'b0;
  assign \A[7][188] [3] = 1'b0;
  assign \A[7][188] [2] = 1'b0;
  assign \A[7][188] [0] = 1'b0;
  assign \A[7][189] [4] = 1'b0;
  assign \A[7][189] [3] = 1'b0;
  assign \A[7][189] [2] = 1'b0;
  assign \A[7][189] [1] = 1'b0;
  assign \A[7][189] [0] = 1'b0;
  assign \A[7][190] [4] = 1'b0;
  assign \A[7][190] [3] = 1'b0;
  assign \A[7][190] [2] = 1'b0;
  assign \A[7][191] [4] = 1'b0;
  assign \A[7][191] [3] = 1'b0;
  assign \A[7][191] [2] = 1'b0;
  assign \A[7][191] [1] = 1'b0;
  assign \A[7][192] [4] = 1'b0;
  assign \A[7][192] [3] = 1'b0;
  assign \A[7][192] [2] = 1'b0;
  assign \A[7][193] [4] = 1'b0;
  assign \A[7][193] [3] = 1'b0;
  assign \A[7][193] [1] = 1'b0;
  assign \A[7][194] [4] = 1'b0;
  assign \A[7][194] [3] = 1'b0;
  assign \A[7][194] [2] = 1'b0;
  assign \A[7][194] [1] = 1'b0;
  assign \A[7][195] [4] = 1'b0;
  assign \A[7][195] [3] = 1'b0;
  assign \A[7][195] [2] = 1'b0;
  assign \A[7][195] [1] = 1'b0;
  assign \A[7][195] [0] = 1'b0;
  assign \A[7][196] [4] = 1'b0;
  assign \A[7][196] [3] = 1'b0;
  assign \A[7][196] [2] = 1'b0;
  assign \A[7][198] [0] = 1'b0;
  assign \A[7][199] [4] = 1'b0;
  assign \A[7][199] [3] = 1'b0;
  assign \A[7][199] [2] = 1'b0;
  assign \A[7][199] [1] = 1'b0;
  assign \A[7][200] [4] = 1'b0;
  assign \A[7][200] [3] = 1'b0;
  assign \A[7][200] [2] = 1'b0;
  assign \A[7][200] [1] = 1'b0;
  assign \A[7][200] [0] = 1'b0;
  assign \A[7][201] [1] = 1'b0;
  assign \A[7][202] [4] = 1'b0;
  assign \A[7][202] [3] = 1'b0;
  assign \A[7][202] [2] = 1'b0;
  assign \A[7][202] [1] = 1'b0;
  assign \A[7][203] [4] = 1'b0;
  assign \A[7][203] [3] = 1'b0;
  assign \A[7][203] [2] = 1'b0;
  assign \A[7][203] [0] = 1'b0;
  assign \A[7][204] [4] = 1'b0;
  assign \A[7][204] [3] = 1'b0;
  assign \A[7][204] [2] = 1'b0;
  assign \A[7][204] [1] = 1'b0;
  assign \A[7][204] [0] = 1'b0;
  assign \A[7][205] [4] = 1'b0;
  assign \A[7][205] [3] = 1'b0;
  assign \A[7][205] [2] = 1'b0;
  assign \A[7][205] [1] = 1'b0;
  assign \A[7][206] [4] = 1'b0;
  assign \A[7][206] [3] = 1'b0;
  assign \A[7][206] [2] = 1'b0;
  assign \A[7][206] [1] = 1'b0;
  assign \A[7][207] [4] = 1'b0;
  assign \A[7][207] [3] = 1'b0;
  assign \A[7][207] [1] = 1'b0;
  assign \A[7][207] [0] = 1'b0;
  assign \A[7][208] [4] = 1'b0;
  assign \A[7][208] [3] = 1'b0;
  assign \A[7][208] [2] = 1'b0;
  assign \A[7][208] [1] = 1'b0;
  assign \A[7][209] [4] = 1'b0;
  assign \A[7][209] [3] = 1'b0;
  assign \A[7][209] [2] = 1'b0;
  assign \A[7][209] [1] = 1'b0;
  assign \A[7][209] [0] = 1'b0;
  assign \A[7][213] [4] = 1'b0;
  assign \A[7][213] [3] = 1'b0;
  assign \A[7][213] [2] = 1'b0;
  assign \A[7][213] [1] = 1'b0;
  assign \A[7][213] [0] = 1'b0;
  assign \A[7][215] [0] = 1'b0;
  assign \A[7][216] [4] = 1'b0;
  assign \A[7][216] [3] = 1'b0;
  assign \A[7][216] [2] = 1'b0;
  assign \A[7][216] [1] = 1'b0;
  assign \A[7][217] [4] = 1'b0;
  assign \A[7][217] [3] = 1'b0;
  assign \A[7][217] [2] = 1'b0;
  assign \A[7][217] [1] = 1'b0;
  assign \A[7][217] [0] = 1'b0;
  assign \A[7][218] [1] = 1'b0;
  assign \A[7][220] [4] = 1'b0;
  assign \A[7][220] [3] = 1'b0;
  assign \A[7][220] [2] = 1'b0;
  assign \A[7][220] [1] = 1'b0;
  assign \A[7][221] [2] = 1'b0;
  assign \A[7][222] [4] = 1'b0;
  assign \A[7][222] [3] = 1'b0;
  assign \A[7][222] [2] = 1'b0;
  assign \A[7][222] [1] = 1'b0;
  assign \A[7][223] [4] = 1'b0;
  assign \A[7][223] [3] = 1'b0;
  assign \A[7][223] [2] = 1'b0;
  assign \A[7][223] [1] = 1'b0;
  assign \A[7][223] [0] = 1'b0;
  assign \A[7][224] [0] = 1'b0;
  assign \A[7][226] [0] = 1'b0;
  assign \A[7][227] [4] = 1'b0;
  assign \A[7][227] [3] = 1'b0;
  assign \A[7][227] [2] = 1'b0;
  assign \A[7][227] [0] = 1'b0;
  assign \A[7][228] [4] = 1'b0;
  assign \A[7][228] [3] = 1'b0;
  assign \A[7][228] [2] = 1'b0;
  assign \A[7][229] [4] = 1'b0;
  assign \A[7][229] [3] = 1'b0;
  assign \A[7][229] [2] = 1'b0;
  assign \A[7][229] [1] = 1'b0;
  assign \A[7][230] [4] = 1'b0;
  assign \A[7][230] [3] = 1'b0;
  assign \A[7][230] [2] = 1'b0;
  assign \A[7][230] [1] = 1'b0;
  assign \A[7][230] [0] = 1'b0;
  assign \A[7][231] [4] = 1'b0;
  assign \A[7][231] [3] = 1'b0;
  assign \A[7][231] [1] = 1'b0;
  assign \A[7][231] [0] = 1'b0;
  assign \A[7][232] [4] = 1'b0;
  assign \A[7][232] [3] = 1'b0;
  assign \A[7][232] [2] = 1'b0;
  assign \A[7][232] [1] = 1'b0;
  assign \A[7][232] [0] = 1'b0;
  assign \A[7][234] [4] = 1'b0;
  assign \A[7][234] [3] = 1'b0;
  assign \A[7][234] [2] = 1'b0;
  assign \A[7][234] [0] = 1'b0;
  assign \A[7][235] [4] = 1'b0;
  assign \A[7][235] [3] = 1'b0;
  assign \A[7][235] [2] = 1'b0;
  assign \A[7][235] [1] = 1'b0;
  assign \A[7][235] [0] = 1'b0;
  assign \A[7][236] [4] = 1'b0;
  assign \A[7][236] [3] = 1'b0;
  assign \A[7][236] [2] = 1'b0;
  assign \A[7][236] [1] = 1'b0;
  assign \A[7][236] [0] = 1'b0;
  assign \A[7][237] [4] = 1'b0;
  assign \A[7][237] [3] = 1'b0;
  assign \A[7][237] [2] = 1'b0;
  assign \A[7][237] [1] = 1'b0;
  assign \A[7][237] [0] = 1'b0;
  assign \A[7][238] [1] = 1'b0;
  assign \A[7][239] [1] = 1'b0;
  assign \A[7][240] [0] = 1'b0;
  assign \A[7][241] [4] = 1'b0;
  assign \A[7][241] [3] = 1'b0;
  assign \A[7][241] [2] = 1'b0;
  assign \A[7][241] [0] = 1'b0;
  assign \A[7][242] [4] = 1'b0;
  assign \A[7][242] [3] = 1'b0;
  assign \A[7][242] [2] = 1'b0;
  assign \A[7][242] [1] = 1'b0;
  assign \A[7][242] [0] = 1'b0;
  assign \A[7][243] [4] = 1'b0;
  assign \A[7][243] [3] = 1'b0;
  assign \A[7][243] [2] = 1'b0;
  assign \A[7][243] [0] = 1'b0;
  assign \A[7][244] [4] = 1'b0;
  assign \A[7][244] [3] = 1'b0;
  assign \A[7][244] [2] = 1'b0;
  assign \A[7][244] [1] = 1'b0;
  assign \A[7][245] [4] = 1'b0;
  assign \A[7][245] [3] = 1'b0;
  assign \A[7][245] [2] = 1'b0;
  assign \A[7][245] [1] = 1'b0;
  assign \A[7][245] [0] = 1'b0;
  assign \A[7][246] [4] = 1'b0;
  assign \A[7][246] [3] = 1'b0;
  assign \A[7][246] [2] = 1'b0;
  assign \A[7][246] [1] = 1'b0;
  assign \A[7][247] [4] = 1'b0;
  assign \A[7][247] [3] = 1'b0;
  assign \A[7][247] [2] = 1'b0;
  assign \A[7][247] [1] = 1'b0;
  assign \A[7][248] [4] = 1'b0;
  assign \A[7][248] [3] = 1'b0;
  assign \A[7][248] [2] = 1'b0;
  assign \A[7][248] [1] = 1'b0;
  assign \A[7][249] [0] = 1'b0;
  assign \A[7][250] [4] = 1'b0;
  assign \A[7][250] [3] = 1'b0;
  assign \A[7][250] [2] = 1'b0;
  assign \A[7][250] [0] = 1'b0;
  assign \A[7][251] [4] = 1'b0;
  assign \A[7][251] [3] = 1'b0;
  assign \A[7][251] [2] = 1'b0;
  assign \A[7][251] [0] = 1'b0;
  assign \A[7][252] [4] = 1'b0;
  assign \A[7][252] [3] = 1'b0;
  assign \A[7][252] [2] = 1'b0;
  assign \A[7][252] [1] = 1'b0;
  assign \A[7][252] [0] = 1'b0;
  assign \A[7][254] [1] = 1'b0;
  assign \A[7][255] [1] = 1'b0;
  assign \A[8][0] [4] = 1'b0;
  assign \A[8][0] [3] = 1'b0;
  assign \A[8][0] [2] = 1'b0;
  assign \A[8][1] [4] = 1'b0;
  assign \A[8][1] [3] = 1'b0;
  assign \A[8][1] [2] = 1'b0;
  assign \A[8][1] [1] = 1'b0;
  assign \A[8][2] [4] = 1'b0;
  assign \A[8][2] [3] = 1'b0;
  assign \A[8][2] [2] = 1'b0;
  assign \A[8][2] [0] = 1'b0;
  assign \A[8][4] [4] = 1'b0;
  assign \A[8][4] [3] = 1'b0;
  assign \A[8][4] [2] = 1'b0;
  assign \A[8][4] [1] = 1'b0;
  assign \A[8][5] [4] = 1'b0;
  assign \A[8][5] [3] = 1'b0;
  assign \A[8][5] [2] = 1'b0;
  assign \A[8][5] [1] = 1'b0;
  assign \A[8][5] [0] = 1'b0;
  assign \A[8][6] [4] = 1'b0;
  assign \A[8][6] [3] = 1'b0;
  assign \A[8][6] [2] = 1'b0;
  assign \A[8][6] [1] = 1'b0;
  assign \A[8][6] [0] = 1'b0;
  assign \A[8][7] [0] = 1'b0;
  assign \A[8][8] [4] = 1'b0;
  assign \A[8][8] [3] = 1'b0;
  assign \A[8][8] [2] = 1'b0;
  assign \A[8][8] [1] = 1'b0;
  assign \A[8][9] [4] = 1'b0;
  assign \A[8][9] [3] = 1'b0;
  assign \A[8][9] [2] = 1'b0;
  assign \A[8][9] [1] = 1'b0;
  assign \A[8][10] [0] = 1'b0;
  assign \A[8][11] [4] = 1'b0;
  assign \A[8][11] [3] = 1'b0;
  assign \A[8][11] [2] = 1'b0;
  assign \A[8][11] [1] = 1'b0;
  assign \A[8][12] [4] = 1'b0;
  assign \A[8][12] [3] = 1'b0;
  assign \A[8][12] [2] = 1'b0;
  assign \A[8][12] [1] = 1'b0;
  assign \A[8][12] [0] = 1'b0;
  assign \A[8][13] [4] = 1'b0;
  assign \A[8][13] [3] = 1'b0;
  assign \A[8][13] [2] = 1'b0;
  assign \A[8][13] [0] = 1'b0;
  assign \A[8][15] [4] = 1'b0;
  assign \A[8][15] [3] = 1'b0;
  assign \A[8][15] [2] = 1'b0;
  assign \A[8][15] [1] = 1'b0;
  assign \A[8][15] [0] = 1'b0;
  assign \A[8][17] [4] = 1'b0;
  assign \A[8][17] [3] = 1'b0;
  assign \A[8][17] [2] = 1'b0;
  assign \A[8][17] [1] = 1'b0;
  assign \A[8][17] [0] = 1'b0;
  assign \A[8][18] [4] = 1'b0;
  assign \A[8][18] [3] = 1'b0;
  assign \A[8][18] [2] = 1'b0;
  assign \A[8][18] [1] = 1'b0;
  assign \A[8][18] [0] = 1'b0;
  assign \A[8][19] [4] = 1'b0;
  assign \A[8][19] [3] = 1'b0;
  assign \A[8][19] [2] = 1'b0;
  assign \A[8][19] [0] = 1'b0;
  assign \A[8][20] [4] = 1'b0;
  assign \A[8][20] [3] = 1'b0;
  assign \A[8][20] [2] = 1'b0;
  assign \A[8][20] [0] = 1'b0;
  assign \A[8][21] [0] = 1'b0;
  assign \A[8][22] [0] = 1'b0;
  assign \A[8][24] [4] = 1'b0;
  assign \A[8][24] [3] = 1'b0;
  assign \A[8][24] [2] = 1'b0;
  assign \A[8][24] [1] = 1'b0;
  assign \A[8][26] [4] = 1'b0;
  assign \A[8][26] [3] = 1'b0;
  assign \A[8][26] [2] = 1'b0;
  assign \A[8][26] [1] = 1'b0;
  assign \A[8][26] [0] = 1'b0;
  assign \A[8][28] [4] = 1'b0;
  assign \A[8][28] [3] = 1'b0;
  assign \A[8][28] [2] = 1'b0;
  assign \A[8][28] [0] = 1'b0;
  assign \A[8][29] [0] = 1'b0;
  assign \A[8][30] [1] = 1'b0;
  assign \A[8][31] [4] = 1'b0;
  assign \A[8][31] [3] = 1'b0;
  assign \A[8][31] [2] = 1'b0;
  assign \A[8][31] [1] = 1'b0;
  assign \A[8][31] [0] = 1'b0;
  assign \A[8][32] [4] = 1'b0;
  assign \A[8][32] [3] = 1'b0;
  assign \A[8][32] [2] = 1'b0;
  assign \A[8][32] [0] = 1'b0;
  assign \A[8][33] [4] = 1'b0;
  assign \A[8][33] [3] = 1'b0;
  assign \A[8][33] [2] = 1'b0;
  assign \A[8][33] [1] = 1'b0;
  assign \A[8][33] [0] = 1'b0;
  assign \A[8][35] [4] = 1'b0;
  assign \A[8][35] [3] = 1'b0;
  assign \A[8][35] [2] = 1'b0;
  assign \A[8][35] [1] = 1'b0;
  assign \A[8][35] [0] = 1'b0;
  assign \A[8][36] [4] = 1'b0;
  assign \A[8][36] [3] = 1'b0;
  assign \A[8][36] [2] = 1'b0;
  assign \A[8][36] [1] = 1'b0;
  assign \A[8][37] [4] = 1'b0;
  assign \A[8][37] [3] = 1'b0;
  assign \A[8][37] [2] = 1'b0;
  assign \A[8][37] [1] = 1'b0;
  assign \A[8][38] [4] = 1'b0;
  assign \A[8][38] [3] = 1'b0;
  assign \A[8][38] [2] = 1'b0;
  assign \A[8][38] [1] = 1'b0;
  assign \A[8][39] [4] = 1'b0;
  assign \A[8][39] [3] = 1'b0;
  assign \A[8][39] [2] = 1'b0;
  assign \A[8][39] [1] = 1'b0;
  assign \A[8][40] [4] = 1'b0;
  assign \A[8][40] [3] = 1'b0;
  assign \A[8][40] [2] = 1'b0;
  assign \A[8][40] [1] = 1'b0;
  assign \A[8][43] [4] = 1'b0;
  assign \A[8][43] [3] = 1'b0;
  assign \A[8][43] [2] = 1'b0;
  assign \A[8][43] [1] = 1'b0;
  assign \A[8][43] [0] = 1'b0;
  assign \A[8][44] [1] = 1'b0;
  assign \A[8][45] [1] = 1'b0;
  assign \A[8][46] [4] = 1'b0;
  assign \A[8][46] [3] = 1'b0;
  assign \A[8][46] [2] = 1'b0;
  assign \A[8][46] [1] = 1'b0;
  assign \A[8][48] [4] = 1'b0;
  assign \A[8][48] [3] = 1'b0;
  assign \A[8][48] [2] = 1'b0;
  assign \A[8][49] [4] = 1'b0;
  assign \A[8][49] [3] = 1'b0;
  assign \A[8][49] [2] = 1'b0;
  assign \A[8][49] [0] = 1'b0;
  assign \A[8][50] [4] = 1'b0;
  assign \A[8][50] [3] = 1'b0;
  assign \A[8][50] [2] = 1'b0;
  assign \A[8][50] [1] = 1'b0;
  assign \A[8][50] [0] = 1'b0;
  assign \A[8][51] [4] = 1'b0;
  assign \A[8][51] [3] = 1'b0;
  assign \A[8][51] [2] = 1'b0;
  assign \A[8][51] [0] = 1'b0;
  assign \A[8][52] [4] = 1'b0;
  assign \A[8][52] [3] = 1'b0;
  assign \A[8][52] [2] = 1'b0;
  assign \A[8][52] [1] = 1'b0;
  assign \A[8][52] [0] = 1'b0;
  assign \A[8][53] [4] = 1'b0;
  assign \A[8][53] [3] = 1'b0;
  assign \A[8][53] [2] = 1'b0;
  assign \A[8][53] [0] = 1'b0;
  assign \A[8][54] [4] = 1'b0;
  assign \A[8][54] [3] = 1'b0;
  assign \A[8][54] [2] = 1'b0;
  assign \A[8][54] [1] = 1'b0;
  assign \A[8][55] [1] = 1'b0;
  assign \A[8][57] [0] = 1'b0;
  assign \A[8][59] [0] = 1'b0;
  assign \A[8][60] [4] = 1'b0;
  assign \A[8][60] [3] = 1'b0;
  assign \A[8][60] [2] = 1'b0;
  assign \A[8][60] [1] = 1'b0;
  assign \A[8][60] [0] = 1'b0;
  assign \A[8][62] [0] = 1'b0;
  assign \A[8][63] [0] = 1'b0;
  assign \A[8][64] [1] = 1'b0;
  assign \A[8][65] [4] = 1'b0;
  assign \A[8][65] [3] = 1'b0;
  assign \A[8][65] [2] = 1'b0;
  assign \A[8][66] [4] = 1'b0;
  assign \A[8][66] [3] = 1'b0;
  assign \A[8][66] [2] = 1'b0;
  assign \A[8][66] [1] = 1'b0;
  assign \A[8][66] [0] = 1'b0;
  assign \A[8][68] [4] = 1'b0;
  assign \A[8][68] [3] = 1'b0;
  assign \A[8][68] [2] = 1'b0;
  assign \A[8][68] [1] = 1'b0;
  assign \A[8][69] [4] = 1'b0;
  assign \A[8][69] [3] = 1'b0;
  assign \A[8][69] [2] = 1'b0;
  assign \A[8][69] [1] = 1'b0;
  assign \A[8][70] [4] = 1'b0;
  assign \A[8][70] [3] = 1'b0;
  assign \A[8][70] [2] = 1'b0;
  assign \A[8][70] [1] = 1'b0;
  assign \A[8][70] [0] = 1'b0;
  assign \A[8][71] [1] = 1'b0;
  assign \A[8][72] [1] = 1'b0;
  assign \A[8][72] [0] = 1'b0;
  assign \A[8][73] [1] = 1'b0;
  assign \A[8][73] [0] = 1'b0;
  assign \A[8][74] [4] = 1'b0;
  assign \A[8][74] [3] = 1'b0;
  assign \A[8][74] [2] = 1'b0;
  assign \A[8][74] [1] = 1'b0;
  assign \A[8][74] [0] = 1'b0;
  assign \A[8][76] [1] = 1'b0;
  assign \A[8][77] [0] = 1'b0;
  assign \A[8][78] [0] = 1'b0;
  assign \A[8][79] [4] = 1'b0;
  assign \A[8][79] [3] = 1'b0;
  assign \A[8][79] [2] = 1'b0;
  assign \A[8][79] [1] = 1'b0;
  assign \A[8][80] [0] = 1'b0;
  assign \A[8][81] [0] = 1'b0;
  assign \A[8][82] [0] = 1'b0;
  assign \A[8][83] [0] = 1'b0;
  assign \A[8][84] [1] = 1'b0;
  assign \A[8][85] [4] = 1'b0;
  assign \A[8][85] [3] = 1'b0;
  assign \A[8][85] [2] = 1'b0;
  assign \A[8][85] [1] = 1'b0;
  assign \A[8][85] [0] = 1'b0;
  assign \A[8][86] [0] = 1'b0;
  assign \A[8][87] [4] = 1'b0;
  assign \A[8][87] [3] = 1'b0;
  assign \A[8][87] [2] = 1'b0;
  assign \A[8][87] [1] = 1'b0;
  assign \A[8][87] [0] = 1'b0;
  assign \A[8][88] [4] = 1'b0;
  assign \A[8][88] [3] = 1'b0;
  assign \A[8][88] [2] = 1'b0;
  assign \A[8][88] [1] = 1'b0;
  assign \A[8][90] [4] = 1'b0;
  assign \A[8][90] [3] = 1'b0;
  assign \A[8][90] [2] = 1'b0;
  assign \A[8][90] [1] = 1'b0;
  assign \A[8][91] [1] = 1'b0;
  assign \A[8][92] [0] = 1'b0;
  assign \A[8][93] [4] = 1'b0;
  assign \A[8][93] [3] = 1'b0;
  assign \A[8][93] [2] = 1'b0;
  assign \A[8][93] [0] = 1'b0;
  assign \A[8][94] [2] = 1'b0;
  assign \A[8][95] [4] = 1'b0;
  assign \A[8][95] [3] = 1'b0;
  assign \A[8][95] [2] = 1'b0;
  assign \A[8][95] [1] = 1'b0;
  assign \A[8][96] [0] = 1'b0;
  assign \A[8][97] [0] = 1'b0;
  assign \A[8][99] [4] = 1'b0;
  assign \A[8][99] [3] = 1'b0;
  assign \A[8][99] [2] = 1'b0;
  assign \A[8][99] [1] = 1'b0;
  assign \A[8][99] [0] = 1'b0;
  assign \A[8][100] [1] = 1'b0;
  assign \A[8][101] [4] = 1'b0;
  assign \A[8][101] [3] = 1'b0;
  assign \A[8][101] [2] = 1'b0;
  assign \A[8][101] [1] = 1'b0;
  assign \A[8][101] [0] = 1'b0;
  assign \A[8][102] [4] = 1'b0;
  assign \A[8][102] [3] = 1'b0;
  assign \A[8][102] [2] = 1'b0;
  assign \A[8][102] [1] = 1'b0;
  assign \A[8][102] [0] = 1'b0;
  assign \A[8][104] [0] = 1'b0;
  assign \A[8][107] [4] = 1'b0;
  assign \A[8][107] [3] = 1'b0;
  assign \A[8][107] [2] = 1'b0;
  assign \A[8][107] [1] = 1'b0;
  assign \A[8][107] [0] = 1'b0;
  assign \A[8][108] [4] = 1'b0;
  assign \A[8][108] [3] = 1'b0;
  assign \A[8][108] [2] = 1'b0;
  assign \A[8][108] [1] = 1'b0;
  assign \A[8][108] [0] = 1'b0;
  assign \A[8][109] [4] = 1'b0;
  assign \A[8][109] [3] = 1'b0;
  assign \A[8][109] [2] = 1'b0;
  assign \A[8][109] [1] = 1'b0;
  assign \A[8][111] [1] = 1'b0;
  assign \A[8][112] [4] = 1'b0;
  assign \A[8][112] [3] = 1'b0;
  assign \A[8][112] [2] = 1'b0;
  assign \A[8][112] [1] = 1'b0;
  assign \A[8][113] [0] = 1'b0;
  assign \A[8][114] [0] = 1'b0;
  assign \A[8][115] [4] = 1'b0;
  assign \A[8][115] [3] = 1'b0;
  assign \A[8][115] [2] = 1'b0;
  assign \A[8][115] [1] = 1'b0;
  assign \A[8][116] [4] = 1'b0;
  assign \A[8][116] [3] = 1'b0;
  assign \A[8][116] [2] = 1'b0;
  assign \A[8][116] [1] = 1'b0;
  assign \A[8][116] [0] = 1'b0;
  assign \A[8][117] [4] = 1'b0;
  assign \A[8][117] [3] = 1'b0;
  assign \A[8][117] [2] = 1'b0;
  assign \A[8][117] [1] = 1'b0;
  assign \A[8][118] [0] = 1'b0;
  assign \A[8][119] [4] = 1'b0;
  assign \A[8][119] [3] = 1'b0;
  assign \A[8][119] [2] = 1'b0;
  assign \A[8][119] [1] = 1'b0;
  assign \A[8][120] [0] = 1'b0;
  assign \A[8][122] [4] = 1'b0;
  assign \A[8][122] [3] = 1'b0;
  assign \A[8][122] [2] = 1'b0;
  assign \A[8][122] [1] = 1'b0;
  assign \A[8][123] [4] = 1'b0;
  assign \A[8][123] [3] = 1'b0;
  assign \A[8][123] [2] = 1'b0;
  assign \A[8][123] [1] = 1'b0;
  assign \A[8][123] [0] = 1'b0;
  assign \A[8][124] [4] = 1'b0;
  assign \A[8][124] [3] = 1'b0;
  assign \A[8][124] [2] = 1'b0;
  assign \A[8][124] [1] = 1'b0;
  assign \A[8][125] [0] = 1'b0;
  assign \A[8][127] [4] = 1'b0;
  assign \A[8][127] [3] = 1'b0;
  assign \A[8][127] [2] = 1'b0;
  assign \A[8][127] [1] = 1'b0;
  assign \A[8][127] [0] = 1'b0;
  assign \A[8][128] [4] = 1'b0;
  assign \A[8][128] [3] = 1'b0;
  assign \A[8][128] [2] = 1'b0;
  assign \A[8][128] [0] = 1'b0;
  assign \A[8][129] [4] = 1'b0;
  assign \A[8][129] [3] = 1'b0;
  assign \A[8][129] [2] = 1'b0;
  assign \A[8][129] [1] = 1'b0;
  assign \A[8][130] [4] = 1'b0;
  assign \A[8][130] [3] = 1'b0;
  assign \A[8][130] [2] = 1'b0;
  assign \A[8][130] [1] = 1'b0;
  assign \A[8][131] [4] = 1'b0;
  assign \A[8][131] [3] = 1'b0;
  assign \A[8][131] [2] = 1'b0;
  assign \A[8][132] [0] = 1'b0;
  assign \A[8][133] [4] = 1'b0;
  assign \A[8][133] [3] = 1'b0;
  assign \A[8][133] [2] = 1'b0;
  assign \A[8][133] [1] = 1'b0;
  assign \A[8][133] [0] = 1'b0;
  assign \A[8][134] [4] = 1'b0;
  assign \A[8][134] [3] = 1'b0;
  assign \A[8][134] [2] = 1'b0;
  assign \A[8][134] [1] = 1'b0;
  assign \A[8][135] [4] = 1'b0;
  assign \A[8][135] [3] = 1'b0;
  assign \A[8][135] [2] = 1'b0;
  assign \A[8][135] [1] = 1'b0;
  assign \A[8][135] [0] = 1'b0;
  assign \A[8][136] [4] = 1'b0;
  assign \A[8][136] [3] = 1'b0;
  assign \A[8][136] [2] = 1'b0;
  assign \A[8][136] [1] = 1'b0;
  assign \A[8][137] [1] = 1'b0;
  assign \A[8][138] [4] = 1'b0;
  assign \A[8][138] [3] = 1'b0;
  assign \A[8][138] [2] = 1'b0;
  assign \A[8][138] [1] = 1'b0;
  assign \A[8][140] [0] = 1'b0;
  assign \A[8][141] [4] = 1'b0;
  assign \A[8][141] [3] = 1'b0;
  assign \A[8][141] [2] = 1'b0;
  assign \A[8][141] [1] = 1'b0;
  assign \A[8][142] [0] = 1'b0;
  assign \A[8][143] [4] = 1'b0;
  assign \A[8][143] [3] = 1'b0;
  assign \A[8][143] [2] = 1'b0;
  assign \A[8][143] [0] = 1'b0;
  assign \A[8][144] [4] = 1'b0;
  assign \A[8][144] [3] = 1'b0;
  assign \A[8][144] [2] = 1'b0;
  assign \A[8][144] [1] = 1'b0;
  assign \A[8][145] [4] = 1'b0;
  assign \A[8][145] [3] = 1'b0;
  assign \A[8][145] [2] = 1'b0;
  assign \A[8][145] [0] = 1'b0;
  assign \A[8][146] [4] = 1'b0;
  assign \A[8][146] [3] = 1'b0;
  assign \A[8][146] [2] = 1'b0;
  assign \A[8][146] [1] = 1'b0;
  assign \A[8][147] [4] = 1'b0;
  assign \A[8][147] [3] = 1'b0;
  assign \A[8][147] [2] = 1'b0;
  assign \A[8][147] [0] = 1'b0;
  assign \A[8][148] [4] = 1'b0;
  assign \A[8][148] [3] = 1'b0;
  assign \A[8][148] [2] = 1'b0;
  assign \A[8][149] [4] = 1'b0;
  assign \A[8][149] [3] = 1'b0;
  assign \A[8][149] [2] = 1'b0;
  assign \A[8][149] [1] = 1'b0;
  assign \A[8][150] [0] = 1'b0;
  assign \A[8][152] [4] = 1'b0;
  assign \A[8][152] [3] = 1'b0;
  assign \A[8][152] [2] = 1'b0;
  assign \A[8][152] [0] = 1'b0;
  assign \A[8][153] [4] = 1'b0;
  assign \A[8][153] [3] = 1'b0;
  assign \A[8][153] [2] = 1'b0;
  assign \A[8][153] [1] = 1'b0;
  assign \A[8][153] [0] = 1'b0;
  assign \A[8][154] [4] = 1'b0;
  assign \A[8][154] [3] = 1'b0;
  assign \A[8][154] [2] = 1'b0;
  assign \A[8][154] [0] = 1'b0;
  assign \A[8][155] [4] = 1'b0;
  assign \A[8][155] [3] = 1'b0;
  assign \A[8][155] [2] = 1'b0;
  assign \A[8][155] [1] = 1'b0;
  assign \A[8][155] [0] = 1'b0;
  assign \A[8][156] [4] = 1'b0;
  assign \A[8][156] [3] = 1'b0;
  assign \A[8][156] [2] = 1'b0;
  assign \A[8][156] [1] = 1'b0;
  assign \A[8][157] [4] = 1'b0;
  assign \A[8][157] [3] = 1'b0;
  assign \A[8][157] [2] = 1'b0;
  assign \A[8][157] [1] = 1'b0;
  assign \A[8][158] [1] = 1'b0;
  assign \A[8][158] [0] = 1'b0;
  assign \A[8][160] [4] = 1'b0;
  assign \A[8][160] [3] = 1'b0;
  assign \A[8][160] [2] = 1'b0;
  assign \A[8][160] [0] = 1'b0;
  assign \A[8][161] [4] = 1'b0;
  assign \A[8][161] [3] = 1'b0;
  assign \A[8][161] [1] = 1'b0;
  assign \A[8][161] [0] = 1'b0;
  assign \A[8][162] [4] = 1'b0;
  assign \A[8][162] [3] = 1'b0;
  assign \A[8][162] [2] = 1'b0;
  assign \A[8][163] [4] = 1'b0;
  assign \A[8][163] [3] = 1'b0;
  assign \A[8][163] [2] = 1'b0;
  assign \A[8][163] [1] = 1'b0;
  assign \A[8][164] [4] = 1'b0;
  assign \A[8][164] [3] = 1'b0;
  assign \A[8][164] [2] = 1'b0;
  assign \A[8][165] [4] = 1'b0;
  assign \A[8][165] [3] = 1'b0;
  assign \A[8][165] [2] = 1'b0;
  assign \A[8][165] [1] = 1'b0;
  assign \A[8][166] [4] = 1'b0;
  assign \A[8][166] [3] = 1'b0;
  assign \A[8][166] [1] = 1'b0;
  assign \A[8][166] [0] = 1'b0;
  assign \A[8][167] [4] = 1'b0;
  assign \A[8][167] [3] = 1'b0;
  assign \A[8][167] [2] = 1'b0;
  assign \A[8][167] [1] = 1'b0;
  assign \A[8][167] [0] = 1'b0;
  assign \A[8][168] [4] = 1'b0;
  assign \A[8][168] [3] = 1'b0;
  assign \A[8][168] [2] = 1'b0;
  assign \A[8][168] [1] = 1'b0;
  assign \A[8][169] [4] = 1'b0;
  assign \A[8][169] [3] = 1'b0;
  assign \A[8][169] [2] = 1'b0;
  assign \A[8][169] [0] = 1'b0;
  assign \A[8][173] [0] = 1'b0;
  assign \A[8][174] [4] = 1'b0;
  assign \A[8][174] [3] = 1'b0;
  assign \A[8][174] [2] = 1'b0;
  assign \A[8][174] [1] = 1'b0;
  assign \A[8][174] [0] = 1'b0;
  assign \A[8][175] [4] = 1'b0;
  assign \A[8][175] [3] = 1'b0;
  assign \A[8][175] [2] = 1'b0;
  assign \A[8][175] [1] = 1'b0;
  assign \A[8][177] [4] = 1'b0;
  assign \A[8][177] [3] = 1'b0;
  assign \A[8][177] [1] = 1'b0;
  assign \A[8][177] [0] = 1'b0;
  assign \A[8][178] [4] = 1'b0;
  assign \A[8][178] [3] = 1'b0;
  assign \A[8][178] [2] = 1'b0;
  assign \A[8][178] [1] = 1'b0;
  assign \A[8][179] [4] = 1'b0;
  assign \A[8][179] [3] = 1'b0;
  assign \A[8][179] [2] = 1'b0;
  assign \A[8][179] [0] = 1'b0;
  assign \A[8][180] [4] = 1'b0;
  assign \A[8][180] [3] = 1'b0;
  assign \A[8][180] [2] = 1'b0;
  assign \A[8][181] [4] = 1'b0;
  assign \A[8][181] [3] = 1'b0;
  assign \A[8][181] [2] = 1'b0;
  assign \A[8][182] [4] = 1'b0;
  assign \A[8][182] [3] = 1'b0;
  assign \A[8][182] [2] = 1'b0;
  assign \A[8][183] [4] = 1'b0;
  assign \A[8][183] [3] = 1'b0;
  assign \A[8][183] [2] = 1'b0;
  assign \A[8][183] [1] = 1'b0;
  assign \A[8][183] [0] = 1'b0;
  assign \A[8][184] [0] = 1'b0;
  assign \A[8][185] [4] = 1'b0;
  assign \A[8][185] [3] = 1'b0;
  assign \A[8][185] [2] = 1'b0;
  assign \A[8][185] [1] = 1'b0;
  assign \A[8][185] [0] = 1'b0;
  assign \A[8][187] [0] = 1'b0;
  assign \A[8][188] [1] = 1'b0;
  assign \A[8][188] [0] = 1'b0;
  assign \A[8][189] [4] = 1'b0;
  assign \A[8][189] [3] = 1'b0;
  assign \A[8][189] [2] = 1'b0;
  assign \A[8][189] [1] = 1'b0;
  assign \A[8][189] [0] = 1'b0;
  assign \A[8][190] [0] = 1'b0;
  assign \A[8][191] [1] = 1'b0;
  assign \A[8][192] [4] = 1'b0;
  assign \A[8][192] [3] = 1'b0;
  assign \A[8][192] [2] = 1'b0;
  assign \A[8][192] [1] = 1'b0;
  assign \A[8][193] [4] = 1'b0;
  assign \A[8][193] [3] = 1'b0;
  assign \A[8][193] [1] = 1'b0;
  assign \A[8][193] [0] = 1'b0;
  assign \A[8][194] [4] = 1'b0;
  assign \A[8][194] [3] = 1'b0;
  assign \A[8][194] [2] = 1'b0;
  assign \A[8][194] [1] = 1'b0;
  assign \A[8][194] [0] = 1'b0;
  assign \A[8][195] [4] = 1'b0;
  assign \A[8][195] [3] = 1'b0;
  assign \A[8][195] [2] = 1'b0;
  assign \A[8][196] [4] = 1'b0;
  assign \A[8][196] [3] = 1'b0;
  assign \A[8][196] [2] = 1'b0;
  assign \A[8][196] [1] = 1'b0;
  assign \A[8][197] [4] = 1'b0;
  assign \A[8][197] [3] = 1'b0;
  assign \A[8][197] [2] = 1'b0;
  assign \A[8][197] [1] = 1'b0;
  assign \A[8][198] [4] = 1'b0;
  assign \A[8][198] [3] = 1'b0;
  assign \A[8][198] [2] = 1'b0;
  assign \A[8][200] [4] = 1'b0;
  assign \A[8][200] [3] = 1'b0;
  assign \A[8][200] [2] = 1'b0;
  assign \A[8][200] [0] = 1'b0;
  assign \A[8][201] [4] = 1'b0;
  assign \A[8][201] [3] = 1'b0;
  assign \A[8][201] [2] = 1'b0;
  assign \A[8][201] [1] = 1'b0;
  assign \A[8][202] [4] = 1'b0;
  assign \A[8][202] [3] = 1'b0;
  assign \A[8][202] [2] = 1'b0;
  assign \A[8][202] [1] = 1'b0;
  assign \A[8][202] [0] = 1'b0;
  assign \A[8][204] [4] = 1'b0;
  assign \A[8][204] [3] = 1'b0;
  assign \A[8][204] [2] = 1'b0;
  assign \A[8][204] [0] = 1'b0;
  assign \A[8][205] [0] = 1'b0;
  assign \A[8][207] [4] = 1'b0;
  assign \A[8][207] [3] = 1'b0;
  assign \A[8][207] [2] = 1'b0;
  assign \A[8][207] [1] = 1'b0;
  assign \A[8][208] [4] = 1'b0;
  assign \A[8][208] [3] = 1'b0;
  assign \A[8][208] [1] = 1'b0;
  assign \A[8][208] [0] = 1'b0;
  assign \A[8][209] [4] = 1'b0;
  assign \A[8][209] [3] = 1'b0;
  assign \A[8][209] [2] = 1'b0;
  assign \A[8][209] [1] = 1'b0;
  assign \A[8][211] [4] = 1'b0;
  assign \A[8][211] [3] = 1'b0;
  assign \A[8][211] [2] = 1'b0;
  assign \A[8][211] [1] = 1'b0;
  assign \A[8][212] [4] = 1'b0;
  assign \A[8][212] [3] = 1'b0;
  assign \A[8][212] [2] = 1'b0;
  assign \A[8][212] [1] = 1'b0;
  assign \A[8][212] [0] = 1'b0;
  assign \A[8][213] [4] = 1'b0;
  assign \A[8][213] [3] = 1'b0;
  assign \A[8][213] [2] = 1'b0;
  assign \A[8][213] [1] = 1'b0;
  assign \A[8][213] [0] = 1'b0;
  assign \A[8][214] [4] = 1'b0;
  assign \A[8][214] [3] = 1'b0;
  assign \A[8][214] [2] = 1'b0;
  assign \A[8][214] [1] = 1'b0;
  assign \A[8][214] [0] = 1'b0;
  assign \A[8][216] [4] = 1'b0;
  assign \A[8][216] [3] = 1'b0;
  assign \A[8][216] [2] = 1'b0;
  assign \A[8][216] [1] = 1'b0;
  assign \A[8][217] [4] = 1'b0;
  assign \A[8][217] [3] = 1'b0;
  assign \A[8][217] [2] = 1'b0;
  assign \A[8][217] [1] = 1'b0;
  assign \A[8][217] [0] = 1'b0;
  assign \A[8][218] [4] = 1'b0;
  assign \A[8][218] [3] = 1'b0;
  assign \A[8][218] [2] = 1'b0;
  assign \A[8][218] [1] = 1'b0;
  assign \A[8][219] [4] = 1'b0;
  assign \A[8][219] [3] = 1'b0;
  assign \A[8][219] [2] = 1'b0;
  assign \A[8][219] [1] = 1'b0;
  assign \A[8][219] [0] = 1'b0;
  assign \A[8][223] [1] = 1'b0;
  assign \A[8][224] [4] = 1'b0;
  assign \A[8][224] [3] = 1'b0;
  assign \A[8][224] [2] = 1'b0;
  assign \A[8][224] [1] = 1'b0;
  assign \A[8][226] [4] = 1'b0;
  assign \A[8][226] [3] = 1'b0;
  assign \A[8][226] [2] = 1'b0;
  assign \A[8][226] [1] = 1'b0;
  assign \A[8][227] [4] = 1'b0;
  assign \A[8][227] [3] = 1'b0;
  assign \A[8][227] [2] = 1'b0;
  assign \A[8][227] [1] = 1'b0;
  assign \A[8][229] [4] = 1'b0;
  assign \A[8][229] [3] = 1'b0;
  assign \A[8][229] [2] = 1'b0;
  assign \A[8][229] [1] = 1'b0;
  assign \A[8][230] [4] = 1'b0;
  assign \A[8][230] [3] = 1'b0;
  assign \A[8][230] [2] = 1'b0;
  assign \A[8][231] [0] = 1'b0;
  assign \A[8][233] [4] = 1'b0;
  assign \A[8][233] [3] = 1'b0;
  assign \A[8][233] [2] = 1'b0;
  assign \A[8][233] [1] = 1'b0;
  assign \A[8][234] [4] = 1'b0;
  assign \A[8][234] [3] = 1'b0;
  assign \A[8][234] [2] = 1'b0;
  assign \A[8][234] [1] = 1'b0;
  assign \A[8][235] [0] = 1'b0;
  assign \A[8][236] [4] = 1'b0;
  assign \A[8][236] [3] = 1'b0;
  assign \A[8][236] [2] = 1'b0;
  assign \A[8][236] [1] = 1'b0;
  assign \A[8][238] [0] = 1'b0;
  assign \A[8][239] [4] = 1'b0;
  assign \A[8][239] [3] = 1'b0;
  assign \A[8][239] [2] = 1'b0;
  assign \A[8][239] [0] = 1'b0;
  assign \A[8][240] [1] = 1'b0;
  assign \A[8][241] [4] = 1'b0;
  assign \A[8][241] [3] = 1'b0;
  assign \A[8][241] [2] = 1'b0;
  assign \A[8][241] [1] = 1'b0;
  assign \A[8][242] [4] = 1'b0;
  assign \A[8][242] [3] = 1'b0;
  assign \A[8][242] [2] = 1'b0;
  assign \A[8][242] [1] = 1'b0;
  assign \A[8][242] [0] = 1'b0;
  assign \A[8][243] [0] = 1'b0;
  assign \A[8][244] [4] = 1'b0;
  assign \A[8][244] [3] = 1'b0;
  assign \A[8][244] [2] = 1'b0;
  assign \A[8][244] [1] = 1'b0;
  assign \A[8][244] [0] = 1'b0;
  assign \A[8][245] [4] = 1'b0;
  assign \A[8][245] [3] = 1'b0;
  assign \A[8][245] [2] = 1'b0;
  assign \A[8][245] [1] = 1'b0;
  assign \A[8][245] [0] = 1'b0;
  assign \A[8][246] [4] = 1'b0;
  assign \A[8][246] [3] = 1'b0;
  assign \A[8][246] [2] = 1'b0;
  assign \A[8][246] [1] = 1'b0;
  assign \A[8][246] [0] = 1'b0;
  assign \A[8][247] [4] = 1'b0;
  assign \A[8][247] [3] = 1'b0;
  assign \A[8][247] [2] = 1'b0;
  assign \A[8][247] [0] = 1'b0;
  assign \A[8][248] [4] = 1'b0;
  assign \A[8][248] [3] = 1'b0;
  assign \A[8][248] [2] = 1'b0;
  assign \A[8][248] [1] = 1'b0;
  assign \A[8][248] [0] = 1'b0;
  assign \A[8][249] [4] = 1'b0;
  assign \A[8][249] [3] = 1'b0;
  assign \A[8][249] [2] = 1'b0;
  assign \A[8][249] [1] = 1'b0;
  assign \A[8][249] [0] = 1'b0;
  assign \A[8][250] [4] = 1'b0;
  assign \A[8][250] [3] = 1'b0;
  assign \A[8][250] [2] = 1'b0;
  assign \A[8][250] [0] = 1'b0;
  assign \A[8][251] [4] = 1'b0;
  assign \A[8][251] [3] = 1'b0;
  assign \A[8][251] [2] = 1'b0;
  assign \A[8][251] [1] = 1'b0;
  assign \A[8][253] [4] = 1'b0;
  assign \A[8][253] [3] = 1'b0;
  assign \A[8][253] [1] = 1'b0;
  assign \A[8][253] [0] = 1'b0;
  assign \A[8][254] [4] = 1'b0;
  assign \A[8][254] [3] = 1'b0;
  assign \A[8][254] [2] = 1'b0;
  assign \A[8][254] [1] = 1'b0;
  assign \A[8][254] [0] = 1'b0;
  assign \A[8][255] [4] = 1'b0;
  assign \A[8][255] [3] = 1'b0;
  assign \A[8][255] [2] = 1'b0;
  assign \A[8][255] [1] = 1'b0;
  assign \A[8][255] [0] = 1'b0;
  assign \A[9][0] [4] = 1'b0;
  assign \A[9][0] [3] = 1'b0;
  assign \A[9][0] [1] = 1'b0;
  assign \A[9][0] [0] = 1'b0;
  assign \A[9][1] [4] = 1'b0;
  assign \A[9][1] [3] = 1'b0;
  assign \A[9][1] [2] = 1'b0;
  assign \A[9][1] [1] = 1'b0;
  assign \A[9][1] [0] = 1'b0;
  assign \A[9][2] [4] = 1'b0;
  assign \A[9][2] [3] = 1'b0;
  assign \A[9][2] [2] = 1'b0;
  assign \A[9][2] [0] = 1'b0;
  assign \A[9][3] [4] = 1'b0;
  assign \A[9][3] [3] = 1'b0;
  assign \A[9][3] [2] = 1'b0;
  assign \A[9][5] [4] = 1'b0;
  assign \A[9][5] [3] = 1'b0;
  assign \A[9][5] [2] = 1'b0;
  assign \A[9][5] [0] = 1'b0;
  assign \A[9][6] [0] = 1'b0;
  assign \A[9][7] [4] = 1'b0;
  assign \A[9][7] [3] = 1'b0;
  assign \A[9][7] [1] = 1'b0;
  assign \A[9][8] [4] = 1'b0;
  assign \A[9][8] [3] = 1'b0;
  assign \A[9][8] [2] = 1'b0;
  assign \A[9][8] [1] = 1'b0;
  assign \A[9][9] [4] = 1'b0;
  assign \A[9][9] [3] = 1'b0;
  assign \A[9][9] [2] = 1'b0;
  assign \A[9][9] [1] = 1'b0;
  assign \A[9][9] [0] = 1'b0;
  assign \A[9][10] [4] = 1'b0;
  assign \A[9][10] [3] = 1'b0;
  assign \A[9][10] [2] = 1'b0;
  assign \A[9][10] [1] = 1'b0;
  assign \A[9][12] [4] = 1'b0;
  assign \A[9][12] [3] = 1'b0;
  assign \A[9][12] [2] = 1'b0;
  assign \A[9][12] [1] = 1'b0;
  assign \A[9][12] [0] = 1'b0;
  assign \A[9][13] [4] = 1'b0;
  assign \A[9][13] [3] = 1'b0;
  assign \A[9][13] [2] = 1'b0;
  assign \A[9][13] [1] = 1'b0;
  assign \A[9][13] [0] = 1'b0;
  assign \A[9][15] [4] = 1'b0;
  assign \A[9][15] [3] = 1'b0;
  assign \A[9][15] [2] = 1'b0;
  assign \A[9][15] [1] = 1'b0;
  assign \A[9][15] [0] = 1'b0;
  assign \A[9][16] [4] = 1'b0;
  assign \A[9][16] [3] = 1'b0;
  assign \A[9][16] [2] = 1'b0;
  assign \A[9][16] [0] = 1'b0;
  assign \A[9][17] [4] = 1'b0;
  assign \A[9][17] [3] = 1'b0;
  assign \A[9][17] [2] = 1'b0;
  assign \A[9][17] [0] = 1'b0;
  assign \A[9][18] [0] = 1'b0;
  assign \A[9][19] [4] = 1'b0;
  assign \A[9][19] [3] = 1'b0;
  assign \A[9][19] [2] = 1'b0;
  assign \A[9][19] [0] = 1'b0;
  assign \A[9][20] [4] = 1'b0;
  assign \A[9][20] [3] = 1'b0;
  assign \A[9][20] [2] = 1'b0;
  assign \A[9][20] [1] = 1'b0;
  assign \A[9][20] [0] = 1'b0;
  assign \A[9][21] [4] = 1'b0;
  assign \A[9][21] [3] = 1'b0;
  assign \A[9][21] [2] = 1'b0;
  assign \A[9][21] [1] = 1'b0;
  assign \A[9][22] [4] = 1'b0;
  assign \A[9][22] [3] = 1'b0;
  assign \A[9][22] [2] = 1'b0;
  assign \A[9][22] [1] = 1'b0;
  assign \A[9][23] [4] = 1'b0;
  assign \A[9][23] [3] = 1'b0;
  assign \A[9][23] [2] = 1'b0;
  assign \A[9][23] [1] = 1'b0;
  assign \A[9][23] [0] = 1'b0;
  assign \A[9][24] [4] = 1'b0;
  assign \A[9][24] [3] = 1'b0;
  assign \A[9][24] [2] = 1'b0;
  assign \A[9][24] [1] = 1'b0;
  assign \A[9][24] [0] = 1'b0;
  assign \A[9][25] [0] = 1'b0;
  assign \A[9][27] [4] = 1'b0;
  assign \A[9][27] [3] = 1'b0;
  assign \A[9][27] [2] = 1'b0;
  assign \A[9][27] [1] = 1'b0;
  assign \A[9][27] [0] = 1'b0;
  assign \A[9][28] [4] = 1'b0;
  assign \A[9][28] [3] = 1'b0;
  assign \A[9][28] [2] = 1'b0;
  assign \A[9][28] [1] = 1'b0;
  assign \A[9][28] [0] = 1'b0;
  assign \A[9][29] [0] = 1'b0;
  assign \A[9][30] [4] = 1'b0;
  assign \A[9][30] [3] = 1'b0;
  assign \A[9][30] [1] = 1'b0;
  assign \A[9][30] [0] = 1'b0;
  assign \A[9][31] [4] = 1'b0;
  assign \A[9][31] [3] = 1'b0;
  assign \A[9][31] [2] = 1'b0;
  assign \A[9][31] [1] = 1'b0;
  assign \A[9][31] [0] = 1'b0;
  assign \A[9][33] [4] = 1'b0;
  assign \A[9][33] [3] = 1'b0;
  assign \A[9][33] [2] = 1'b0;
  assign \A[9][33] [0] = 1'b0;
  assign \A[9][34] [4] = 1'b0;
  assign \A[9][34] [3] = 1'b0;
  assign \A[9][34] [2] = 1'b0;
  assign \A[9][34] [1] = 1'b0;
  assign \A[9][35] [4] = 1'b0;
  assign \A[9][35] [3] = 1'b0;
  assign \A[9][35] [2] = 1'b0;
  assign \A[9][35] [1] = 1'b0;
  assign \A[9][35] [0] = 1'b0;
  assign \A[9][36] [4] = 1'b0;
  assign \A[9][36] [3] = 1'b0;
  assign \A[9][36] [2] = 1'b0;
  assign \A[9][36] [1] = 1'b0;
  assign \A[9][37] [4] = 1'b0;
  assign \A[9][37] [3] = 1'b0;
  assign \A[9][37] [2] = 1'b0;
  assign \A[9][37] [1] = 1'b0;
  assign \A[9][37] [0] = 1'b0;
  assign \A[9][38] [4] = 1'b0;
  assign \A[9][38] [3] = 1'b0;
  assign \A[9][38] [2] = 1'b0;
  assign \A[9][38] [0] = 1'b0;
  assign \A[9][39] [4] = 1'b0;
  assign \A[9][39] [3] = 1'b0;
  assign \A[9][39] [2] = 1'b0;
  assign \A[9][39] [0] = 1'b0;
  assign \A[9][40] [4] = 1'b0;
  assign \A[9][40] [3] = 1'b0;
  assign \A[9][40] [2] = 1'b0;
  assign \A[9][40] [1] = 1'b0;
  assign \A[9][40] [0] = 1'b0;
  assign \A[9][41] [4] = 1'b0;
  assign \A[9][41] [3] = 1'b0;
  assign \A[9][41] [2] = 1'b0;
  assign \A[9][41] [1] = 1'b0;
  assign \A[9][41] [0] = 1'b0;
  assign \A[9][43] [4] = 1'b0;
  assign \A[9][43] [3] = 1'b0;
  assign \A[9][43] [2] = 1'b0;
  assign \A[9][43] [0] = 1'b0;
  assign \A[9][44] [4] = 1'b0;
  assign \A[9][44] [3] = 1'b0;
  assign \A[9][44] [2] = 1'b0;
  assign \A[9][44] [1] = 1'b0;
  assign \A[9][44] [0] = 1'b0;
  assign \A[9][45] [4] = 1'b0;
  assign \A[9][45] [3] = 1'b0;
  assign \A[9][45] [2] = 1'b0;
  assign \A[9][45] [0] = 1'b0;
  assign \A[9][46] [4] = 1'b0;
  assign \A[9][46] [3] = 1'b0;
  assign \A[9][46] [2] = 1'b0;
  assign \A[9][46] [0] = 1'b0;
  assign \A[9][47] [4] = 1'b0;
  assign \A[9][47] [3] = 1'b0;
  assign \A[9][47] [2] = 1'b0;
  assign \A[9][47] [0] = 1'b0;
  assign \A[9][49] [0] = 1'b0;
  assign \A[9][50] [4] = 1'b0;
  assign \A[9][50] [3] = 1'b0;
  assign \A[9][50] [2] = 1'b0;
  assign \A[9][50] [0] = 1'b0;
  assign \A[9][51] [4] = 1'b0;
  assign \A[9][51] [3] = 1'b0;
  assign \A[9][51] [2] = 1'b0;
  assign \A[9][51] [1] = 1'b0;
  assign \A[9][51] [0] = 1'b0;
  assign \A[9][52] [0] = 1'b0;
  assign \A[9][53] [4] = 1'b0;
  assign \A[9][53] [3] = 1'b0;
  assign \A[9][53] [2] = 1'b0;
  assign \A[9][53] [1] = 1'b0;
  assign \A[9][53] [0] = 1'b0;
  assign \A[9][55] [4] = 1'b0;
  assign \A[9][55] [3] = 1'b0;
  assign \A[9][55] [2] = 1'b0;
  assign \A[9][55] [1] = 1'b0;
  assign \A[9][56] [4] = 1'b0;
  assign \A[9][56] [3] = 1'b0;
  assign \A[9][56] [2] = 1'b0;
  assign \A[9][56] [0] = 1'b0;
  assign \A[9][57] [4] = 1'b0;
  assign \A[9][57] [3] = 1'b0;
  assign \A[9][57] [2] = 1'b0;
  assign \A[9][57] [0] = 1'b0;
  assign \A[9][59] [4] = 1'b0;
  assign \A[9][59] [3] = 1'b0;
  assign \A[9][59] [2] = 1'b0;
  assign \A[9][59] [1] = 1'b0;
  assign \A[9][59] [0] = 1'b0;
  assign \A[9][60] [4] = 1'b0;
  assign \A[9][60] [3] = 1'b0;
  assign \A[9][60] [2] = 1'b0;
  assign \A[9][60] [0] = 1'b0;
  assign \A[9][61] [4] = 1'b0;
  assign \A[9][61] [3] = 1'b0;
  assign \A[9][61] [2] = 1'b0;
  assign \A[9][61] [1] = 1'b0;
  assign \A[9][62] [4] = 1'b0;
  assign \A[9][62] [3] = 1'b0;
  assign \A[9][62] [2] = 1'b0;
  assign \A[9][62] [0] = 1'b0;
  assign \A[9][63] [4] = 1'b0;
  assign \A[9][63] [3] = 1'b0;
  assign \A[9][63] [2] = 1'b0;
  assign \A[9][63] [1] = 1'b0;
  assign \A[9][63] [0] = 1'b0;
  assign \A[9][65] [1] = 1'b0;
  assign \A[9][66] [0] = 1'b0;
  assign \A[9][67] [4] = 1'b0;
  assign \A[9][67] [3] = 1'b0;
  assign \A[9][67] [2] = 1'b0;
  assign \A[9][67] [1] = 1'b0;
  assign \A[9][67] [0] = 1'b0;
  assign \A[9][69] [4] = 1'b0;
  assign \A[9][69] [3] = 1'b0;
  assign \A[9][69] [2] = 1'b0;
  assign \A[9][69] [1] = 1'b0;
  assign \A[9][70] [0] = 1'b0;
  assign \A[9][71] [4] = 1'b0;
  assign \A[9][71] [3] = 1'b0;
  assign \A[9][71] [2] = 1'b0;
  assign \A[9][71] [0] = 1'b0;
  assign \A[9][72] [4] = 1'b0;
  assign \A[9][72] [3] = 1'b0;
  assign \A[9][72] [2] = 1'b0;
  assign \A[9][73] [4] = 1'b0;
  assign \A[9][73] [3] = 1'b0;
  assign \A[9][73] [2] = 1'b0;
  assign \A[9][73] [1] = 1'b0;
  assign \A[9][73] [0] = 1'b0;
  assign \A[9][74] [4] = 1'b0;
  assign \A[9][74] [3] = 1'b0;
  assign \A[9][74] [2] = 1'b0;
  assign \A[9][75] [4] = 1'b0;
  assign \A[9][75] [3] = 1'b0;
  assign \A[9][75] [2] = 1'b0;
  assign \A[9][75] [1] = 1'b0;
  assign \A[9][76] [4] = 1'b0;
  assign \A[9][76] [3] = 1'b0;
  assign \A[9][76] [2] = 1'b0;
  assign \A[9][77] [4] = 1'b0;
  assign \A[9][77] [3] = 1'b0;
  assign \A[9][77] [2] = 1'b0;
  assign \A[9][77] [0] = 1'b0;
  assign \A[9][78] [4] = 1'b0;
  assign \A[9][78] [3] = 1'b0;
  assign \A[9][78] [2] = 1'b0;
  assign \A[9][78] [1] = 1'b0;
  assign \A[9][78] [0] = 1'b0;
  assign \A[9][79] [4] = 1'b0;
  assign \A[9][79] [3] = 1'b0;
  assign \A[9][79] [2] = 1'b0;
  assign \A[9][79] [1] = 1'b0;
  assign \A[9][80] [0] = 1'b0;
  assign \A[9][81] [0] = 1'b0;
  assign \A[9][82] [4] = 1'b0;
  assign \A[9][82] [3] = 1'b0;
  assign \A[9][82] [2] = 1'b0;
  assign \A[9][83] [4] = 1'b0;
  assign \A[9][83] [3] = 1'b0;
  assign \A[9][83] [2] = 1'b0;
  assign \A[9][83] [1] = 1'b0;
  assign \A[9][83] [0] = 1'b0;
  assign \A[9][84] [0] = 1'b0;
  assign \A[9][85] [4] = 1'b0;
  assign \A[9][85] [3] = 1'b0;
  assign \A[9][85] [2] = 1'b0;
  assign \A[9][85] [1] = 1'b0;
  assign \A[9][85] [0] = 1'b0;
  assign \A[9][86] [4] = 1'b0;
  assign \A[9][86] [3] = 1'b0;
  assign \A[9][86] [2] = 1'b0;
  assign \A[9][86] [0] = 1'b0;
  assign \A[9][87] [4] = 1'b0;
  assign \A[9][87] [3] = 1'b0;
  assign \A[9][87] [2] = 1'b0;
  assign \A[9][87] [1] = 1'b0;
  assign \A[9][88] [4] = 1'b0;
  assign \A[9][88] [3] = 1'b0;
  assign \A[9][88] [2] = 1'b0;
  assign \A[9][88] [1] = 1'b0;
  assign \A[9][89] [4] = 1'b0;
  assign \A[9][89] [3] = 1'b0;
  assign \A[9][89] [2] = 1'b0;
  assign \A[9][89] [1] = 1'b0;
  assign \A[9][89] [0] = 1'b0;
  assign \A[9][90] [4] = 1'b0;
  assign \A[9][90] [3] = 1'b0;
  assign \A[9][90] [2] = 1'b0;
  assign \A[9][90] [1] = 1'b0;
  assign \A[9][90] [0] = 1'b0;
  assign \A[9][92] [4] = 1'b0;
  assign \A[9][92] [3] = 1'b0;
  assign \A[9][92] [2] = 1'b0;
  assign \A[9][92] [1] = 1'b0;
  assign \A[9][92] [0] = 1'b0;
  assign \A[9][93] [0] = 1'b0;
  assign \A[9][94] [0] = 1'b0;
  assign \A[9][95] [4] = 1'b0;
  assign \A[9][95] [3] = 1'b0;
  assign \A[9][95] [2] = 1'b0;
  assign \A[9][95] [1] = 1'b0;
  assign \A[9][96] [4] = 1'b0;
  assign \A[9][96] [3] = 1'b0;
  assign \A[9][96] [2] = 1'b0;
  assign \A[9][96] [1] = 1'b0;
  assign \A[9][96] [0] = 1'b0;
  assign \A[9][97] [0] = 1'b0;
  assign \A[9][98] [1] = 1'b0;
  assign \A[9][99] [4] = 1'b0;
  assign \A[9][99] [3] = 1'b0;
  assign \A[9][99] [2] = 1'b0;
  assign \A[9][99] [1] = 1'b0;
  assign \A[9][99] [0] = 1'b0;
  assign \A[9][100] [4] = 1'b0;
  assign \A[9][100] [3] = 1'b0;
  assign \A[9][100] [2] = 1'b0;
  assign \A[9][100] [0] = 1'b0;
  assign \A[9][101] [4] = 1'b0;
  assign \A[9][101] [3] = 1'b0;
  assign \A[9][101] [2] = 1'b0;
  assign \A[9][101] [0] = 1'b0;
  assign \A[9][102] [4] = 1'b0;
  assign \A[9][102] [3] = 1'b0;
  assign \A[9][102] [2] = 1'b0;
  assign \A[9][102] [1] = 1'b0;
  assign \A[9][103] [4] = 1'b0;
  assign \A[9][103] [3] = 1'b0;
  assign \A[9][103] [2] = 1'b0;
  assign \A[9][103] [1] = 1'b0;
  assign \A[9][104] [4] = 1'b0;
  assign \A[9][104] [3] = 1'b0;
  assign \A[9][104] [2] = 1'b0;
  assign \A[9][104] [1] = 1'b0;
  assign \A[9][104] [0] = 1'b0;
  assign \A[9][105] [4] = 1'b0;
  assign \A[9][105] [3] = 1'b0;
  assign \A[9][105] [2] = 1'b0;
  assign \A[9][105] [1] = 1'b0;
  assign \A[9][106] [4] = 1'b0;
  assign \A[9][106] [3] = 1'b0;
  assign \A[9][106] [2] = 1'b0;
  assign \A[9][106] [1] = 1'b0;
  assign \A[9][107] [4] = 1'b0;
  assign \A[9][107] [3] = 1'b0;
  assign \A[9][107] [2] = 1'b0;
  assign \A[9][107] [1] = 1'b0;
  assign \A[9][107] [0] = 1'b0;
  assign \A[9][108] [4] = 1'b0;
  assign \A[9][108] [3] = 1'b0;
  assign \A[9][108] [2] = 1'b0;
  assign \A[9][108] [0] = 1'b0;
  assign \A[9][109] [4] = 1'b0;
  assign \A[9][109] [3] = 1'b0;
  assign \A[9][109] [2] = 1'b0;
  assign \A[9][109] [1] = 1'b0;
  assign \A[9][109] [0] = 1'b0;
  assign \A[9][110] [0] = 1'b0;
  assign \A[9][111] [4] = 1'b0;
  assign \A[9][111] [3] = 1'b0;
  assign \A[9][111] [2] = 1'b0;
  assign \A[9][111] [1] = 1'b0;
  assign \A[9][111] [0] = 1'b0;
  assign \A[9][112] [4] = 1'b0;
  assign \A[9][112] [3] = 1'b0;
  assign \A[9][112] [2] = 1'b0;
  assign \A[9][112] [1] = 1'b0;
  assign \A[9][112] [0] = 1'b0;
  assign \A[9][113] [4] = 1'b0;
  assign \A[9][113] [3] = 1'b0;
  assign \A[9][113] [2] = 1'b0;
  assign \A[9][113] [0] = 1'b0;
  assign \A[9][114] [4] = 1'b0;
  assign \A[9][114] [3] = 1'b0;
  assign \A[9][114] [2] = 1'b0;
  assign \A[9][114] [1] = 1'b0;
  assign \A[9][115] [4] = 1'b0;
  assign \A[9][115] [3] = 1'b0;
  assign \A[9][115] [2] = 1'b0;
  assign \A[9][115] [1] = 1'b0;
  assign \A[9][115] [0] = 1'b0;
  assign \A[9][116] [4] = 1'b0;
  assign \A[9][116] [3] = 1'b0;
  assign \A[9][116] [2] = 1'b0;
  assign \A[9][116] [1] = 1'b0;
  assign \A[9][117] [4] = 1'b0;
  assign \A[9][117] [3] = 1'b0;
  assign \A[9][117] [2] = 1'b0;
  assign \A[9][117] [1] = 1'b0;
  assign \A[9][117] [0] = 1'b0;
  assign \A[9][118] [4] = 1'b0;
  assign \A[9][118] [3] = 1'b0;
  assign \A[9][118] [2] = 1'b0;
  assign \A[9][118] [1] = 1'b0;
  assign \A[9][119] [4] = 1'b0;
  assign \A[9][119] [3] = 1'b0;
  assign \A[9][119] [2] = 1'b0;
  assign \A[9][119] [1] = 1'b0;
  assign \A[9][120] [4] = 1'b0;
  assign \A[9][120] [3] = 1'b0;
  assign \A[9][120] [2] = 1'b0;
  assign \A[9][120] [0] = 1'b0;
  assign \A[9][121] [4] = 1'b0;
  assign \A[9][121] [3] = 1'b0;
  assign \A[9][121] [2] = 1'b0;
  assign \A[9][121] [1] = 1'b0;
  assign \A[9][122] [4] = 1'b0;
  assign \A[9][122] [3] = 1'b0;
  assign \A[9][122] [2] = 1'b0;
  assign \A[9][122] [1] = 1'b0;
  assign \A[9][122] [0] = 1'b0;
  assign \A[9][123] [4] = 1'b0;
  assign \A[9][123] [3] = 1'b0;
  assign \A[9][123] [2] = 1'b0;
  assign \A[9][123] [0] = 1'b0;
  assign \A[9][124] [4] = 1'b0;
  assign \A[9][124] [3] = 1'b0;
  assign \A[9][124] [2] = 1'b0;
  assign \A[9][125] [4] = 1'b0;
  assign \A[9][125] [3] = 1'b0;
  assign \A[9][125] [2] = 1'b0;
  assign \A[9][125] [1] = 1'b0;
  assign \A[9][125] [0] = 1'b0;
  assign \A[9][126] [0] = 1'b0;
  assign \A[9][127] [4] = 1'b0;
  assign \A[9][127] [3] = 1'b0;
  assign \A[9][127] [2] = 1'b0;
  assign \A[9][127] [1] = 1'b0;
  assign \A[9][128] [0] = 1'b0;
  assign \A[9][129] [0] = 1'b0;
  assign \A[9][130] [4] = 1'b0;
  assign \A[9][130] [3] = 1'b0;
  assign \A[9][130] [2] = 1'b0;
  assign \A[9][130] [1] = 1'b0;
  assign \A[9][131] [4] = 1'b0;
  assign \A[9][131] [3] = 1'b0;
  assign \A[9][131] [2] = 1'b0;
  assign \A[9][131] [1] = 1'b0;
  assign \A[9][132] [4] = 1'b0;
  assign \A[9][132] [3] = 1'b0;
  assign \A[9][132] [2] = 1'b0;
  assign \A[9][132] [1] = 1'b0;
  assign \A[9][132] [0] = 1'b0;
  assign \A[9][134] [4] = 1'b0;
  assign \A[9][134] [3] = 1'b0;
  assign \A[9][134] [2] = 1'b0;
  assign \A[9][134] [0] = 1'b0;
  assign \A[9][136] [4] = 1'b0;
  assign \A[9][136] [3] = 1'b0;
  assign \A[9][136] [2] = 1'b0;
  assign \A[9][136] [1] = 1'b0;
  assign \A[9][136] [0] = 1'b0;
  assign \A[9][137] [4] = 1'b0;
  assign \A[9][137] [3] = 1'b0;
  assign \A[9][137] [2] = 1'b0;
  assign \A[9][137] [0] = 1'b0;
  assign \A[9][138] [4] = 1'b0;
  assign \A[9][138] [3] = 1'b0;
  assign \A[9][138] [2] = 1'b0;
  assign \A[9][138] [1] = 1'b0;
  assign \A[9][139] [4] = 1'b0;
  assign \A[9][139] [3] = 1'b0;
  assign \A[9][139] [2] = 1'b0;
  assign \A[9][139] [1] = 1'b0;
  assign \A[9][141] [4] = 1'b0;
  assign \A[9][141] [3] = 1'b0;
  assign \A[9][141] [2] = 1'b0;
  assign \A[9][141] [1] = 1'b0;
  assign \A[9][142] [4] = 1'b0;
  assign \A[9][142] [3] = 1'b0;
  assign \A[9][142] [2] = 1'b0;
  assign \A[9][142] [1] = 1'b0;
  assign \A[9][142] [0] = 1'b0;
  assign \A[9][143] [4] = 1'b0;
  assign \A[9][143] [3] = 1'b0;
  assign \A[9][143] [2] = 1'b0;
  assign \A[9][144] [4] = 1'b0;
  assign \A[9][144] [3] = 1'b0;
  assign \A[9][144] [2] = 1'b0;
  assign \A[9][144] [1] = 1'b0;
  assign \A[9][144] [0] = 1'b0;
  assign \A[9][145] [4] = 1'b0;
  assign \A[9][145] [3] = 1'b0;
  assign \A[9][145] [2] = 1'b0;
  assign \A[9][145] [1] = 1'b0;
  assign \A[9][145] [0] = 1'b0;
  assign \A[9][146] [1] = 1'b0;
  assign \A[9][147] [4] = 1'b0;
  assign \A[9][147] [3] = 1'b0;
  assign \A[9][147] [2] = 1'b0;
  assign \A[9][147] [1] = 1'b0;
  assign \A[9][147] [0] = 1'b0;
  assign \A[9][148] [0] = 1'b0;
  assign \A[9][149] [4] = 1'b0;
  assign \A[9][149] [3] = 1'b0;
  assign \A[9][149] [2] = 1'b0;
  assign \A[9][149] [0] = 1'b0;
  assign \A[9][150] [4] = 1'b0;
  assign \A[9][150] [3] = 1'b0;
  assign \A[9][150] [2] = 1'b0;
  assign \A[9][150] [1] = 1'b0;
  assign \A[9][151] [4] = 1'b0;
  assign \A[9][151] [3] = 1'b0;
  assign \A[9][151] [2] = 1'b0;
  assign \A[9][151] [1] = 1'b0;
  assign \A[9][153] [4] = 1'b0;
  assign \A[9][153] [3] = 1'b0;
  assign \A[9][153] [2] = 1'b0;
  assign \A[9][153] [0] = 1'b0;
  assign \A[9][154] [4] = 1'b0;
  assign \A[9][154] [3] = 1'b0;
  assign \A[9][154] [2] = 1'b0;
  assign \A[9][154] [1] = 1'b0;
  assign \A[9][155] [4] = 1'b0;
  assign \A[9][155] [3] = 1'b0;
  assign \A[9][155] [2] = 1'b0;
  assign \A[9][155] [1] = 1'b0;
  assign \A[9][156] [4] = 1'b0;
  assign \A[9][156] [3] = 1'b0;
  assign \A[9][156] [2] = 1'b0;
  assign \A[9][158] [4] = 1'b0;
  assign \A[9][158] [3] = 1'b0;
  assign \A[9][158] [2] = 1'b0;
  assign \A[9][158] [1] = 1'b0;
  assign \A[9][158] [0] = 1'b0;
  assign \A[9][159] [4] = 1'b0;
  assign \A[9][159] [3] = 1'b0;
  assign \A[9][159] [2] = 1'b0;
  assign \A[9][160] [4] = 1'b0;
  assign \A[9][160] [3] = 1'b0;
  assign \A[9][160] [2] = 1'b0;
  assign \A[9][160] [1] = 1'b0;
  assign \A[9][160] [0] = 1'b0;
  assign \A[9][162] [4] = 1'b0;
  assign \A[9][162] [3] = 1'b0;
  assign \A[9][162] [2] = 1'b0;
  assign \A[9][162] [1] = 1'b0;
  assign \A[9][162] [0] = 1'b0;
  assign \A[9][163] [1] = 1'b0;
  assign \A[9][165] [4] = 1'b0;
  assign \A[9][165] [3] = 1'b0;
  assign \A[9][165] [2] = 1'b0;
  assign \A[9][165] [1] = 1'b0;
  assign \A[9][165] [0] = 1'b0;
  assign \A[9][166] [4] = 1'b0;
  assign \A[9][166] [3] = 1'b0;
  assign \A[9][166] [2] = 1'b0;
  assign \A[9][166] [1] = 1'b0;
  assign \A[9][167] [4] = 1'b0;
  assign \A[9][167] [3] = 1'b0;
  assign \A[9][167] [2] = 1'b0;
  assign \A[9][167] [1] = 1'b0;
  assign \A[9][167] [0] = 1'b0;
  assign \A[9][168] [4] = 1'b0;
  assign \A[9][168] [3] = 1'b0;
  assign \A[9][168] [2] = 1'b0;
  assign \A[9][168] [0] = 1'b0;
  assign \A[9][169] [0] = 1'b0;
  assign \A[9][170] [4] = 1'b0;
  assign \A[9][170] [3] = 1'b0;
  assign \A[9][170] [2] = 1'b0;
  assign \A[9][170] [1] = 1'b0;
  assign \A[9][171] [4] = 1'b0;
  assign \A[9][171] [3] = 1'b0;
  assign \A[9][171] [2] = 1'b0;
  assign \A[9][171] [1] = 1'b0;
  assign \A[9][171] [0] = 1'b0;
  assign \A[9][172] [4] = 1'b0;
  assign \A[9][172] [3] = 1'b0;
  assign \A[9][172] [2] = 1'b0;
  assign \A[9][172] [1] = 1'b0;
  assign \A[9][173] [4] = 1'b0;
  assign \A[9][173] [3] = 1'b0;
  assign \A[9][173] [2] = 1'b0;
  assign \A[9][173] [0] = 1'b0;
  assign \A[9][174] [4] = 1'b0;
  assign \A[9][174] [3] = 1'b0;
  assign \A[9][174] [2] = 1'b0;
  assign \A[9][174] [1] = 1'b0;
  assign \A[9][175] [4] = 1'b0;
  assign \A[9][175] [3] = 1'b0;
  assign \A[9][175] [2] = 1'b0;
  assign \A[9][175] [0] = 1'b0;
  assign \A[9][176] [1] = 1'b0;
  assign \A[9][177] [0] = 1'b0;
  assign \A[9][180] [4] = 1'b0;
  assign \A[9][180] [3] = 1'b0;
  assign \A[9][180] [2] = 1'b0;
  assign \A[9][180] [1] = 1'b0;
  assign \A[9][181] [0] = 1'b0;
  assign \A[9][182] [1] = 1'b0;
  assign \A[9][182] [0] = 1'b0;
  assign \A[9][183] [4] = 1'b0;
  assign \A[9][183] [3] = 1'b0;
  assign \A[9][183] [2] = 1'b0;
  assign \A[9][183] [0] = 1'b0;
  assign \A[9][184] [4] = 1'b0;
  assign \A[9][184] [3] = 1'b0;
  assign \A[9][184] [2] = 1'b0;
  assign \A[9][184] [0] = 1'b0;
  assign \A[9][185] [4] = 1'b0;
  assign \A[9][185] [3] = 1'b0;
  assign \A[9][185] [2] = 1'b0;
  assign \A[9][185] [1] = 1'b0;
  assign \A[9][186] [4] = 1'b0;
  assign \A[9][186] [3] = 1'b0;
  assign \A[9][186] [2] = 1'b0;
  assign \A[9][186] [1] = 1'b0;
  assign \A[9][186] [0] = 1'b0;
  assign \A[9][187] [0] = 1'b0;
  assign \A[9][189] [4] = 1'b0;
  assign \A[9][189] [3] = 1'b0;
  assign \A[9][189] [2] = 1'b0;
  assign \A[9][189] [1] = 1'b0;
  assign \A[9][189] [0] = 1'b0;
  assign \A[9][191] [4] = 1'b0;
  assign \A[9][191] [3] = 1'b0;
  assign \A[9][191] [2] = 1'b0;
  assign \A[9][191] [1] = 1'b0;
  assign \A[9][192] [0] = 1'b0;
  assign \A[9][193] [0] = 1'b0;
  assign \A[9][194] [4] = 1'b0;
  assign \A[9][194] [3] = 1'b0;
  assign \A[9][194] [2] = 1'b0;
  assign \A[9][194] [1] = 1'b0;
  assign \A[9][194] [0] = 1'b0;
  assign \A[9][197] [4] = 1'b0;
  assign \A[9][197] [3] = 1'b0;
  assign \A[9][197] [2] = 1'b0;
  assign \A[9][199] [0] = 1'b0;
  assign \A[9][200] [0] = 1'b0;
  assign \A[9][202] [0] = 1'b0;
  assign \A[9][203] [4] = 1'b0;
  assign \A[9][203] [3] = 1'b0;
  assign \A[9][203] [2] = 1'b0;
  assign \A[9][203] [1] = 1'b0;
  assign \A[9][205] [4] = 1'b0;
  assign \A[9][205] [3] = 1'b0;
  assign \A[9][205] [2] = 1'b0;
  assign \A[9][205] [1] = 1'b0;
  assign \A[9][207] [4] = 1'b0;
  assign \A[9][207] [3] = 1'b0;
  assign \A[9][207] [2] = 1'b0;
  assign \A[9][207] [1] = 1'b0;
  assign \A[9][207] [0] = 1'b0;
  assign \A[9][209] [4] = 1'b0;
  assign \A[9][209] [3] = 1'b0;
  assign \A[9][209] [2] = 1'b0;
  assign \A[9][210] [0] = 1'b0;
  assign \A[9][211] [0] = 1'b0;
  assign \A[9][212] [0] = 1'b0;
  assign \A[9][213] [0] = 1'b0;
  assign \A[9][214] [0] = 1'b0;
  assign \A[9][215] [0] = 1'b0;
  assign \A[9][217] [1] = 1'b0;
  assign \A[9][219] [4] = 1'b0;
  assign \A[9][219] [3] = 1'b0;
  assign \A[9][219] [2] = 1'b0;
  assign \A[9][219] [0] = 1'b0;
  assign \A[9][221] [1] = 1'b0;
  assign \A[9][222] [4] = 1'b0;
  assign \A[9][222] [3] = 1'b0;
  assign \A[9][222] [2] = 1'b0;
  assign \A[9][222] [1] = 1'b0;
  assign \A[9][224] [4] = 1'b0;
  assign \A[9][224] [3] = 1'b0;
  assign \A[9][224] [2] = 1'b0;
  assign \A[9][224] [1] = 1'b0;
  assign \A[9][226] [1] = 1'b0;
  assign \A[9][227] [1] = 1'b0;
  assign \A[9][230] [1] = 1'b0;
  assign \A[9][232] [0] = 1'b0;
  assign \A[9][233] [0] = 1'b0;
  assign \A[9][234] [1] = 1'b0;
  assign \A[9][234] [0] = 1'b0;
  assign \A[9][236] [4] = 1'b0;
  assign \A[9][236] [3] = 1'b0;
  assign \A[9][236] [2] = 1'b0;
  assign \A[9][236] [1] = 1'b0;
  assign \A[9][237] [4] = 1'b0;
  assign \A[9][237] [3] = 1'b0;
  assign \A[9][237] [2] = 1'b0;
  assign \A[9][237] [1] = 1'b0;
  assign \A[9][237] [0] = 1'b0;
  assign \A[9][238] [0] = 1'b0;
  assign \A[9][241] [1] = 1'b0;
  assign \A[9][242] [4] = 1'b0;
  assign \A[9][242] [3] = 1'b0;
  assign \A[9][242] [2] = 1'b0;
  assign \A[9][242] [0] = 1'b0;
  assign \A[9][243] [4] = 1'b0;
  assign \A[9][243] [3] = 1'b0;
  assign \A[9][243] [2] = 1'b0;
  assign \A[9][243] [1] = 1'b0;
  assign \A[9][243] [0] = 1'b0;
  assign \A[9][244] [0] = 1'b0;
  assign \A[9][245] [2] = 1'b0;
  assign \A[9][249] [4] = 1'b0;
  assign \A[9][249] [3] = 1'b0;
  assign \A[9][249] [2] = 1'b0;
  assign \A[9][249] [1] = 1'b0;
  assign \A[9][249] [0] = 1'b0;
  assign \A[9][250] [0] = 1'b0;
  assign \A[9][253] [2] = 1'b0;
  assign \A[9][254] [1] = 1'b0;
  assign \A[9][255] [4] = 1'b0;
  assign \A[9][255] [3] = 1'b0;
  assign \A[9][255] [2] = 1'b0;
  assign \A[9][255] [0] = 1'b0;
  assign \A[10][0] [0] = 1'b0;
  assign \A[10][1] [4] = 1'b0;
  assign \A[10][1] [3] = 1'b0;
  assign \A[10][1] [2] = 1'b0;
  assign \A[10][1] [1] = 1'b0;
  assign \A[10][4] [0] = 1'b0;
  assign \A[10][5] [1] = 1'b0;
  assign \A[10][7] [4] = 1'b0;
  assign \A[10][7] [3] = 1'b0;
  assign \A[10][7] [2] = 1'b0;
  assign \A[10][7] [1] = 1'b0;
  assign \A[10][8] [0] = 1'b0;
  assign \A[10][9] [4] = 1'b0;
  assign \A[10][9] [3] = 1'b0;
  assign \A[10][9] [2] = 1'b0;
  assign \A[10][9] [1] = 1'b0;
  assign \A[10][9] [0] = 1'b0;
  assign \A[10][11] [4] = 1'b0;
  assign \A[10][11] [3] = 1'b0;
  assign \A[10][11] [2] = 1'b0;
  assign \A[10][11] [1] = 1'b0;
  assign \A[10][11] [0] = 1'b0;
  assign \A[10][13] [4] = 1'b0;
  assign \A[10][13] [3] = 1'b0;
  assign \A[10][13] [2] = 1'b0;
  assign \A[10][13] [1] = 1'b0;
  assign \A[10][13] [0] = 1'b0;
  assign \A[10][14] [4] = 1'b0;
  assign \A[10][14] [3] = 1'b0;
  assign \A[10][14] [2] = 1'b0;
  assign \A[10][14] [1] = 1'b0;
  assign \A[10][14] [0] = 1'b0;
  assign \A[10][15] [4] = 1'b0;
  assign \A[10][15] [3] = 1'b0;
  assign \A[10][15] [2] = 1'b0;
  assign \A[10][15] [1] = 1'b0;
  assign \A[10][17] [4] = 1'b0;
  assign \A[10][17] [3] = 1'b0;
  assign \A[10][17] [2] = 1'b0;
  assign \A[10][17] [1] = 1'b0;
  assign \A[10][18] [0] = 1'b0;
  assign \A[10][20] [4] = 1'b0;
  assign \A[10][20] [3] = 1'b0;
  assign \A[10][20] [2] = 1'b0;
  assign \A[10][20] [0] = 1'b0;
  assign \A[10][21] [4] = 1'b0;
  assign \A[10][21] [3] = 1'b0;
  assign \A[10][21] [2] = 1'b0;
  assign \A[10][21] [1] = 1'b0;
  assign \A[10][22] [4] = 1'b0;
  assign \A[10][22] [3] = 1'b0;
  assign \A[10][22] [2] = 1'b0;
  assign \A[10][22] [1] = 1'b0;
  assign \A[10][22] [0] = 1'b0;
  assign \A[10][25] [0] = 1'b0;
  assign \A[10][26] [4] = 1'b0;
  assign \A[10][26] [3] = 1'b0;
  assign \A[10][26] [2] = 1'b0;
  assign \A[10][26] [1] = 1'b0;
  assign \A[10][26] [0] = 1'b0;
  assign \A[10][28] [4] = 1'b0;
  assign \A[10][28] [3] = 1'b0;
  assign \A[10][28] [2] = 1'b0;
  assign \A[10][28] [1] = 1'b0;
  assign \A[10][30] [4] = 1'b0;
  assign \A[10][30] [3] = 1'b0;
  assign \A[10][30] [2] = 1'b0;
  assign \A[10][30] [1] = 1'b0;
  assign \A[10][31] [4] = 1'b0;
  assign \A[10][31] [3] = 1'b0;
  assign \A[10][31] [2] = 1'b0;
  assign \A[10][31] [1] = 1'b0;
  assign \A[10][31] [0] = 1'b0;
  assign \A[10][32] [0] = 1'b0;
  assign \A[10][33] [4] = 1'b0;
  assign \A[10][33] [3] = 1'b0;
  assign \A[10][33] [2] = 1'b0;
  assign \A[10][33] [1] = 1'b0;
  assign \A[10][34] [4] = 1'b0;
  assign \A[10][34] [3] = 1'b0;
  assign \A[10][34] [2] = 1'b0;
  assign \A[10][34] [1] = 1'b0;
  assign \A[10][34] [0] = 1'b0;
  assign \A[10][35] [0] = 1'b0;
  assign \A[10][36] [4] = 1'b0;
  assign \A[10][36] [3] = 1'b0;
  assign \A[10][36] [2] = 1'b0;
  assign \A[10][36] [1] = 1'b0;
  assign \A[10][36] [0] = 1'b0;
  assign \A[10][37] [4] = 1'b0;
  assign \A[10][37] [3] = 1'b0;
  assign \A[10][37] [2] = 1'b0;
  assign \A[10][37] [0] = 1'b0;
  assign \A[10][38] [0] = 1'b0;
  assign \A[10][39] [0] = 1'b0;
  assign \A[10][40] [4] = 1'b0;
  assign \A[10][40] [3] = 1'b0;
  assign \A[10][40] [2] = 1'b0;
  assign \A[10][40] [1] = 1'b0;
  assign \A[10][41] [4] = 1'b0;
  assign \A[10][41] [3] = 1'b0;
  assign \A[10][41] [2] = 1'b0;
  assign \A[10][41] [1] = 1'b0;
  assign \A[10][42] [0] = 1'b0;
  assign \A[10][45] [4] = 1'b0;
  assign \A[10][45] [3] = 1'b0;
  assign \A[10][45] [2] = 1'b0;
  assign \A[10][45] [1] = 1'b0;
  assign \A[10][45] [0] = 1'b0;
  assign \A[10][47] [4] = 1'b0;
  assign \A[10][47] [3] = 1'b0;
  assign \A[10][47] [2] = 1'b0;
  assign \A[10][47] [1] = 1'b0;
  assign \A[10][47] [0] = 1'b0;
  assign \A[10][50] [4] = 1'b0;
  assign \A[10][50] [3] = 1'b0;
  assign \A[10][50] [2] = 1'b0;
  assign \A[10][50] [1] = 1'b0;
  assign \A[10][50] [0] = 1'b0;
  assign \A[10][51] [4] = 1'b0;
  assign \A[10][51] [3] = 1'b0;
  assign \A[10][51] [2] = 1'b0;
  assign \A[10][51] [0] = 1'b0;
  assign \A[10][52] [4] = 1'b0;
  assign \A[10][52] [3] = 1'b0;
  assign \A[10][52] [2] = 1'b0;
  assign \A[10][52] [0] = 1'b0;
  assign \A[10][53] [4] = 1'b0;
  assign \A[10][53] [3] = 1'b0;
  assign \A[10][53] [2] = 1'b0;
  assign \A[10][53] [0] = 1'b0;
  assign \A[10][54] [4] = 1'b0;
  assign \A[10][54] [3] = 1'b0;
  assign \A[10][54] [2] = 1'b0;
  assign \A[10][54] [1] = 1'b0;
  assign \A[10][54] [0] = 1'b0;
  assign \A[10][55] [0] = 1'b0;
  assign \A[10][56] [4] = 1'b0;
  assign \A[10][56] [3] = 1'b0;
  assign \A[10][56] [2] = 1'b0;
  assign \A[10][56] [1] = 1'b0;
  assign \A[10][57] [1] = 1'b0;
  assign \A[10][58] [4] = 1'b0;
  assign \A[10][58] [3] = 1'b0;
  assign \A[10][58] [2] = 1'b0;
  assign \A[10][58] [1] = 1'b0;
  assign \A[10][58] [0] = 1'b0;
  assign \A[10][59] [4] = 1'b0;
  assign \A[10][59] [3] = 1'b0;
  assign \A[10][59] [2] = 1'b0;
  assign \A[10][59] [1] = 1'b0;
  assign \A[10][59] [0] = 1'b0;
  assign \A[10][60] [4] = 1'b0;
  assign \A[10][60] [3] = 1'b0;
  assign \A[10][60] [2] = 1'b0;
  assign \A[10][60] [1] = 1'b0;
  assign \A[10][62] [4] = 1'b0;
  assign \A[10][62] [3] = 1'b0;
  assign \A[10][62] [2] = 1'b0;
  assign \A[10][62] [1] = 1'b0;
  assign \A[10][62] [0] = 1'b0;
  assign \A[10][63] [0] = 1'b0;
  assign \A[10][64] [4] = 1'b0;
  assign \A[10][64] [3] = 1'b0;
  assign \A[10][64] [2] = 1'b0;
  assign \A[10][64] [1] = 1'b0;
  assign \A[10][64] [0] = 1'b0;
  assign \A[10][65] [4] = 1'b0;
  assign \A[10][65] [3] = 1'b0;
  assign \A[10][65] [2] = 1'b0;
  assign \A[10][65] [1] = 1'b0;
  assign \A[10][66] [4] = 1'b0;
  assign \A[10][66] [3] = 1'b0;
  assign \A[10][66] [2] = 1'b0;
  assign \A[10][66] [1] = 1'b0;
  assign \A[10][68] [4] = 1'b0;
  assign \A[10][68] [3] = 1'b0;
  assign \A[10][68] [2] = 1'b0;
  assign \A[10][68] [1] = 1'b0;
  assign \A[10][68] [0] = 1'b0;
  assign \A[10][69] [4] = 1'b0;
  assign \A[10][69] [3] = 1'b0;
  assign \A[10][69] [2] = 1'b0;
  assign \A[10][69] [1] = 1'b0;
  assign \A[10][69] [0] = 1'b0;
  assign \A[10][70] [4] = 1'b0;
  assign \A[10][70] [3] = 1'b0;
  assign \A[10][70] [2] = 1'b0;
  assign \A[10][70] [1] = 1'b0;
  assign \A[10][71] [4] = 1'b0;
  assign \A[10][71] [3] = 1'b0;
  assign \A[10][71] [2] = 1'b0;
  assign \A[10][71] [1] = 1'b0;
  assign \A[10][71] [0] = 1'b0;
  assign \A[10][73] [0] = 1'b0;
  assign \A[10][74] [4] = 1'b0;
  assign \A[10][74] [3] = 1'b0;
  assign \A[10][74] [2] = 1'b0;
  assign \A[10][74] [1] = 1'b0;
  assign \A[10][74] [0] = 1'b0;
  assign \A[10][75] [4] = 1'b0;
  assign \A[10][75] [3] = 1'b0;
  assign \A[10][75] [2] = 1'b0;
  assign \A[10][75] [0] = 1'b0;
  assign \A[10][77] [4] = 1'b0;
  assign \A[10][77] [3] = 1'b0;
  assign \A[10][77] [2] = 1'b0;
  assign \A[10][77] [1] = 1'b0;
  assign \A[10][77] [0] = 1'b0;
  assign \A[10][78] [4] = 1'b0;
  assign \A[10][78] [3] = 1'b0;
  assign \A[10][78] [2] = 1'b0;
  assign \A[10][78] [0] = 1'b0;
  assign \A[10][79] [4] = 1'b0;
  assign \A[10][79] [3] = 1'b0;
  assign \A[10][79] [2] = 1'b0;
  assign \A[10][79] [1] = 1'b0;
  assign \A[10][80] [4] = 1'b0;
  assign \A[10][80] [3] = 1'b0;
  assign \A[10][80] [2] = 1'b0;
  assign \A[10][80] [1] = 1'b0;
  assign \A[10][81] [4] = 1'b0;
  assign \A[10][81] [3] = 1'b0;
  assign \A[10][81] [2] = 1'b0;
  assign \A[10][81] [1] = 1'b0;
  assign \A[10][81] [0] = 1'b0;
  assign \A[10][82] [4] = 1'b0;
  assign \A[10][82] [3] = 1'b0;
  assign \A[10][82] [2] = 1'b0;
  assign \A[10][82] [1] = 1'b0;
  assign \A[10][85] [0] = 1'b0;
  assign \A[10][86] [4] = 1'b0;
  assign \A[10][86] [3] = 1'b0;
  assign \A[10][86] [2] = 1'b0;
  assign \A[10][86] [1] = 1'b0;
  assign \A[10][87] [4] = 1'b0;
  assign \A[10][87] [3] = 1'b0;
  assign \A[10][87] [2] = 1'b0;
  assign \A[10][87] [1] = 1'b0;
  assign \A[10][87] [0] = 1'b0;
  assign \A[10][88] [4] = 1'b0;
  assign \A[10][88] [3] = 1'b0;
  assign \A[10][88] [2] = 1'b0;
  assign \A[10][88] [1] = 1'b0;
  assign \A[10][88] [0] = 1'b0;
  assign \A[10][89] [4] = 1'b0;
  assign \A[10][89] [3] = 1'b0;
  assign \A[10][89] [2] = 1'b0;
  assign \A[10][89] [1] = 1'b0;
  assign \A[10][89] [0] = 1'b0;
  assign \A[10][90] [4] = 1'b0;
  assign \A[10][90] [3] = 1'b0;
  assign \A[10][90] [2] = 1'b0;
  assign \A[10][90] [1] = 1'b0;
  assign \A[10][90] [0] = 1'b0;
  assign \A[10][91] [4] = 1'b0;
  assign \A[10][91] [3] = 1'b0;
  assign \A[10][91] [2] = 1'b0;
  assign \A[10][91] [1] = 1'b0;
  assign \A[10][93] [4] = 1'b0;
  assign \A[10][93] [3] = 1'b0;
  assign \A[10][93] [2] = 1'b0;
  assign \A[10][93] [1] = 1'b0;
  assign \A[10][93] [0] = 1'b0;
  assign \A[10][94] [4] = 1'b0;
  assign \A[10][94] [3] = 1'b0;
  assign \A[10][94] [2] = 1'b0;
  assign \A[10][94] [1] = 1'b0;
  assign \A[10][95] [4] = 1'b0;
  assign \A[10][95] [3] = 1'b0;
  assign \A[10][95] [2] = 1'b0;
  assign \A[10][95] [1] = 1'b0;
  assign \A[10][96] [4] = 1'b0;
  assign \A[10][96] [3] = 1'b0;
  assign \A[10][96] [2] = 1'b0;
  assign \A[10][96] [0] = 1'b0;
  assign \A[10][98] [4] = 1'b0;
  assign \A[10][98] [3] = 1'b0;
  assign \A[10][98] [2] = 1'b0;
  assign \A[10][98] [1] = 1'b0;
  assign \A[10][99] [4] = 1'b0;
  assign \A[10][99] [3] = 1'b0;
  assign \A[10][99] [2] = 1'b0;
  assign \A[10][99] [1] = 1'b0;
  assign \A[10][99] [0] = 1'b0;
  assign \A[10][100] [4] = 1'b0;
  assign \A[10][100] [3] = 1'b0;
  assign \A[10][100] [2] = 1'b0;
  assign \A[10][100] [1] = 1'b0;
  assign \A[10][100] [0] = 1'b0;
  assign \A[10][101] [4] = 1'b0;
  assign \A[10][101] [3] = 1'b0;
  assign \A[10][101] [2] = 1'b0;
  assign \A[10][102] [4] = 1'b0;
  assign \A[10][102] [3] = 1'b0;
  assign \A[10][102] [2] = 1'b0;
  assign \A[10][104] [4] = 1'b0;
  assign \A[10][104] [3] = 1'b0;
  assign \A[10][104] [2] = 1'b0;
  assign \A[10][104] [1] = 1'b0;
  assign \A[10][104] [0] = 1'b0;
  assign \A[10][105] [4] = 1'b0;
  assign \A[10][105] [3] = 1'b0;
  assign \A[10][105] [2] = 1'b0;
  assign \A[10][105] [1] = 1'b0;
  assign \A[10][105] [0] = 1'b0;
  assign \A[10][106] [0] = 1'b0;
  assign \A[10][107] [1] = 1'b0;
  assign \A[10][110] [1] = 1'b0;
  assign \A[10][111] [4] = 1'b0;
  assign \A[10][111] [3] = 1'b0;
  assign \A[10][111] [2] = 1'b0;
  assign \A[10][111] [1] = 1'b0;
  assign \A[10][111] [0] = 1'b0;
  assign \A[10][112] [0] = 1'b0;
  assign \A[10][113] [4] = 1'b0;
  assign \A[10][113] [3] = 1'b0;
  assign \A[10][113] [2] = 1'b0;
  assign \A[10][113] [1] = 1'b0;
  assign \A[10][113] [0] = 1'b0;
  assign \A[10][114] [4] = 1'b0;
  assign \A[10][114] [3] = 1'b0;
  assign \A[10][114] [2] = 1'b0;
  assign \A[10][114] [1] = 1'b0;
  assign \A[10][115] [1] = 1'b0;
  assign \A[10][116] [4] = 1'b0;
  assign \A[10][116] [3] = 1'b0;
  assign \A[10][116] [2] = 1'b0;
  assign \A[10][116] [1] = 1'b0;
  assign \A[10][120] [4] = 1'b0;
  assign \A[10][120] [3] = 1'b0;
  assign \A[10][120] [2] = 1'b0;
  assign \A[10][120] [1] = 1'b0;
  assign \A[10][122] [1] = 1'b0;
  assign \A[10][124] [4] = 1'b0;
  assign \A[10][124] [3] = 1'b0;
  assign \A[10][124] [2] = 1'b0;
  assign \A[10][124] [0] = 1'b0;
  assign \A[10][125] [4] = 1'b0;
  assign \A[10][125] [3] = 1'b0;
  assign \A[10][125] [2] = 1'b0;
  assign \A[10][125] [1] = 1'b0;
  assign \A[10][126] [4] = 1'b0;
  assign \A[10][126] [3] = 1'b0;
  assign \A[10][126] [2] = 1'b0;
  assign \A[10][126] [1] = 1'b0;
  assign \A[10][127] [4] = 1'b0;
  assign \A[10][127] [3] = 1'b0;
  assign \A[10][127] [2] = 1'b0;
  assign \A[10][127] [1] = 1'b0;
  assign \A[10][128] [4] = 1'b0;
  assign \A[10][128] [3] = 1'b0;
  assign \A[10][128] [2] = 1'b0;
  assign \A[10][128] [1] = 1'b0;
  assign \A[10][129] [4] = 1'b0;
  assign \A[10][129] [3] = 1'b0;
  assign \A[10][129] [2] = 1'b0;
  assign \A[10][129] [1] = 1'b0;
  assign \A[10][129] [0] = 1'b0;
  assign \A[10][130] [4] = 1'b0;
  assign \A[10][130] [3] = 1'b0;
  assign \A[10][130] [2] = 1'b0;
  assign \A[10][130] [1] = 1'b0;
  assign \A[10][130] [0] = 1'b0;
  assign \A[10][131] [4] = 1'b0;
  assign \A[10][131] [3] = 1'b0;
  assign \A[10][131] [2] = 1'b0;
  assign \A[10][131] [1] = 1'b0;
  assign \A[10][132] [4] = 1'b0;
  assign \A[10][132] [3] = 1'b0;
  assign \A[10][132] [2] = 1'b0;
  assign \A[10][132] [1] = 1'b0;
  assign \A[10][132] [0] = 1'b0;
  assign \A[10][133] [4] = 1'b0;
  assign \A[10][133] [3] = 1'b0;
  assign \A[10][133] [2] = 1'b0;
  assign \A[10][133] [1] = 1'b0;
  assign \A[10][134] [4] = 1'b0;
  assign \A[10][134] [3] = 1'b0;
  assign \A[10][134] [2] = 1'b0;
  assign \A[10][134] [1] = 1'b0;
  assign \A[10][136] [0] = 1'b0;
  assign \A[10][137] [4] = 1'b0;
  assign \A[10][137] [3] = 1'b0;
  assign \A[10][137] [2] = 1'b0;
  assign \A[10][137] [1] = 1'b0;
  assign \A[10][137] [0] = 1'b0;
  assign \A[10][138] [4] = 1'b0;
  assign \A[10][138] [3] = 1'b0;
  assign \A[10][138] [2] = 1'b0;
  assign \A[10][138] [1] = 1'b0;
  assign \A[10][138] [0] = 1'b0;
  assign \A[10][139] [4] = 1'b0;
  assign \A[10][139] [3] = 1'b0;
  assign \A[10][139] [2] = 1'b0;
  assign \A[10][139] [0] = 1'b0;
  assign \A[10][140] [0] = 1'b0;
  assign \A[10][141] [4] = 1'b0;
  assign \A[10][141] [3] = 1'b0;
  assign \A[10][141] [2] = 1'b0;
  assign \A[10][141] [1] = 1'b0;
  assign \A[10][141] [0] = 1'b0;
  assign \A[10][142] [4] = 1'b0;
  assign \A[10][142] [3] = 1'b0;
  assign \A[10][142] [2] = 1'b0;
  assign \A[10][142] [1] = 1'b0;
  assign \A[10][143] [4] = 1'b0;
  assign \A[10][143] [3] = 1'b0;
  assign \A[10][143] [2] = 1'b0;
  assign \A[10][143] [1] = 1'b0;
  assign \A[10][143] [0] = 1'b0;
  assign \A[10][145] [1] = 1'b0;
  assign \A[10][148] [4] = 1'b0;
  assign \A[10][148] [3] = 1'b0;
  assign \A[10][148] [2] = 1'b0;
  assign \A[10][148] [1] = 1'b0;
  assign \A[10][148] [0] = 1'b0;
  assign \A[10][151] [4] = 1'b0;
  assign \A[10][151] [3] = 1'b0;
  assign \A[10][151] [2] = 1'b0;
  assign \A[10][151] [1] = 1'b0;
  assign \A[10][152] [4] = 1'b0;
  assign \A[10][152] [3] = 1'b0;
  assign \A[10][152] [2] = 1'b0;
  assign \A[10][152] [0] = 1'b0;
  assign \A[10][153] [4] = 1'b0;
  assign \A[10][153] [3] = 1'b0;
  assign \A[10][153] [2] = 1'b0;
  assign \A[10][153] [1] = 1'b0;
  assign \A[10][153] [0] = 1'b0;
  assign \A[10][154] [4] = 1'b0;
  assign \A[10][154] [3] = 1'b0;
  assign \A[10][154] [2] = 1'b0;
  assign \A[10][154] [1] = 1'b0;
  assign \A[10][154] [0] = 1'b0;
  assign \A[10][155] [4] = 1'b0;
  assign \A[10][155] [3] = 1'b0;
  assign \A[10][155] [2] = 1'b0;
  assign \A[10][155] [1] = 1'b0;
  assign \A[10][156] [4] = 1'b0;
  assign \A[10][156] [3] = 1'b0;
  assign \A[10][156] [2] = 1'b0;
  assign \A[10][156] [1] = 1'b0;
  assign \A[10][156] [0] = 1'b0;
  assign \A[10][157] [4] = 1'b0;
  assign \A[10][157] [3] = 1'b0;
  assign \A[10][157] [2] = 1'b0;
  assign \A[10][157] [0] = 1'b0;
  assign \A[10][158] [4] = 1'b0;
  assign \A[10][158] [3] = 1'b0;
  assign \A[10][158] [2] = 1'b0;
  assign \A[10][158] [1] = 1'b0;
  assign \A[10][158] [0] = 1'b0;
  assign \A[10][159] [4] = 1'b0;
  assign \A[10][159] [3] = 1'b0;
  assign \A[10][159] [2] = 1'b0;
  assign \A[10][159] [0] = 1'b0;
  assign \A[10][160] [4] = 1'b0;
  assign \A[10][160] [3] = 1'b0;
  assign \A[10][160] [2] = 1'b0;
  assign \A[10][160] [1] = 1'b0;
  assign \A[10][160] [0] = 1'b0;
  assign \A[10][161] [4] = 1'b0;
  assign \A[10][161] [3] = 1'b0;
  assign \A[10][161] [2] = 1'b0;
  assign \A[10][161] [1] = 1'b0;
  assign \A[10][161] [0] = 1'b0;
  assign \A[10][162] [4] = 1'b0;
  assign \A[10][162] [3] = 1'b0;
  assign \A[10][162] [2] = 1'b0;
  assign \A[10][162] [0] = 1'b0;
  assign \A[10][163] [4] = 1'b0;
  assign \A[10][163] [3] = 1'b0;
  assign \A[10][163] [2] = 1'b0;
  assign \A[10][164] [4] = 1'b0;
  assign \A[10][164] [3] = 1'b0;
  assign \A[10][164] [2] = 1'b0;
  assign \A[10][164] [1] = 1'b0;
  assign \A[10][164] [0] = 1'b0;
  assign \A[10][166] [4] = 1'b0;
  assign \A[10][166] [3] = 1'b0;
  assign \A[10][166] [2] = 1'b0;
  assign \A[10][166] [0] = 1'b0;
  assign \A[10][167] [4] = 1'b0;
  assign \A[10][167] [3] = 1'b0;
  assign \A[10][167] [2] = 1'b0;
  assign \A[10][167] [1] = 1'b0;
  assign \A[10][168] [1] = 1'b0;
  assign \A[10][169] [4] = 1'b0;
  assign \A[10][169] [3] = 1'b0;
  assign \A[10][169] [2] = 1'b0;
  assign \A[10][169] [1] = 1'b0;
  assign \A[10][169] [0] = 1'b0;
  assign \A[10][171] [4] = 1'b0;
  assign \A[10][171] [3] = 1'b0;
  assign \A[10][171] [2] = 1'b0;
  assign \A[10][171] [1] = 1'b0;
  assign \A[10][172] [0] = 1'b0;
  assign \A[10][173] [4] = 1'b0;
  assign \A[10][173] [3] = 1'b0;
  assign \A[10][173] [2] = 1'b0;
  assign \A[10][173] [1] = 1'b0;
  assign \A[10][173] [0] = 1'b0;
  assign \A[10][174] [4] = 1'b0;
  assign \A[10][174] [3] = 1'b0;
  assign \A[10][174] [2] = 1'b0;
  assign \A[10][174] [1] = 1'b0;
  assign \A[10][174] [0] = 1'b0;
  assign \A[10][176] [4] = 1'b0;
  assign \A[10][176] [3] = 1'b0;
  assign \A[10][176] [2] = 1'b0;
  assign \A[10][176] [1] = 1'b0;
  assign \A[10][176] [0] = 1'b0;
  assign \A[10][177] [4] = 1'b0;
  assign \A[10][177] [3] = 1'b0;
  assign \A[10][177] [2] = 1'b0;
  assign \A[10][177] [1] = 1'b0;
  assign \A[10][179] [4] = 1'b0;
  assign \A[10][179] [3] = 1'b0;
  assign \A[10][179] [2] = 1'b0;
  assign \A[10][179] [0] = 1'b0;
  assign \A[10][181] [0] = 1'b0;
  assign \A[10][184] [4] = 1'b0;
  assign \A[10][184] [3] = 1'b0;
  assign \A[10][184] [2] = 1'b0;
  assign \A[10][184] [1] = 1'b0;
  assign \A[10][184] [0] = 1'b0;
  assign \A[10][185] [4] = 1'b0;
  assign \A[10][185] [3] = 1'b0;
  assign \A[10][185] [2] = 1'b0;
  assign \A[10][185] [1] = 1'b0;
  assign \A[10][185] [0] = 1'b0;
  assign \A[10][186] [1] = 1'b0;
  assign \A[10][187] [0] = 1'b0;
  assign \A[10][188] [4] = 1'b0;
  assign \A[10][188] [3] = 1'b0;
  assign \A[10][188] [2] = 1'b0;
  assign \A[10][188] [1] = 1'b0;
  assign \A[10][189] [4] = 1'b0;
  assign \A[10][189] [3] = 1'b0;
  assign \A[10][189] [2] = 1'b0;
  assign \A[10][189] [1] = 1'b0;
  assign \A[10][190] [4] = 1'b0;
  assign \A[10][190] [3] = 1'b0;
  assign \A[10][190] [2] = 1'b0;
  assign \A[10][190] [1] = 1'b0;
  assign \A[10][191] [4] = 1'b0;
  assign \A[10][191] [3] = 1'b0;
  assign \A[10][191] [2] = 1'b0;
  assign \A[10][191] [1] = 1'b0;
  assign \A[10][191] [0] = 1'b0;
  assign \A[10][192] [4] = 1'b0;
  assign \A[10][192] [3] = 1'b0;
  assign \A[10][192] [2] = 1'b0;
  assign \A[10][192] [1] = 1'b0;
  assign \A[10][192] [0] = 1'b0;
  assign \A[10][193] [4] = 1'b0;
  assign \A[10][193] [3] = 1'b0;
  assign \A[10][193] [2] = 1'b0;
  assign \A[10][193] [1] = 1'b0;
  assign \A[10][195] [4] = 1'b0;
  assign \A[10][195] [3] = 1'b0;
  assign \A[10][195] [2] = 1'b0;
  assign \A[10][195] [1] = 1'b0;
  assign \A[10][196] [0] = 1'b0;
  assign \A[10][197] [0] = 1'b0;
  assign \A[10][198] [4] = 1'b0;
  assign \A[10][198] [3] = 1'b0;
  assign \A[10][198] [2] = 1'b0;
  assign \A[10][198] [1] = 1'b0;
  assign \A[10][199] [4] = 1'b0;
  assign \A[10][199] [3] = 1'b0;
  assign \A[10][199] [2] = 1'b0;
  assign \A[10][199] [1] = 1'b0;
  assign \A[10][199] [0] = 1'b0;
  assign \A[10][201] [4] = 1'b0;
  assign \A[10][201] [3] = 1'b0;
  assign \A[10][201] [2] = 1'b0;
  assign \A[10][201] [1] = 1'b0;
  assign \A[10][201] [0] = 1'b0;
  assign \A[10][203] [4] = 1'b0;
  assign \A[10][203] [3] = 1'b0;
  assign \A[10][203] [2] = 1'b0;
  assign \A[10][203] [1] = 1'b0;
  assign \A[10][204] [4] = 1'b0;
  assign \A[10][204] [3] = 1'b0;
  assign \A[10][204] [2] = 1'b0;
  assign \A[10][204] [1] = 1'b0;
  assign \A[10][205] [4] = 1'b0;
  assign \A[10][205] [3] = 1'b0;
  assign \A[10][205] [2] = 1'b0;
  assign \A[10][205] [1] = 1'b0;
  assign \A[10][205] [0] = 1'b0;
  assign \A[10][206] [4] = 1'b0;
  assign \A[10][206] [3] = 1'b0;
  assign \A[10][206] [2] = 1'b0;
  assign \A[10][206] [1] = 1'b0;
  assign \A[10][207] [4] = 1'b0;
  assign \A[10][207] [3] = 1'b0;
  assign \A[10][207] [2] = 1'b0;
  assign \A[10][207] [1] = 1'b0;
  assign \A[10][208] [4] = 1'b0;
  assign \A[10][208] [3] = 1'b0;
  assign \A[10][208] [2] = 1'b0;
  assign \A[10][208] [1] = 1'b0;
  assign \A[10][209] [0] = 1'b0;
  assign \A[10][212] [4] = 1'b0;
  assign \A[10][212] [3] = 1'b0;
  assign \A[10][212] [2] = 1'b0;
  assign \A[10][212] [0] = 1'b0;
  assign \A[10][214] [4] = 1'b0;
  assign \A[10][214] [3] = 1'b0;
  assign \A[10][214] [2] = 1'b0;
  assign \A[10][214] [1] = 1'b0;
  assign \A[10][214] [0] = 1'b0;
  assign \A[10][215] [4] = 1'b0;
  assign \A[10][215] [3] = 1'b0;
  assign \A[10][215] [2] = 1'b0;
  assign \A[10][215] [0] = 1'b0;
  assign \A[10][216] [0] = 1'b0;
  assign \A[10][217] [4] = 1'b0;
  assign \A[10][217] [3] = 1'b0;
  assign \A[10][217] [2] = 1'b0;
  assign \A[10][217] [1] = 1'b0;
  assign \A[10][217] [0] = 1'b0;
  assign \A[10][218] [4] = 1'b0;
  assign \A[10][218] [3] = 1'b0;
  assign \A[10][218] [2] = 1'b0;
  assign \A[10][218] [1] = 1'b0;
  assign \A[10][218] [0] = 1'b0;
  assign \A[10][219] [4] = 1'b0;
  assign \A[10][219] [3] = 1'b0;
  assign \A[10][219] [2] = 1'b0;
  assign \A[10][219] [0] = 1'b0;
  assign \A[10][220] [4] = 1'b0;
  assign \A[10][220] [3] = 1'b0;
  assign \A[10][220] [2] = 1'b0;
  assign \A[10][222] [4] = 1'b0;
  assign \A[10][222] [3] = 1'b0;
  assign \A[10][222] [2] = 1'b0;
  assign \A[10][222] [1] = 1'b0;
  assign \A[10][222] [0] = 1'b0;
  assign \A[10][223] [4] = 1'b0;
  assign \A[10][223] [3] = 1'b0;
  assign \A[10][223] [2] = 1'b0;
  assign \A[10][223] [0] = 1'b0;
  assign \A[10][224] [4] = 1'b0;
  assign \A[10][224] [3] = 1'b0;
  assign \A[10][224] [2] = 1'b0;
  assign \A[10][224] [1] = 1'b0;
  assign \A[10][225] [4] = 1'b0;
  assign \A[10][225] [3] = 1'b0;
  assign \A[10][225] [2] = 1'b0;
  assign \A[10][225] [1] = 1'b0;
  assign \A[10][225] [0] = 1'b0;
  assign \A[10][226] [4] = 1'b0;
  assign \A[10][226] [3] = 1'b0;
  assign \A[10][226] [2] = 1'b0;
  assign \A[10][226] [0] = 1'b0;
  assign \A[10][228] [4] = 1'b0;
  assign \A[10][228] [3] = 1'b0;
  assign \A[10][228] [2] = 1'b0;
  assign \A[10][228] [0] = 1'b0;
  assign \A[10][230] [4] = 1'b0;
  assign \A[10][230] [3] = 1'b0;
  assign \A[10][230] [2] = 1'b0;
  assign \A[10][230] [1] = 1'b0;
  assign \A[10][232] [0] = 1'b0;
  assign \A[10][233] [0] = 1'b0;
  assign \A[10][234] [4] = 1'b0;
  assign \A[10][234] [3] = 1'b0;
  assign \A[10][234] [2] = 1'b0;
  assign \A[10][234] [1] = 1'b0;
  assign \A[10][234] [0] = 1'b0;
  assign \A[10][235] [4] = 1'b0;
  assign \A[10][235] [3] = 1'b0;
  assign \A[10][235] [2] = 1'b0;
  assign \A[10][235] [1] = 1'b0;
  assign \A[10][235] [0] = 1'b0;
  assign \A[10][236] [1] = 1'b0;
  assign \A[10][237] [4] = 1'b0;
  assign \A[10][237] [3] = 1'b0;
  assign \A[10][237] [2] = 1'b0;
  assign \A[10][237] [1] = 1'b0;
  assign \A[10][237] [0] = 1'b0;
  assign \A[10][238] [4] = 1'b0;
  assign \A[10][238] [3] = 1'b0;
  assign \A[10][238] [2] = 1'b0;
  assign \A[10][238] [1] = 1'b0;
  assign \A[10][238] [0] = 1'b0;
  assign \A[10][241] [4] = 1'b0;
  assign \A[10][241] [3] = 1'b0;
  assign \A[10][241] [2] = 1'b0;
  assign \A[10][241] [1] = 1'b0;
  assign \A[10][242] [4] = 1'b0;
  assign \A[10][242] [3] = 1'b0;
  assign \A[10][242] [2] = 1'b0;
  assign \A[10][242] [1] = 1'b0;
  assign \A[10][243] [4] = 1'b0;
  assign \A[10][243] [3] = 1'b0;
  assign \A[10][243] [2] = 1'b0;
  assign \A[10][243] [1] = 1'b0;
  assign \A[10][245] [4] = 1'b0;
  assign \A[10][245] [3] = 1'b0;
  assign \A[10][245] [2] = 1'b0;
  assign \A[10][245] [1] = 1'b0;
  assign \A[10][245] [0] = 1'b0;
  assign \A[10][247] [4] = 1'b0;
  assign \A[10][247] [3] = 1'b0;
  assign \A[10][247] [2] = 1'b0;
  assign \A[10][247] [1] = 1'b0;
  assign \A[10][248] [0] = 1'b0;
  assign \A[10][249] [4] = 1'b0;
  assign \A[10][249] [3] = 1'b0;
  assign \A[10][249] [2] = 1'b0;
  assign \A[10][249] [1] = 1'b0;
  assign \A[10][249] [0] = 1'b0;
  assign \A[10][252] [4] = 1'b0;
  assign \A[10][252] [3] = 1'b0;
  assign \A[10][252] [2] = 1'b0;
  assign \A[10][252] [1] = 1'b0;
  assign \A[10][254] [4] = 1'b0;
  assign \A[10][254] [3] = 1'b0;
  assign \A[10][254] [2] = 1'b0;
  assign \A[10][254] [1] = 1'b0;
  assign \A[10][254] [0] = 1'b0;
  assign \A[10][255] [4] = 1'b0;
  assign \A[10][255] [3] = 1'b0;
  assign \A[10][255] [2] = 1'b0;
  assign \A[10][255] [1] = 1'b0;
  assign \A[10][255] [0] = 1'b0;
  assign \A[11][0] [4] = 1'b0;
  assign \A[11][0] [3] = 1'b0;
  assign \A[11][0] [1] = 1'b0;
  assign \A[11][0] [0] = 1'b0;
  assign \A[11][1] [0] = 1'b0;
  assign \A[11][3] [4] = 1'b0;
  assign \A[11][3] [3] = 1'b0;
  assign \A[11][3] [2] = 1'b0;
  assign \A[11][3] [1] = 1'b0;
  assign \A[11][3] [0] = 1'b0;
  assign \A[11][5] [1] = 1'b0;
  assign \A[11][6] [4] = 1'b0;
  assign \A[11][6] [3] = 1'b0;
  assign \A[11][6] [2] = 1'b0;
  assign \A[11][6] [1] = 1'b0;
  assign \A[11][6] [0] = 1'b0;
  assign \A[11][7] [4] = 1'b0;
  assign \A[11][7] [3] = 1'b0;
  assign \A[11][7] [2] = 1'b0;
  assign \A[11][7] [1] = 1'b0;
  assign \A[11][8] [2] = 1'b0;
  assign \A[11][9] [0] = 1'b0;
  assign \A[11][10] [4] = 1'b0;
  assign \A[11][10] [3] = 1'b0;
  assign \A[11][10] [2] = 1'b0;
  assign \A[11][10] [1] = 1'b0;
  assign \A[11][10] [0] = 1'b0;
  assign \A[11][11] [1] = 1'b0;
  assign \A[11][12] [0] = 1'b0;
  assign \A[11][13] [4] = 1'b0;
  assign \A[11][13] [3] = 1'b0;
  assign \A[11][13] [2] = 1'b0;
  assign \A[11][13] [1] = 1'b0;
  assign \A[11][14] [0] = 1'b0;
  assign \A[11][15] [4] = 1'b0;
  assign \A[11][15] [3] = 1'b0;
  assign \A[11][15] [2] = 1'b0;
  assign \A[11][15] [1] = 1'b0;
  assign \A[11][16] [1] = 1'b0;
  assign \A[11][17] [4] = 1'b0;
  assign \A[11][17] [3] = 1'b0;
  assign \A[11][17] [2] = 1'b0;
  assign \A[11][17] [1] = 1'b0;
  assign \A[11][17] [0] = 1'b0;
  assign \A[11][19] [4] = 1'b0;
  assign \A[11][19] [3] = 1'b0;
  assign \A[11][19] [2] = 1'b0;
  assign \A[11][19] [1] = 1'b0;
  assign \A[11][19] [0] = 1'b0;
  assign \A[11][22] [2] = 1'b0;
  assign \A[11][24] [1] = 1'b0;
  assign \A[11][26] [4] = 1'b0;
  assign \A[11][26] [3] = 1'b0;
  assign \A[11][26] [2] = 1'b0;
  assign \A[11][26] [1] = 1'b0;
  assign \A[11][26] [0] = 1'b0;
  assign \A[11][27] [4] = 1'b0;
  assign \A[11][27] [3] = 1'b0;
  assign \A[11][27] [2] = 1'b0;
  assign \A[11][27] [0] = 1'b0;
  assign \A[11][28] [4] = 1'b0;
  assign \A[11][28] [3] = 1'b0;
  assign \A[11][28] [2] = 1'b0;
  assign \A[11][28] [1] = 1'b0;
  assign \A[11][28] [0] = 1'b0;
  assign \A[11][30] [4] = 1'b0;
  assign \A[11][30] [3] = 1'b0;
  assign \A[11][30] [2] = 1'b0;
  assign \A[11][30] [0] = 1'b0;
  assign \A[11][32] [0] = 1'b0;
  assign \A[11][34] [4] = 1'b0;
  assign \A[11][34] [3] = 1'b0;
  assign \A[11][34] [2] = 1'b0;
  assign \A[11][34] [1] = 1'b0;
  assign \A[11][37] [4] = 1'b0;
  assign \A[11][37] [3] = 1'b0;
  assign \A[11][37] [2] = 1'b0;
  assign \A[11][37] [0] = 1'b0;
  assign \A[11][38] [4] = 1'b0;
  assign \A[11][38] [3] = 1'b0;
  assign \A[11][38] [2] = 1'b0;
  assign \A[11][38] [1] = 1'b0;
  assign \A[11][38] [0] = 1'b0;
  assign \A[11][39] [4] = 1'b0;
  assign \A[11][39] [3] = 1'b0;
  assign \A[11][39] [2] = 1'b0;
  assign \A[11][39] [1] = 1'b0;
  assign \A[11][39] [0] = 1'b0;
  assign \A[11][40] [0] = 1'b0;
  assign \A[11][41] [0] = 1'b0;
  assign \A[11][42] [4] = 1'b0;
  assign \A[11][42] [3] = 1'b0;
  assign \A[11][42] [2] = 1'b0;
  assign \A[11][42] [1] = 1'b0;
  assign \A[11][42] [0] = 1'b0;
  assign \A[11][43] [4] = 1'b0;
  assign \A[11][43] [3] = 1'b0;
  assign \A[11][43] [2] = 1'b0;
  assign \A[11][43] [1] = 1'b0;
  assign \A[11][43] [0] = 1'b0;
  assign \A[11][44] [4] = 1'b0;
  assign \A[11][44] [3] = 1'b0;
  assign \A[11][44] [2] = 1'b0;
  assign \A[11][44] [0] = 1'b0;
  assign \A[11][45] [4] = 1'b0;
  assign \A[11][45] [3] = 1'b0;
  assign \A[11][45] [2] = 1'b0;
  assign \A[11][45] [1] = 1'b0;
  assign \A[11][46] [1] = 1'b0;
  assign \A[11][47] [4] = 1'b0;
  assign \A[11][47] [3] = 1'b0;
  assign \A[11][47] [2] = 1'b0;
  assign \A[11][47] [1] = 1'b0;
  assign \A[11][47] [0] = 1'b0;
  assign \A[11][48] [4] = 1'b0;
  assign \A[11][48] [3] = 1'b0;
  assign \A[11][48] [2] = 1'b0;
  assign \A[11][48] [1] = 1'b0;
  assign \A[11][48] [0] = 1'b0;
  assign \A[11][50] [1] = 1'b0;
  assign \A[11][51] [4] = 1'b0;
  assign \A[11][51] [3] = 1'b0;
  assign \A[11][51] [2] = 1'b0;
  assign \A[11][51] [1] = 1'b0;
  assign \A[11][51] [0] = 1'b0;
  assign \A[11][52] [4] = 1'b0;
  assign \A[11][52] [3] = 1'b0;
  assign \A[11][52] [2] = 1'b0;
  assign \A[11][52] [1] = 1'b0;
  assign \A[11][53] [4] = 1'b0;
  assign \A[11][53] [3] = 1'b0;
  assign \A[11][53] [2] = 1'b0;
  assign \A[11][53] [1] = 1'b0;
  assign \A[11][53] [0] = 1'b0;
  assign \A[11][54] [4] = 1'b0;
  assign \A[11][54] [3] = 1'b0;
  assign \A[11][54] [2] = 1'b0;
  assign \A[11][54] [1] = 1'b0;
  assign \A[11][54] [0] = 1'b0;
  assign \A[11][55] [0] = 1'b0;
  assign \A[11][56] [4] = 1'b0;
  assign \A[11][56] [3] = 1'b0;
  assign \A[11][56] [2] = 1'b0;
  assign \A[11][56] [0] = 1'b0;
  assign \A[11][57] [4] = 1'b0;
  assign \A[11][57] [3] = 1'b0;
  assign \A[11][57] [2] = 1'b0;
  assign \A[11][57] [1] = 1'b0;
  assign \A[11][58] [4] = 1'b0;
  assign \A[11][58] [3] = 1'b0;
  assign \A[11][58] [2] = 1'b0;
  assign \A[11][58] [1] = 1'b0;
  assign \A[11][60] [2] = 1'b0;
  assign \A[11][62] [0] = 1'b0;
  assign \A[11][63] [2] = 1'b0;
  assign \A[11][64] [4] = 1'b0;
  assign \A[11][64] [3] = 1'b0;
  assign \A[11][64] [2] = 1'b0;
  assign \A[11][64] [1] = 1'b0;
  assign \A[11][64] [0] = 1'b0;
  assign \A[11][65] [0] = 1'b0;
  assign \A[11][67] [4] = 1'b0;
  assign \A[11][67] [3] = 1'b0;
  assign \A[11][67] [2] = 1'b0;
  assign \A[11][67] [1] = 1'b0;
  assign \A[11][67] [0] = 1'b0;
  assign \A[11][68] [4] = 1'b0;
  assign \A[11][68] [3] = 1'b0;
  assign \A[11][68] [2] = 1'b0;
  assign \A[11][68] [0] = 1'b0;
  assign \A[11][69] [4] = 1'b0;
  assign \A[11][69] [3] = 1'b0;
  assign \A[11][69] [2] = 1'b0;
  assign \A[11][69] [0] = 1'b0;
  assign \A[11][70] [4] = 1'b0;
  assign \A[11][70] [3] = 1'b0;
  assign \A[11][70] [2] = 1'b0;
  assign \A[11][70] [1] = 1'b0;
  assign \A[11][71] [1] = 1'b0;
  assign \A[11][72] [4] = 1'b0;
  assign \A[11][72] [3] = 1'b0;
  assign \A[11][72] [2] = 1'b0;
  assign \A[11][72] [1] = 1'b0;
  assign \A[11][72] [0] = 1'b0;
  assign \A[11][73] [4] = 1'b0;
  assign \A[11][73] [3] = 1'b0;
  assign \A[11][73] [1] = 1'b0;
  assign \A[11][73] [0] = 1'b0;
  assign \A[11][74] [0] = 1'b0;
  assign \A[11][75] [0] = 1'b0;
  assign \A[11][76] [1] = 1'b0;
  assign \A[11][77] [0] = 1'b0;
  assign \A[11][79] [0] = 1'b0;
  assign \A[11][80] [4] = 1'b0;
  assign \A[11][80] [3] = 1'b0;
  assign \A[11][80] [2] = 1'b0;
  assign \A[11][80] [1] = 1'b0;
  assign \A[11][81] [4] = 1'b0;
  assign \A[11][81] [3] = 1'b0;
  assign \A[11][81] [2] = 1'b0;
  assign \A[11][81] [0] = 1'b0;
  assign \A[11][82] [4] = 1'b0;
  assign \A[11][82] [3] = 1'b0;
  assign \A[11][82] [2] = 1'b0;
  assign \A[11][82] [1] = 1'b0;
  assign \A[11][82] [0] = 1'b0;
  assign \A[11][84] [4] = 1'b0;
  assign \A[11][84] [3] = 1'b0;
  assign \A[11][84] [2] = 1'b0;
  assign \A[11][84] [1] = 1'b0;
  assign \A[11][85] [0] = 1'b0;
  assign \A[11][87] [4] = 1'b0;
  assign \A[11][87] [3] = 1'b0;
  assign \A[11][87] [2] = 1'b0;
  assign \A[11][87] [1] = 1'b0;
  assign \A[11][87] [0] = 1'b0;
  assign \A[11][89] [1] = 1'b0;
  assign \A[11][89] [0] = 1'b0;
  assign \A[11][91] [1] = 1'b0;
  assign \A[11][92] [1] = 1'b0;
  assign \A[11][92] [0] = 1'b0;
  assign \A[11][93] [4] = 1'b0;
  assign \A[11][93] [3] = 1'b0;
  assign \A[11][93] [2] = 1'b0;
  assign \A[11][93] [1] = 1'b0;
  assign \A[11][93] [0] = 1'b0;
  assign \A[11][94] [1] = 1'b0;
  assign \A[11][95] [4] = 1'b0;
  assign \A[11][95] [3] = 1'b0;
  assign \A[11][95] [2] = 1'b0;
  assign \A[11][95] [1] = 1'b0;
  assign \A[11][95] [0] = 1'b0;
  assign \A[11][96] [4] = 1'b0;
  assign \A[11][96] [3] = 1'b0;
  assign \A[11][96] [2] = 1'b0;
  assign \A[11][96] [0] = 1'b0;
  assign \A[11][97] [4] = 1'b0;
  assign \A[11][97] [3] = 1'b0;
  assign \A[11][97] [2] = 1'b0;
  assign \A[11][97] [0] = 1'b0;
  assign \A[11][98] [0] = 1'b0;
  assign \A[11][100] [4] = 1'b0;
  assign \A[11][100] [3] = 1'b0;
  assign \A[11][100] [2] = 1'b0;
  assign \A[11][101] [1] = 1'b0;
  assign \A[11][102] [0] = 1'b0;
  assign \A[11][106] [4] = 1'b0;
  assign \A[11][106] [3] = 1'b0;
  assign \A[11][106] [2] = 1'b0;
  assign \A[11][106] [1] = 1'b0;
  assign \A[11][106] [0] = 1'b0;
  assign \A[11][107] [1] = 1'b0;
  assign \A[11][108] [4] = 1'b0;
  assign \A[11][108] [3] = 1'b0;
  assign \A[11][108] [2] = 1'b0;
  assign \A[11][108] [0] = 1'b0;
  assign \A[11][109] [4] = 1'b0;
  assign \A[11][109] [3] = 1'b0;
  assign \A[11][109] [2] = 1'b0;
  assign \A[11][109] [1] = 1'b0;
  assign \A[11][109] [0] = 1'b0;
  assign \A[11][110] [0] = 1'b0;
  assign \A[11][111] [4] = 1'b0;
  assign \A[11][111] [3] = 1'b0;
  assign \A[11][111] [2] = 1'b0;
  assign \A[11][111] [1] = 1'b0;
  assign \A[11][111] [0] = 1'b0;
  assign \A[11][112] [4] = 1'b0;
  assign \A[11][112] [3] = 1'b0;
  assign \A[11][112] [2] = 1'b0;
  assign \A[11][112] [1] = 1'b0;
  assign \A[11][113] [4] = 1'b0;
  assign \A[11][113] [3] = 1'b0;
  assign \A[11][113] [2] = 1'b0;
  assign \A[11][113] [1] = 1'b0;
  assign \A[11][113] [0] = 1'b0;
  assign \A[11][114] [4] = 1'b0;
  assign \A[11][114] [3] = 1'b0;
  assign \A[11][114] [2] = 1'b0;
  assign \A[11][114] [1] = 1'b0;
  assign \A[11][115] [4] = 1'b0;
  assign \A[11][115] [3] = 1'b0;
  assign \A[11][115] [2] = 1'b0;
  assign \A[11][115] [0] = 1'b0;
  assign \A[11][116] [4] = 1'b0;
  assign \A[11][116] [3] = 1'b0;
  assign \A[11][116] [2] = 1'b0;
  assign \A[11][116] [1] = 1'b0;
  assign \A[11][117] [4] = 1'b0;
  assign \A[11][117] [3] = 1'b0;
  assign \A[11][117] [2] = 1'b0;
  assign \A[11][117] [1] = 1'b0;
  assign \A[11][119] [4] = 1'b0;
  assign \A[11][119] [3] = 1'b0;
  assign \A[11][119] [2] = 1'b0;
  assign \A[11][119] [1] = 1'b0;
  assign \A[11][119] [0] = 1'b0;
  assign \A[11][120] [4] = 1'b0;
  assign \A[11][120] [3] = 1'b0;
  assign \A[11][120] [2] = 1'b0;
  assign \A[11][120] [1] = 1'b0;
  assign \A[11][122] [4] = 1'b0;
  assign \A[11][122] [3] = 1'b0;
  assign \A[11][122] [2] = 1'b0;
  assign \A[11][122] [1] = 1'b0;
  assign \A[11][124] [4] = 1'b0;
  assign \A[11][124] [3] = 1'b0;
  assign \A[11][124] [1] = 1'b0;
  assign \A[11][124] [0] = 1'b0;
  assign \A[11][125] [4] = 1'b0;
  assign \A[11][125] [3] = 1'b0;
  assign \A[11][125] [2] = 1'b0;
  assign \A[11][125] [1] = 1'b0;
  assign \A[11][125] [0] = 1'b0;
  assign \A[11][126] [1] = 1'b0;
  assign \A[11][127] [0] = 1'b0;
  assign \A[11][128] [4] = 1'b0;
  assign \A[11][128] [3] = 1'b0;
  assign \A[11][128] [2] = 1'b0;
  assign \A[11][129] [4] = 1'b0;
  assign \A[11][129] [3] = 1'b0;
  assign \A[11][129] [1] = 1'b0;
  assign \A[11][129] [0] = 1'b0;
  assign \A[11][130] [4] = 1'b0;
  assign \A[11][130] [3] = 1'b0;
  assign \A[11][130] [2] = 1'b0;
  assign \A[11][130] [1] = 1'b0;
  assign \A[11][130] [0] = 1'b0;
  assign \A[11][132] [4] = 1'b0;
  assign \A[11][132] [3] = 1'b0;
  assign \A[11][132] [2] = 1'b0;
  assign \A[11][132] [1] = 1'b0;
  assign \A[11][134] [4] = 1'b0;
  assign \A[11][134] [3] = 1'b0;
  assign \A[11][134] [2] = 1'b0;
  assign \A[11][134] [1] = 1'b0;
  assign \A[11][135] [4] = 1'b0;
  assign \A[11][135] [3] = 1'b0;
  assign \A[11][135] [2] = 1'b0;
  assign \A[11][135] [1] = 1'b0;
  assign \A[11][135] [0] = 1'b0;
  assign \A[11][136] [4] = 1'b0;
  assign \A[11][136] [3] = 1'b0;
  assign \A[11][136] [2] = 1'b0;
  assign \A[11][136] [0] = 1'b0;
  assign \A[11][137] [4] = 1'b0;
  assign \A[11][137] [3] = 1'b0;
  assign \A[11][137] [2] = 1'b0;
  assign \A[11][137] [0] = 1'b0;
  assign \A[11][139] [4] = 1'b0;
  assign \A[11][139] [3] = 1'b0;
  assign \A[11][139] [2] = 1'b0;
  assign \A[11][139] [1] = 1'b0;
  assign \A[11][140] [0] = 1'b0;
  assign \A[11][141] [4] = 1'b0;
  assign \A[11][141] [3] = 1'b0;
  assign \A[11][141] [2] = 1'b0;
  assign \A[11][142] [4] = 1'b0;
  assign \A[11][142] [3] = 1'b0;
  assign \A[11][142] [2] = 1'b0;
  assign \A[11][142] [0] = 1'b0;
  assign \A[11][143] [4] = 1'b0;
  assign \A[11][143] [3] = 1'b0;
  assign \A[11][143] [2] = 1'b0;
  assign \A[11][143] [0] = 1'b0;
  assign \A[11][144] [4] = 1'b0;
  assign \A[11][144] [3] = 1'b0;
  assign \A[11][144] [2] = 1'b0;
  assign \A[11][144] [1] = 1'b0;
  assign \A[11][144] [0] = 1'b0;
  assign \A[11][145] [4] = 1'b0;
  assign \A[11][145] [3] = 1'b0;
  assign \A[11][145] [2] = 1'b0;
  assign \A[11][146] [4] = 1'b0;
  assign \A[11][146] [3] = 1'b0;
  assign \A[11][146] [1] = 1'b0;
  assign \A[11][147] [4] = 1'b0;
  assign \A[11][147] [3] = 1'b0;
  assign \A[11][147] [2] = 1'b0;
  assign \A[11][147] [0] = 1'b0;
  assign \A[11][148] [4] = 1'b0;
  assign \A[11][148] [3] = 1'b0;
  assign \A[11][148] [2] = 1'b0;
  assign \A[11][148] [1] = 1'b0;
  assign \A[11][150] [0] = 1'b0;
  assign \A[11][151] [4] = 1'b0;
  assign \A[11][151] [3] = 1'b0;
  assign \A[11][151] [2] = 1'b0;
  assign \A[11][151] [0] = 1'b0;
  assign \A[11][152] [4] = 1'b0;
  assign \A[11][152] [3] = 1'b0;
  assign \A[11][152] [2] = 1'b0;
  assign \A[11][152] [1] = 1'b0;
  assign \A[11][153] [0] = 1'b0;
  assign \A[11][154] [4] = 1'b0;
  assign \A[11][154] [3] = 1'b0;
  assign \A[11][154] [2] = 1'b0;
  assign \A[11][154] [1] = 1'b0;
  assign \A[11][154] [0] = 1'b0;
  assign \A[11][155] [4] = 1'b0;
  assign \A[11][155] [3] = 1'b0;
  assign \A[11][155] [2] = 1'b0;
  assign \A[11][155] [0] = 1'b0;
  assign \A[11][157] [4] = 1'b0;
  assign \A[11][157] [3] = 1'b0;
  assign \A[11][157] [2] = 1'b0;
  assign \A[11][157] [0] = 1'b0;
  assign \A[11][159] [4] = 1'b0;
  assign \A[11][159] [3] = 1'b0;
  assign \A[11][159] [2] = 1'b0;
  assign \A[11][159] [1] = 1'b0;
  assign \A[11][161] [4] = 1'b0;
  assign \A[11][161] [3] = 1'b0;
  assign \A[11][162] [4] = 1'b0;
  assign \A[11][162] [3] = 1'b0;
  assign \A[11][162] [2] = 1'b0;
  assign \A[11][162] [1] = 1'b0;
  assign \A[11][163] [4] = 1'b0;
  assign \A[11][163] [3] = 1'b0;
  assign \A[11][163] [2] = 1'b0;
  assign \A[11][163] [0] = 1'b0;
  assign \A[11][164] [0] = 1'b0;
  assign \A[11][167] [4] = 1'b0;
  assign \A[11][167] [3] = 1'b0;
  assign \A[11][167] [2] = 1'b0;
  assign \A[11][168] [4] = 1'b0;
  assign \A[11][168] [3] = 1'b0;
  assign \A[11][168] [2] = 1'b0;
  assign \A[11][169] [4] = 1'b0;
  assign \A[11][169] [3] = 1'b0;
  assign \A[11][169] [2] = 1'b0;
  assign \A[11][169] [1] = 1'b0;
  assign \A[11][170] [4] = 1'b0;
  assign \A[11][170] [3] = 1'b0;
  assign \A[11][170] [1] = 1'b0;
  assign \A[11][170] [0] = 1'b0;
  assign \A[11][171] [4] = 1'b0;
  assign \A[11][171] [3] = 1'b0;
  assign \A[11][171] [2] = 1'b0;
  assign \A[11][171] [1] = 1'b0;
  assign \A[11][172] [4] = 1'b0;
  assign \A[11][172] [3] = 1'b0;
  assign \A[11][172] [2] = 1'b0;
  assign \A[11][172] [1] = 1'b0;
  assign \A[11][173] [4] = 1'b0;
  assign \A[11][173] [3] = 1'b0;
  assign \A[11][173] [2] = 1'b0;
  assign \A[11][173] [0] = 1'b0;
  assign \A[11][174] [4] = 1'b0;
  assign \A[11][174] [3] = 1'b0;
  assign \A[11][174] [2] = 1'b0;
  assign \A[11][174] [0] = 1'b0;
  assign \A[11][175] [4] = 1'b0;
  assign \A[11][175] [3] = 1'b0;
  assign \A[11][175] [2] = 1'b0;
  assign \A[11][175] [0] = 1'b0;
  assign \A[11][176] [4] = 1'b0;
  assign \A[11][176] [3] = 1'b0;
  assign \A[11][176] [2] = 1'b0;
  assign \A[11][176] [0] = 1'b0;
  assign \A[11][177] [4] = 1'b0;
  assign \A[11][177] [3] = 1'b0;
  assign \A[11][177] [2] = 1'b0;
  assign \A[11][177] [0] = 1'b0;
  assign \A[11][178] [4] = 1'b0;
  assign \A[11][178] [3] = 1'b0;
  assign \A[11][178] [2] = 1'b0;
  assign \A[11][178] [1] = 1'b0;
  assign \A[11][178] [0] = 1'b0;
  assign \A[11][179] [4] = 1'b0;
  assign \A[11][179] [3] = 1'b0;
  assign \A[11][179] [2] = 1'b0;
  assign \A[11][179] [1] = 1'b0;
  assign \A[11][180] [4] = 1'b0;
  assign \A[11][180] [3] = 1'b0;
  assign \A[11][180] [2] = 1'b0;
  assign \A[11][180] [0] = 1'b0;
  assign \A[11][181] [4] = 1'b0;
  assign \A[11][181] [3] = 1'b0;
  assign \A[11][181] [2] = 1'b0;
  assign \A[11][181] [1] = 1'b0;
  assign \A[11][183] [4] = 1'b0;
  assign \A[11][183] [3] = 1'b0;
  assign \A[11][183] [2] = 1'b0;
  assign \A[11][183] [1] = 1'b0;
  assign \A[11][184] [4] = 1'b0;
  assign \A[11][184] [3] = 1'b0;
  assign \A[11][184] [2] = 1'b0;
  assign \A[11][184] [1] = 1'b0;
  assign \A[11][184] [0] = 1'b0;
  assign \A[11][185] [4] = 1'b0;
  assign \A[11][185] [3] = 1'b0;
  assign \A[11][185] [2] = 1'b0;
  assign \A[11][185] [0] = 1'b0;
  assign \A[11][186] [4] = 1'b0;
  assign \A[11][186] [3] = 1'b0;
  assign \A[11][186] [2] = 1'b0;
  assign \A[11][186] [1] = 1'b0;
  assign \A[11][186] [0] = 1'b0;
  assign \A[11][187] [4] = 1'b0;
  assign \A[11][187] [3] = 1'b0;
  assign \A[11][187] [2] = 1'b0;
  assign \A[11][187] [0] = 1'b0;
  assign \A[11][189] [4] = 1'b0;
  assign \A[11][189] [3] = 1'b0;
  assign \A[11][189] [2] = 1'b0;
  assign \A[11][189] [0] = 1'b0;
  assign \A[11][190] [4] = 1'b0;
  assign \A[11][190] [3] = 1'b0;
  assign \A[11][190] [2] = 1'b0;
  assign \A[11][190] [1] = 1'b0;
  assign \A[11][191] [4] = 1'b0;
  assign \A[11][191] [3] = 1'b0;
  assign \A[11][191] [2] = 1'b0;
  assign \A[11][191] [1] = 1'b0;
  assign \A[11][191] [0] = 1'b0;
  assign \A[11][192] [4] = 1'b0;
  assign \A[11][192] [3] = 1'b0;
  assign \A[11][192] [2] = 1'b0;
  assign \A[11][192] [1] = 1'b0;
  assign \A[11][192] [0] = 1'b0;
  assign \A[11][193] [4] = 1'b0;
  assign \A[11][193] [3] = 1'b0;
  assign \A[11][193] [2] = 1'b0;
  assign \A[11][193] [1] = 1'b0;
  assign \A[11][194] [4] = 1'b0;
  assign \A[11][194] [3] = 1'b0;
  assign \A[11][194] [2] = 1'b0;
  assign \A[11][195] [4] = 1'b0;
  assign \A[11][195] [3] = 1'b0;
  assign \A[11][195] [2] = 1'b0;
  assign \A[11][195] [1] = 1'b0;
  assign \A[11][196] [4] = 1'b0;
  assign \A[11][196] [3] = 1'b0;
  assign \A[11][196] [2] = 1'b0;
  assign \A[11][196] [1] = 1'b0;
  assign \A[11][197] [4] = 1'b0;
  assign \A[11][197] [3] = 1'b0;
  assign \A[11][197] [2] = 1'b0;
  assign \A[11][197] [0] = 1'b0;
  assign \A[11][198] [0] = 1'b0;
  assign \A[11][199] [4] = 1'b0;
  assign \A[11][199] [3] = 1'b0;
  assign \A[11][199] [2] = 1'b0;
  assign \A[11][200] [0] = 1'b0;
  assign \A[11][201] [4] = 1'b0;
  assign \A[11][201] [3] = 1'b0;
  assign \A[11][201] [2] = 1'b0;
  assign \A[11][201] [1] = 1'b0;
  assign \A[11][201] [0] = 1'b0;
  assign \A[11][202] [4] = 1'b0;
  assign \A[11][202] [3] = 1'b0;
  assign \A[11][202] [2] = 1'b0;
  assign \A[11][202] [0] = 1'b0;
  assign \A[11][203] [4] = 1'b0;
  assign \A[11][203] [3] = 1'b0;
  assign \A[11][203] [2] = 1'b0;
  assign \A[11][203] [1] = 1'b0;
  assign \A[11][203] [0] = 1'b0;
  assign \A[11][204] [4] = 1'b0;
  assign \A[11][204] [3] = 1'b0;
  assign \A[11][204] [2] = 1'b0;
  assign \A[11][204] [1] = 1'b0;
  assign \A[11][204] [0] = 1'b0;
  assign \A[11][206] [4] = 1'b0;
  assign \A[11][206] [3] = 1'b0;
  assign \A[11][206] [2] = 1'b0;
  assign \A[11][206] [1] = 1'b0;
  assign \A[11][206] [0] = 1'b0;
  assign \A[11][207] [4] = 1'b0;
  assign \A[11][207] [3] = 1'b0;
  assign \A[11][207] [2] = 1'b0;
  assign \A[11][207] [1] = 1'b0;
  assign \A[11][208] [4] = 1'b0;
  assign \A[11][208] [3] = 1'b0;
  assign \A[11][208] [2] = 1'b0;
  assign \A[11][208] [1] = 1'b0;
  assign \A[11][211] [4] = 1'b0;
  assign \A[11][211] [3] = 1'b0;
  assign \A[11][211] [2] = 1'b0;
  assign \A[11][211] [1] = 1'b0;
  assign \A[11][212] [1] = 1'b0;
  assign \A[11][212] [0] = 1'b0;
  assign \A[11][214] [4] = 1'b0;
  assign \A[11][214] [3] = 1'b0;
  assign \A[11][214] [2] = 1'b0;
  assign \A[11][214] [1] = 1'b0;
  assign \A[11][214] [0] = 1'b0;
  assign \A[11][215] [4] = 1'b0;
  assign \A[11][215] [3] = 1'b0;
  assign \A[11][215] [2] = 1'b0;
  assign \A[11][215] [1] = 1'b0;
  assign \A[11][217] [4] = 1'b0;
  assign \A[11][217] [3] = 1'b0;
  assign \A[11][217] [2] = 1'b0;
  assign \A[11][217] [1] = 1'b0;
  assign \A[11][218] [0] = 1'b0;
  assign \A[11][219] [4] = 1'b0;
  assign \A[11][219] [3] = 1'b0;
  assign \A[11][219] [2] = 1'b0;
  assign \A[11][219] [1] = 1'b0;
  assign \A[11][219] [0] = 1'b0;
  assign \A[11][221] [4] = 1'b0;
  assign \A[11][221] [3] = 1'b0;
  assign \A[11][221] [2] = 1'b0;
  assign \A[11][221] [1] = 1'b0;
  assign \A[11][222] [1] = 1'b0;
  assign \A[11][224] [4] = 1'b0;
  assign \A[11][224] [3] = 1'b0;
  assign \A[11][224] [2] = 1'b0;
  assign \A[11][224] [1] = 1'b0;
  assign \A[11][225] [4] = 1'b0;
  assign \A[11][225] [3] = 1'b0;
  assign \A[11][225] [2] = 1'b0;
  assign \A[11][225] [1] = 1'b0;
  assign \A[11][226] [0] = 1'b0;
  assign \A[11][228] [4] = 1'b0;
  assign \A[11][228] [3] = 1'b0;
  assign \A[11][228] [2] = 1'b0;
  assign \A[11][228] [1] = 1'b0;
  assign \A[11][228] [0] = 1'b0;
  assign \A[11][229] [4] = 1'b0;
  assign \A[11][229] [3] = 1'b0;
  assign \A[11][229] [2] = 1'b0;
  assign \A[11][230] [0] = 1'b0;
  assign \A[11][231] [4] = 1'b0;
  assign \A[11][231] [3] = 1'b0;
  assign \A[11][231] [2] = 1'b0;
  assign \A[11][231] [1] = 1'b0;
  assign \A[11][231] [0] = 1'b0;
  assign \A[11][232] [4] = 1'b0;
  assign \A[11][232] [3] = 1'b0;
  assign \A[11][232] [2] = 1'b0;
  assign \A[11][232] [1] = 1'b0;
  assign \A[11][232] [0] = 1'b0;
  assign \A[11][234] [4] = 1'b0;
  assign \A[11][234] [3] = 1'b0;
  assign \A[11][234] [2] = 1'b0;
  assign \A[11][234] [1] = 1'b0;
  assign \A[11][234] [0] = 1'b0;
  assign \A[11][235] [4] = 1'b0;
  assign \A[11][235] [3] = 1'b0;
  assign \A[11][235] [2] = 1'b0;
  assign \A[11][235] [1] = 1'b0;
  assign \A[11][236] [4] = 1'b0;
  assign \A[11][236] [3] = 1'b0;
  assign \A[11][236] [2] = 1'b0;
  assign \A[11][236] [1] = 1'b0;
  assign \A[11][236] [0] = 1'b0;
  assign \A[11][237] [4] = 1'b0;
  assign \A[11][237] [3] = 1'b0;
  assign \A[11][237] [2] = 1'b0;
  assign \A[11][237] [1] = 1'b0;
  assign \A[11][237] [0] = 1'b0;
  assign \A[11][239] [0] = 1'b0;
  assign \A[11][242] [4] = 1'b0;
  assign \A[11][242] [3] = 1'b0;
  assign \A[11][242] [2] = 1'b0;
  assign \A[11][242] [1] = 1'b0;
  assign \A[11][244] [1] = 1'b0;
  assign \A[11][247] [4] = 1'b0;
  assign \A[11][247] [3] = 1'b0;
  assign \A[11][247] [2] = 1'b0;
  assign \A[11][247] [1] = 1'b0;
  assign \A[11][248] [4] = 1'b0;
  assign \A[11][248] [3] = 1'b0;
  assign \A[11][248] [2] = 1'b0;
  assign \A[11][248] [1] = 1'b0;
  assign \A[11][248] [0] = 1'b0;
  assign \A[11][249] [4] = 1'b0;
  assign \A[11][249] [3] = 1'b0;
  assign \A[11][249] [2] = 1'b0;
  assign \A[11][249] [1] = 1'b0;
  assign \A[11][249] [0] = 1'b0;
  assign \A[11][250] [4] = 1'b0;
  assign \A[11][250] [3] = 1'b0;
  assign \A[11][250] [2] = 1'b0;
  assign \A[11][250] [1] = 1'b0;
  assign \A[11][250] [0] = 1'b0;
  assign \A[11][251] [0] = 1'b0;
  assign \A[11][253] [4] = 1'b0;
  assign \A[11][253] [3] = 1'b0;
  assign \A[11][253] [2] = 1'b0;
  assign \A[11][253] [1] = 1'b0;
  assign \A[11][253] [0] = 1'b0;
  assign \A[11][254] [0] = 1'b0;
  assign \A[12][0] [4] = 1'b0;
  assign \A[12][0] [3] = 1'b0;
  assign \A[12][0] [2] = 1'b0;
  assign \A[12][0] [1] = 1'b0;
  assign \A[12][1] [0] = 1'b0;
  assign \A[12][2] [0] = 1'b0;
  assign \A[12][3] [4] = 1'b0;
  assign \A[12][3] [3] = 1'b0;
  assign \A[12][3] [2] = 1'b0;
  assign \A[12][3] [1] = 1'b0;
  assign \A[12][3] [0] = 1'b0;
  assign \A[12][4] [4] = 1'b0;
  assign \A[12][4] [3] = 1'b0;
  assign \A[12][4] [2] = 1'b0;
  assign \A[12][4] [1] = 1'b0;
  assign \A[12][5] [4] = 1'b0;
  assign \A[12][5] [3] = 1'b0;
  assign \A[12][5] [2] = 1'b0;
  assign \A[12][5] [0] = 1'b0;
  assign \A[12][6] [0] = 1'b0;
  assign \A[12][7] [4] = 1'b0;
  assign \A[12][7] [3] = 1'b0;
  assign \A[12][7] [2] = 1'b0;
  assign \A[12][7] [1] = 1'b0;
  assign \A[12][7] [0] = 1'b0;
  assign \A[12][8] [1] = 1'b0;
  assign \A[12][10] [0] = 1'b0;
  assign \A[12][12] [4] = 1'b0;
  assign \A[12][12] [3] = 1'b0;
  assign \A[12][12] [2] = 1'b0;
  assign \A[12][12] [1] = 1'b0;
  assign \A[12][12] [0] = 1'b0;
  assign \A[12][13] [4] = 1'b0;
  assign \A[12][13] [3] = 1'b0;
  assign \A[12][13] [2] = 1'b0;
  assign \A[12][13] [0] = 1'b0;
  assign \A[12][14] [4] = 1'b0;
  assign \A[12][14] [3] = 1'b0;
  assign \A[12][14] [2] = 1'b0;
  assign \A[12][14] [1] = 1'b0;
  assign \A[12][19] [4] = 1'b0;
  assign \A[12][19] [3] = 1'b0;
  assign \A[12][19] [2] = 1'b0;
  assign \A[12][19] [1] = 1'b0;
  assign \A[12][19] [0] = 1'b0;
  assign \A[12][20] [4] = 1'b0;
  assign \A[12][20] [3] = 1'b0;
  assign \A[12][20] [2] = 1'b0;
  assign \A[12][20] [1] = 1'b0;
  assign \A[12][20] [0] = 1'b0;
  assign \A[12][21] [4] = 1'b0;
  assign \A[12][21] [3] = 1'b0;
  assign \A[12][21] [2] = 1'b0;
  assign \A[12][21] [1] = 1'b0;
  assign \A[12][23] [4] = 1'b0;
  assign \A[12][23] [3] = 1'b0;
  assign \A[12][23] [2] = 1'b0;
  assign \A[12][23] [1] = 1'b0;
  assign \A[12][24] [4] = 1'b0;
  assign \A[12][24] [3] = 1'b0;
  assign \A[12][24] [2] = 1'b0;
  assign \A[12][24] [1] = 1'b0;
  assign \A[12][24] [0] = 1'b0;
  assign \A[12][27] [4] = 1'b0;
  assign \A[12][27] [3] = 1'b0;
  assign \A[12][27] [2] = 1'b0;
  assign \A[12][27] [1] = 1'b0;
  assign \A[12][28] [4] = 1'b0;
  assign \A[12][28] [3] = 1'b0;
  assign \A[12][28] [2] = 1'b0;
  assign \A[12][28] [1] = 1'b0;
  assign \A[12][28] [0] = 1'b0;
  assign \A[12][29] [4] = 1'b0;
  assign \A[12][29] [3] = 1'b0;
  assign \A[12][29] [2] = 1'b0;
  assign \A[12][29] [1] = 1'b0;
  assign \A[12][30] [0] = 1'b0;
  assign \A[12][31] [0] = 1'b0;
  assign \A[12][32] [4] = 1'b0;
  assign \A[12][32] [3] = 1'b0;
  assign \A[12][32] [2] = 1'b0;
  assign \A[12][32] [1] = 1'b0;
  assign \A[12][33] [4] = 1'b0;
  assign \A[12][33] [3] = 1'b0;
  assign \A[12][33] [2] = 1'b0;
  assign \A[12][33] [1] = 1'b0;
  assign \A[12][34] [4] = 1'b0;
  assign \A[12][34] [3] = 1'b0;
  assign \A[12][34] [2] = 1'b0;
  assign \A[12][34] [1] = 1'b0;
  assign \A[12][34] [0] = 1'b0;
  assign \A[12][35] [4] = 1'b0;
  assign \A[12][35] [3] = 1'b0;
  assign \A[12][35] [2] = 1'b0;
  assign \A[12][35] [1] = 1'b0;
  assign \A[12][35] [0] = 1'b0;
  assign \A[12][36] [4] = 1'b0;
  assign \A[12][36] [3] = 1'b0;
  assign \A[12][36] [2] = 1'b0;
  assign \A[12][36] [1] = 1'b0;
  assign \A[12][36] [0] = 1'b0;
  assign \A[12][37] [4] = 1'b0;
  assign \A[12][37] [3] = 1'b0;
  assign \A[12][37] [2] = 1'b0;
  assign \A[12][37] [1] = 1'b0;
  assign \A[12][38] [4] = 1'b0;
  assign \A[12][38] [3] = 1'b0;
  assign \A[12][38] [2] = 1'b0;
  assign \A[12][38] [1] = 1'b0;
  assign \A[12][38] [0] = 1'b0;
  assign \A[12][41] [4] = 1'b0;
  assign \A[12][41] [3] = 1'b0;
  assign \A[12][41] [2] = 1'b0;
  assign \A[12][41] [1] = 1'b0;
  assign \A[12][42] [4] = 1'b0;
  assign \A[12][42] [3] = 1'b0;
  assign \A[12][42] [2] = 1'b0;
  assign \A[12][42] [1] = 1'b0;
  assign \A[12][43] [4] = 1'b0;
  assign \A[12][43] [3] = 1'b0;
  assign \A[12][43] [2] = 1'b0;
  assign \A[12][43] [1] = 1'b0;
  assign \A[12][45] [4] = 1'b0;
  assign \A[12][45] [3] = 1'b0;
  assign \A[12][45] [2] = 1'b0;
  assign \A[12][45] [1] = 1'b0;
  assign \A[12][45] [0] = 1'b0;
  assign \A[12][46] [4] = 1'b0;
  assign \A[12][46] [3] = 1'b0;
  assign \A[12][46] [2] = 1'b0;
  assign \A[12][46] [0] = 1'b0;
  assign \A[12][49] [4] = 1'b0;
  assign \A[12][49] [3] = 1'b0;
  assign \A[12][49] [2] = 1'b0;
  assign \A[12][49] [1] = 1'b0;
  assign \A[12][50] [1] = 1'b0;
  assign \A[12][51] [0] = 1'b0;
  assign \A[12][52] [4] = 1'b0;
  assign \A[12][52] [3] = 1'b0;
  assign \A[12][52] [2] = 1'b0;
  assign \A[12][52] [1] = 1'b0;
  assign \A[12][53] [4] = 1'b0;
  assign \A[12][53] [3] = 1'b0;
  assign \A[12][53] [2] = 1'b0;
  assign \A[12][54] [0] = 1'b0;
  assign \A[12][55] [4] = 1'b0;
  assign \A[12][55] [3] = 1'b0;
  assign \A[12][55] [2] = 1'b0;
  assign \A[12][55] [1] = 1'b0;
  assign \A[12][56] [4] = 1'b0;
  assign \A[12][56] [3] = 1'b0;
  assign \A[12][56] [2] = 1'b0;
  assign \A[12][56] [0] = 1'b0;
  assign \A[12][57] [4] = 1'b0;
  assign \A[12][57] [3] = 1'b0;
  assign \A[12][57] [2] = 1'b0;
  assign \A[12][57] [1] = 1'b0;
  assign \A[12][57] [0] = 1'b0;
  assign \A[12][58] [4] = 1'b0;
  assign \A[12][58] [3] = 1'b0;
  assign \A[12][58] [2] = 1'b0;
  assign \A[12][58] [1] = 1'b0;
  assign \A[12][61] [4] = 1'b0;
  assign \A[12][61] [3] = 1'b0;
  assign \A[12][61] [2] = 1'b0;
  assign \A[12][61] [1] = 1'b0;
  assign \A[12][61] [0] = 1'b0;
  assign \A[12][62] [4] = 1'b0;
  assign \A[12][62] [3] = 1'b0;
  assign \A[12][62] [2] = 1'b0;
  assign \A[12][62] [0] = 1'b0;
  assign \A[12][63] [4] = 1'b0;
  assign \A[12][63] [3] = 1'b0;
  assign \A[12][63] [2] = 1'b0;
  assign \A[12][63] [1] = 1'b0;
  assign \A[12][64] [4] = 1'b0;
  assign \A[12][64] [3] = 1'b0;
  assign \A[12][64] [2] = 1'b0;
  assign \A[12][65] [4] = 1'b0;
  assign \A[12][65] [3] = 1'b0;
  assign \A[12][65] [2] = 1'b0;
  assign \A[12][65] [1] = 1'b0;
  assign \A[12][65] [0] = 1'b0;
  assign \A[12][66] [4] = 1'b0;
  assign \A[12][66] [3] = 1'b0;
  assign \A[12][66] [2] = 1'b0;
  assign \A[12][66] [1] = 1'b0;
  assign \A[12][67] [4] = 1'b0;
  assign \A[12][67] [3] = 1'b0;
  assign \A[12][67] [2] = 1'b0;
  assign \A[12][67] [1] = 1'b0;
  assign \A[12][67] [0] = 1'b0;
  assign \A[12][68] [4] = 1'b0;
  assign \A[12][68] [3] = 1'b0;
  assign \A[12][68] [2] = 1'b0;
  assign \A[12][68] [1] = 1'b0;
  assign \A[12][69] [4] = 1'b0;
  assign \A[12][69] [3] = 1'b0;
  assign \A[12][69] [2] = 1'b0;
  assign \A[12][70] [0] = 1'b0;
  assign \A[12][71] [1] = 1'b0;
  assign \A[12][72] [4] = 1'b0;
  assign \A[12][72] [3] = 1'b0;
  assign \A[12][72] [2] = 1'b0;
  assign \A[12][72] [1] = 1'b0;
  assign \A[12][73] [4] = 1'b0;
  assign \A[12][73] [3] = 1'b0;
  assign \A[12][73] [2] = 1'b0;
  assign \A[12][73] [1] = 1'b0;
  assign \A[12][73] [0] = 1'b0;
  assign \A[12][74] [1] = 1'b0;
  assign \A[12][77] [4] = 1'b0;
  assign \A[12][77] [3] = 1'b0;
  assign \A[12][77] [2] = 1'b0;
  assign \A[12][77] [1] = 1'b0;
  assign \A[12][78] [0] = 1'b0;
  assign \A[12][80] [4] = 1'b0;
  assign \A[12][80] [3] = 1'b0;
  assign \A[12][80] [2] = 1'b0;
  assign \A[12][80] [1] = 1'b0;
  assign \A[12][81] [0] = 1'b0;
  assign \A[12][83] [0] = 1'b0;
  assign \A[12][84] [4] = 1'b0;
  assign \A[12][84] [3] = 1'b0;
  assign \A[12][84] [2] = 1'b0;
  assign \A[12][85] [4] = 1'b0;
  assign \A[12][85] [3] = 1'b0;
  assign \A[12][85] [2] = 1'b0;
  assign \A[12][85] [0] = 1'b0;
  assign \A[12][86] [4] = 1'b0;
  assign \A[12][86] [3] = 1'b0;
  assign \A[12][86] [2] = 1'b0;
  assign \A[12][86] [1] = 1'b0;
  assign \A[12][88] [4] = 1'b0;
  assign \A[12][88] [3] = 1'b0;
  assign \A[12][88] [2] = 1'b0;
  assign \A[12][88] [1] = 1'b0;
  assign \A[12][89] [4] = 1'b0;
  assign \A[12][89] [3] = 1'b0;
  assign \A[12][89] [2] = 1'b0;
  assign \A[12][89] [1] = 1'b0;
  assign \A[12][89] [0] = 1'b0;
  assign \A[12][90] [4] = 1'b0;
  assign \A[12][90] [3] = 1'b0;
  assign \A[12][90] [2] = 1'b0;
  assign \A[12][90] [1] = 1'b0;
  assign \A[12][92] [0] = 1'b0;
  assign \A[12][94] [4] = 1'b0;
  assign \A[12][94] [3] = 1'b0;
  assign \A[12][94] [2] = 1'b0;
  assign \A[12][94] [1] = 1'b0;
  assign \A[12][97] [4] = 1'b0;
  assign \A[12][97] [3] = 1'b0;
  assign \A[12][97] [2] = 1'b0;
  assign \A[12][97] [1] = 1'b0;
  assign \A[12][97] [0] = 1'b0;
  assign \A[12][99] [4] = 1'b0;
  assign \A[12][99] [3] = 1'b0;
  assign \A[12][99] [2] = 1'b0;
  assign \A[12][99] [1] = 1'b0;
  assign \A[12][99] [0] = 1'b0;
  assign \A[12][100] [0] = 1'b0;
  assign \A[12][102] [4] = 1'b0;
  assign \A[12][102] [3] = 1'b0;
  assign \A[12][102] [2] = 1'b0;
  assign \A[12][102] [1] = 1'b0;
  assign \A[12][103] [4] = 1'b0;
  assign \A[12][103] [3] = 1'b0;
  assign \A[12][103] [2] = 1'b0;
  assign \A[12][103] [1] = 1'b0;
  assign \A[12][103] [0] = 1'b0;
  assign \A[12][104] [4] = 1'b0;
  assign \A[12][104] [3] = 1'b0;
  assign \A[12][104] [2] = 1'b0;
  assign \A[12][104] [1] = 1'b0;
  assign \A[12][105] [4] = 1'b0;
  assign \A[12][105] [3] = 1'b0;
  assign \A[12][105] [2] = 1'b0;
  assign \A[12][105] [0] = 1'b0;
  assign \A[12][106] [0] = 1'b0;
  assign \A[12][107] [4] = 1'b0;
  assign \A[12][107] [3] = 1'b0;
  assign \A[12][107] [2] = 1'b0;
  assign \A[12][107] [1] = 1'b0;
  assign \A[12][107] [0] = 1'b0;
  assign \A[12][108] [4] = 1'b0;
  assign \A[12][108] [3] = 1'b0;
  assign \A[12][108] [2] = 1'b0;
  assign \A[12][108] [1] = 1'b0;
  assign \A[12][109] [4] = 1'b0;
  assign \A[12][109] [3] = 1'b0;
  assign \A[12][109] [2] = 1'b0;
  assign \A[12][109] [1] = 1'b0;
  assign \A[12][109] [0] = 1'b0;
  assign \A[12][110] [4] = 1'b0;
  assign \A[12][110] [3] = 1'b0;
  assign \A[12][110] [2] = 1'b0;
  assign \A[12][110] [1] = 1'b0;
  assign \A[12][111] [4] = 1'b0;
  assign \A[12][111] [3] = 1'b0;
  assign \A[12][111] [2] = 1'b0;
  assign \A[12][111] [0] = 1'b0;
  assign \A[12][112] [4] = 1'b0;
  assign \A[12][112] [3] = 1'b0;
  assign \A[12][112] [2] = 1'b0;
  assign \A[12][112] [1] = 1'b0;
  assign \A[12][113] [4] = 1'b0;
  assign \A[12][113] [3] = 1'b0;
  assign \A[12][113] [2] = 1'b0;
  assign \A[12][113] [0] = 1'b0;
  assign \A[12][114] [4] = 1'b0;
  assign \A[12][114] [3] = 1'b0;
  assign \A[12][114] [2] = 1'b0;
  assign \A[12][114] [0] = 1'b0;
  assign \A[12][115] [0] = 1'b0;
  assign \A[12][116] [1] = 1'b0;
  assign \A[12][117] [4] = 1'b0;
  assign \A[12][117] [3] = 1'b0;
  assign \A[12][117] [2] = 1'b0;
  assign \A[12][117] [1] = 1'b0;
  assign \A[12][119] [4] = 1'b0;
  assign \A[12][119] [3] = 1'b0;
  assign \A[12][119] [2] = 1'b0;
  assign \A[12][119] [1] = 1'b0;
  assign \A[12][119] [0] = 1'b0;
  assign \A[12][120] [4] = 1'b0;
  assign \A[12][120] [3] = 1'b0;
  assign \A[12][120] [2] = 1'b0;
  assign \A[12][120] [0] = 1'b0;
  assign \A[12][121] [4] = 1'b0;
  assign \A[12][121] [3] = 1'b0;
  assign \A[12][121] [2] = 1'b0;
  assign \A[12][121] [1] = 1'b0;
  assign \A[12][122] [1] = 1'b0;
  assign \A[12][124] [0] = 1'b0;
  assign \A[12][125] [0] = 1'b0;
  assign \A[12][126] [4] = 1'b0;
  assign \A[12][126] [3] = 1'b0;
  assign \A[12][126] [2] = 1'b0;
  assign \A[12][126] [0] = 1'b0;
  assign \A[12][127] [0] = 1'b0;
  assign \A[12][128] [1] = 1'b0;
  assign \A[12][129] [0] = 1'b0;
  assign \A[12][132] [0] = 1'b0;
  assign \A[12][133] [4] = 1'b0;
  assign \A[12][133] [3] = 1'b0;
  assign \A[12][133] [2] = 1'b0;
  assign \A[12][133] [1] = 1'b0;
  assign \A[12][133] [0] = 1'b0;
  assign \A[12][134] [4] = 1'b0;
  assign \A[12][134] [3] = 1'b0;
  assign \A[12][134] [2] = 1'b0;
  assign \A[12][135] [4] = 1'b0;
  assign \A[12][135] [3] = 1'b0;
  assign \A[12][135] [2] = 1'b0;
  assign \A[12][135] [0] = 1'b0;
  assign \A[12][136] [4] = 1'b0;
  assign \A[12][136] [3] = 1'b0;
  assign \A[12][136] [2] = 1'b0;
  assign \A[12][136] [1] = 1'b0;
  assign \A[12][136] [0] = 1'b0;
  assign \A[12][137] [4] = 1'b0;
  assign \A[12][137] [3] = 1'b0;
  assign \A[12][137] [2] = 1'b0;
  assign \A[12][137] [1] = 1'b0;
  assign \A[12][137] [0] = 1'b0;
  assign \A[12][138] [4] = 1'b0;
  assign \A[12][138] [3] = 1'b0;
  assign \A[12][138] [2] = 1'b0;
  assign \A[12][138] [1] = 1'b0;
  assign \A[12][138] [0] = 1'b0;
  assign \A[12][139] [4] = 1'b0;
  assign \A[12][139] [3] = 1'b0;
  assign \A[12][139] [2] = 1'b0;
  assign \A[12][139] [1] = 1'b0;
  assign \A[12][139] [0] = 1'b0;
  assign \A[12][140] [4] = 1'b0;
  assign \A[12][140] [3] = 1'b0;
  assign \A[12][140] [2] = 1'b0;
  assign \A[12][141] [4] = 1'b0;
  assign \A[12][141] [3] = 1'b0;
  assign \A[12][141] [2] = 1'b0;
  assign \A[12][142] [4] = 1'b0;
  assign \A[12][142] [3] = 1'b0;
  assign \A[12][142] [2] = 1'b0;
  assign \A[12][142] [1] = 1'b0;
  assign \A[12][143] [4] = 1'b0;
  assign \A[12][143] [3] = 1'b0;
  assign \A[12][143] [2] = 1'b0;
  assign \A[12][143] [0] = 1'b0;
  assign \A[12][144] [4] = 1'b0;
  assign \A[12][144] [3] = 1'b0;
  assign \A[12][144] [2] = 1'b0;
  assign \A[12][144] [1] = 1'b0;
  assign \A[12][145] [4] = 1'b0;
  assign \A[12][145] [3] = 1'b0;
  assign \A[12][145] [2] = 1'b0;
  assign \A[12][145] [1] = 1'b0;
  assign \A[12][145] [0] = 1'b0;
  assign \A[12][146] [4] = 1'b0;
  assign \A[12][146] [3] = 1'b0;
  assign \A[12][146] [2] = 1'b0;
  assign \A[12][146] [1] = 1'b0;
  assign \A[12][147] [4] = 1'b0;
  assign \A[12][147] [3] = 1'b0;
  assign \A[12][147] [2] = 1'b0;
  assign \A[12][147] [1] = 1'b0;
  assign \A[12][149] [4] = 1'b0;
  assign \A[12][149] [3] = 1'b0;
  assign \A[12][149] [2] = 1'b0;
  assign \A[12][149] [1] = 1'b0;
  assign \A[12][149] [0] = 1'b0;
  assign \A[12][150] [4] = 1'b0;
  assign \A[12][150] [3] = 1'b0;
  assign \A[12][150] [1] = 1'b0;
  assign \A[12][150] [0] = 1'b0;
  assign \A[12][151] [4] = 1'b0;
  assign \A[12][151] [3] = 1'b0;
  assign \A[12][151] [2] = 1'b0;
  assign \A[12][153] [4] = 1'b0;
  assign \A[12][153] [3] = 1'b0;
  assign \A[12][153] [2] = 1'b0;
  assign \A[12][153] [0] = 1'b0;
  assign \A[12][154] [4] = 1'b0;
  assign \A[12][154] [3] = 1'b0;
  assign \A[12][154] [2] = 1'b0;
  assign \A[12][154] [0] = 1'b0;
  assign \A[12][155] [1] = 1'b0;
  assign \A[12][156] [4] = 1'b0;
  assign \A[12][156] [3] = 1'b0;
  assign \A[12][156] [2] = 1'b0;
  assign \A[12][156] [1] = 1'b0;
  assign \A[12][157] [4] = 1'b0;
  assign \A[12][157] [3] = 1'b0;
  assign \A[12][157] [2] = 1'b0;
  assign \A[12][157] [1] = 1'b0;
  assign \A[12][157] [0] = 1'b0;
  assign \A[12][158] [0] = 1'b0;
  assign \A[12][159] [4] = 1'b0;
  assign \A[12][159] [3] = 1'b0;
  assign \A[12][159] [2] = 1'b0;
  assign \A[12][159] [1] = 1'b0;
  assign \A[12][159] [0] = 1'b0;
  assign \A[12][160] [4] = 1'b0;
  assign \A[12][160] [3] = 1'b0;
  assign \A[12][160] [2] = 1'b0;
  assign \A[12][160] [1] = 1'b0;
  assign \A[12][161] [4] = 1'b0;
  assign \A[12][161] [3] = 1'b0;
  assign \A[12][161] [2] = 1'b0;
  assign \A[12][161] [1] = 1'b0;
  assign \A[12][161] [0] = 1'b0;
  assign \A[12][162] [4] = 1'b0;
  assign \A[12][162] [3] = 1'b0;
  assign \A[12][162] [2] = 1'b0;
  assign \A[12][162] [1] = 1'b0;
  assign \A[12][162] [0] = 1'b0;
  assign \A[12][163] [0] = 1'b0;
  assign \A[12][164] [4] = 1'b0;
  assign \A[12][164] [3] = 1'b0;
  assign \A[12][164] [2] = 1'b0;
  assign \A[12][164] [0] = 1'b0;
  assign \A[12][165] [4] = 1'b0;
  assign \A[12][165] [3] = 1'b0;
  assign \A[12][165] [2] = 1'b0;
  assign \A[12][165] [0] = 1'b0;
  assign \A[12][166] [4] = 1'b0;
  assign \A[12][166] [3] = 1'b0;
  assign \A[12][166] [2] = 1'b0;
  assign \A[12][166] [1] = 1'b0;
  assign \A[12][166] [0] = 1'b0;
  assign \A[12][167] [4] = 1'b0;
  assign \A[12][167] [3] = 1'b0;
  assign \A[12][167] [2] = 1'b0;
  assign \A[12][167] [0] = 1'b0;
  assign \A[12][168] [4] = 1'b0;
  assign \A[12][168] [3] = 1'b0;
  assign \A[12][168] [2] = 1'b0;
  assign \A[12][168] [1] = 1'b0;
  assign \A[12][169] [4] = 1'b0;
  assign \A[12][169] [3] = 1'b0;
  assign \A[12][169] [2] = 1'b0;
  assign \A[12][169] [1] = 1'b0;
  assign \A[12][169] [0] = 1'b0;
  assign \A[12][170] [4] = 1'b0;
  assign \A[12][170] [3] = 1'b0;
  assign \A[12][170] [2] = 1'b0;
  assign \A[12][170] [0] = 1'b0;
  assign \A[12][171] [4] = 1'b0;
  assign \A[12][171] [3] = 1'b0;
  assign \A[12][171] [2] = 1'b0;
  assign \A[12][171] [1] = 1'b0;
  assign \A[12][171] [0] = 1'b0;
  assign \A[12][174] [4] = 1'b0;
  assign \A[12][174] [3] = 1'b0;
  assign \A[12][174] [2] = 1'b0;
  assign \A[12][174] [1] = 1'b0;
  assign \A[12][174] [0] = 1'b0;
  assign \A[12][175] [4] = 1'b0;
  assign \A[12][175] [3] = 1'b0;
  assign \A[12][175] [2] = 1'b0;
  assign \A[12][175] [1] = 1'b0;
  assign \A[12][175] [0] = 1'b0;
  assign \A[12][176] [0] = 1'b0;
  assign \A[12][178] [4] = 1'b0;
  assign \A[12][178] [3] = 1'b0;
  assign \A[12][178] [2] = 1'b0;
  assign \A[12][178] [1] = 1'b0;
  assign \A[12][179] [0] = 1'b0;
  assign \A[12][182] [4] = 1'b0;
  assign \A[12][182] [3] = 1'b0;
  assign \A[12][182] [2] = 1'b0;
  assign \A[12][182] [1] = 1'b0;
  assign \A[12][182] [0] = 1'b0;
  assign \A[12][183] [4] = 1'b0;
  assign \A[12][183] [3] = 1'b0;
  assign \A[12][183] [2] = 1'b0;
  assign \A[12][183] [1] = 1'b0;
  assign \A[12][183] [0] = 1'b0;
  assign \A[12][184] [4] = 1'b0;
  assign \A[12][184] [3] = 1'b0;
  assign \A[12][184] [2] = 1'b0;
  assign \A[12][184] [1] = 1'b0;
  assign \A[12][184] [0] = 1'b0;
  assign \A[12][185] [4] = 1'b0;
  assign \A[12][185] [3] = 1'b0;
  assign \A[12][185] [2] = 1'b0;
  assign \A[12][185] [0] = 1'b0;
  assign \A[12][186] [4] = 1'b0;
  assign \A[12][186] [3] = 1'b0;
  assign \A[12][186] [2] = 1'b0;
  assign \A[12][186] [1] = 1'b0;
  assign \A[12][186] [0] = 1'b0;
  assign \A[12][187] [0] = 1'b0;
  assign \A[12][188] [4] = 1'b0;
  assign \A[12][188] [3] = 1'b0;
  assign \A[12][188] [2] = 1'b0;
  assign \A[12][188] [0] = 1'b0;
  assign \A[12][190] [1] = 1'b0;
  assign \A[12][192] [4] = 1'b0;
  assign \A[12][192] [3] = 1'b0;
  assign \A[12][192] [2] = 1'b0;
  assign \A[12][192] [0] = 1'b0;
  assign \A[12][193] [4] = 1'b0;
  assign \A[12][193] [3] = 1'b0;
  assign \A[12][193] [2] = 1'b0;
  assign \A[12][193] [1] = 1'b0;
  assign \A[12][193] [0] = 1'b0;
  assign \A[12][194] [4] = 1'b0;
  assign \A[12][194] [3] = 1'b0;
  assign \A[12][194] [2] = 1'b0;
  assign \A[12][194] [1] = 1'b0;
  assign \A[12][195] [4] = 1'b0;
  assign \A[12][195] [3] = 1'b0;
  assign \A[12][195] [2] = 1'b0;
  assign \A[12][195] [1] = 1'b0;
  assign \A[12][196] [1] = 1'b0;
  assign \A[12][197] [4] = 1'b0;
  assign \A[12][197] [3] = 1'b0;
  assign \A[12][197] [2] = 1'b0;
  assign \A[12][197] [1] = 1'b0;
  assign \A[12][197] [0] = 1'b0;
  assign \A[12][198] [4] = 1'b0;
  assign \A[12][198] [3] = 1'b0;
  assign \A[12][198] [2] = 1'b0;
  assign \A[12][198] [0] = 1'b0;
  assign \A[12][200] [4] = 1'b0;
  assign \A[12][200] [3] = 1'b0;
  assign \A[12][200] [2] = 1'b0;
  assign \A[12][200] [1] = 1'b0;
  assign \A[12][201] [4] = 1'b0;
  assign \A[12][201] [3] = 1'b0;
  assign \A[12][201] [2] = 1'b0;
  assign \A[12][201] [1] = 1'b0;
  assign \A[12][201] [0] = 1'b0;
  assign \A[12][202] [4] = 1'b0;
  assign \A[12][202] [3] = 1'b0;
  assign \A[12][202] [2] = 1'b0;
  assign \A[12][202] [1] = 1'b0;
  assign \A[12][204] [4] = 1'b0;
  assign \A[12][204] [3] = 1'b0;
  assign \A[12][204] [2] = 1'b0;
  assign \A[12][204] [1] = 1'b0;
  assign \A[12][204] [0] = 1'b0;
  assign \A[12][205] [0] = 1'b0;
  assign \A[12][207] [4] = 1'b0;
  assign \A[12][207] [3] = 1'b0;
  assign \A[12][207] [2] = 1'b0;
  assign \A[12][208] [4] = 1'b0;
  assign \A[12][208] [3] = 1'b0;
  assign \A[12][208] [2] = 1'b0;
  assign \A[12][208] [1] = 1'b0;
  assign \A[12][208] [0] = 1'b0;
  assign \A[12][209] [4] = 1'b0;
  assign \A[12][209] [3] = 1'b0;
  assign \A[12][209] [2] = 1'b0;
  assign \A[12][209] [1] = 1'b0;
  assign \A[12][209] [0] = 1'b0;
  assign \A[12][210] [1] = 1'b0;
  assign \A[12][211] [4] = 1'b0;
  assign \A[12][211] [3] = 1'b0;
  assign \A[12][211] [2] = 1'b0;
  assign \A[12][211] [1] = 1'b0;
  assign \A[12][211] [0] = 1'b0;
  assign \A[12][212] [4] = 1'b0;
  assign \A[12][212] [3] = 1'b0;
  assign \A[12][212] [2] = 1'b0;
  assign \A[12][212] [1] = 1'b0;
  assign \A[12][212] [0] = 1'b0;
  assign \A[12][213] [0] = 1'b0;
  assign \A[12][214] [4] = 1'b0;
  assign \A[12][214] [3] = 1'b0;
  assign \A[12][214] [2] = 1'b0;
  assign \A[12][214] [1] = 1'b0;
  assign \A[12][216] [4] = 1'b0;
  assign \A[12][216] [3] = 1'b0;
  assign \A[12][216] [2] = 1'b0;
  assign \A[12][216] [1] = 1'b0;
  assign \A[12][216] [0] = 1'b0;
  assign \A[12][217] [4] = 1'b0;
  assign \A[12][217] [3] = 1'b0;
  assign \A[12][217] [2] = 1'b0;
  assign \A[12][217] [1] = 1'b0;
  assign \A[12][218] [0] = 1'b0;
  assign \A[12][220] [4] = 1'b0;
  assign \A[12][220] [3] = 1'b0;
  assign \A[12][220] [2] = 1'b0;
  assign \A[12][220] [0] = 1'b0;
  assign \A[12][221] [4] = 1'b0;
  assign \A[12][221] [3] = 1'b0;
  assign \A[12][221] [2] = 1'b0;
  assign \A[12][222] [4] = 1'b0;
  assign \A[12][222] [3] = 1'b0;
  assign \A[12][222] [2] = 1'b0;
  assign \A[12][222] [1] = 1'b0;
  assign \A[12][222] [0] = 1'b0;
  assign \A[12][224] [4] = 1'b0;
  assign \A[12][224] [3] = 1'b0;
  assign \A[12][224] [2] = 1'b0;
  assign \A[12][224] [1] = 1'b0;
  assign \A[12][227] [4] = 1'b0;
  assign \A[12][227] [3] = 1'b0;
  assign \A[12][227] [2] = 1'b0;
  assign \A[12][227] [1] = 1'b0;
  assign \A[12][228] [4] = 1'b0;
  assign \A[12][228] [3] = 1'b0;
  assign \A[12][228] [2] = 1'b0;
  assign \A[12][228] [1] = 1'b0;
  assign \A[12][228] [0] = 1'b0;
  assign \A[12][230] [4] = 1'b0;
  assign \A[12][230] [3] = 1'b0;
  assign \A[12][230] [2] = 1'b0;
  assign \A[12][230] [1] = 1'b0;
  assign \A[12][230] [0] = 1'b0;
  assign \A[12][232] [1] = 1'b0;
  assign \A[12][233] [4] = 1'b0;
  assign \A[12][233] [3] = 1'b0;
  assign \A[12][233] [2] = 1'b0;
  assign \A[12][233] [1] = 1'b0;
  assign \A[12][234] [0] = 1'b0;
  assign \A[12][235] [4] = 1'b0;
  assign \A[12][235] [3] = 1'b0;
  assign \A[12][235] [2] = 1'b0;
  assign \A[12][235] [1] = 1'b0;
  assign \A[12][237] [0] = 1'b0;
  assign \A[12][238] [4] = 1'b0;
  assign \A[12][238] [3] = 1'b0;
  assign \A[12][238] [2] = 1'b0;
  assign \A[12][238] [1] = 1'b0;
  assign \A[12][238] [0] = 1'b0;
  assign \A[12][239] [0] = 1'b0;
  assign \A[12][241] [4] = 1'b0;
  assign \A[12][241] [3] = 1'b0;
  assign \A[12][241] [2] = 1'b0;
  assign \A[12][241] [1] = 1'b0;
  assign \A[12][241] [0] = 1'b0;
  assign \A[12][242] [4] = 1'b0;
  assign \A[12][242] [3] = 1'b0;
  assign \A[12][242] [2] = 1'b0;
  assign \A[12][242] [0] = 1'b0;
  assign \A[12][243] [4] = 1'b0;
  assign \A[12][243] [3] = 1'b0;
  assign \A[12][243] [2] = 1'b0;
  assign \A[12][243] [1] = 1'b0;
  assign \A[12][244] [4] = 1'b0;
  assign \A[12][244] [3] = 1'b0;
  assign \A[12][244] [2] = 1'b0;
  assign \A[12][244] [1] = 1'b0;
  assign \A[12][245] [4] = 1'b0;
  assign \A[12][245] [3] = 1'b0;
  assign \A[12][245] [2] = 1'b0;
  assign \A[12][245] [1] = 1'b0;
  assign \A[12][245] [0] = 1'b0;
  assign \A[12][246] [4] = 1'b0;
  assign \A[12][246] [3] = 1'b0;
  assign \A[12][246] [2] = 1'b0;
  assign \A[12][246] [1] = 1'b0;
  assign \A[12][246] [0] = 1'b0;
  assign \A[12][247] [4] = 1'b0;
  assign \A[12][247] [3] = 1'b0;
  assign \A[12][247] [2] = 1'b0;
  assign \A[12][247] [1] = 1'b0;
  assign \A[12][247] [0] = 1'b0;
  assign \A[12][248] [4] = 1'b0;
  assign \A[12][248] [3] = 1'b0;
  assign \A[12][248] [2] = 1'b0;
  assign \A[12][248] [1] = 1'b0;
  assign \A[12][248] [0] = 1'b0;
  assign \A[12][249] [0] = 1'b0;
  assign \A[12][250] [4] = 1'b0;
  assign \A[12][250] [3] = 1'b0;
  assign \A[12][250] [2] = 1'b0;
  assign \A[12][250] [0] = 1'b0;
  assign \A[12][251] [4] = 1'b0;
  assign \A[12][251] [3] = 1'b0;
  assign \A[12][251] [1] = 1'b0;
  assign \A[12][251] [0] = 1'b0;
  assign \A[12][253] [0] = 1'b0;
  assign \A[12][254] [4] = 1'b0;
  assign \A[12][254] [3] = 1'b0;
  assign \A[12][254] [2] = 1'b0;
  assign \A[12][254] [1] = 1'b0;
  assign \A[12][254] [0] = 1'b0;
  assign \A[12][255] [4] = 1'b0;
  assign \A[12][255] [3] = 1'b0;
  assign \A[12][255] [2] = 1'b0;
  assign \A[12][255] [1] = 1'b0;
  assign \A[12][255] [0] = 1'b0;
  assign \A[13][0] [4] = 1'b0;
  assign \A[13][0] [3] = 1'b0;
  assign \A[13][0] [2] = 1'b0;
  assign \A[13][0] [1] = 1'b0;
  assign \A[13][0] [0] = 1'b0;
  assign \A[13][3] [4] = 1'b0;
  assign \A[13][3] [3] = 1'b0;
  assign \A[13][3] [2] = 1'b0;
  assign \A[13][3] [1] = 1'b0;
  assign \A[13][4] [4] = 1'b0;
  assign \A[13][4] [3] = 1'b0;
  assign \A[13][4] [1] = 1'b0;
  assign \A[13][4] [0] = 1'b0;
  assign \A[13][5] [0] = 1'b0;
  assign \A[13][6] [4] = 1'b0;
  assign \A[13][6] [3] = 1'b0;
  assign \A[13][6] [2] = 1'b0;
  assign \A[13][6] [1] = 1'b0;
  assign \A[13][8] [4] = 1'b0;
  assign \A[13][8] [3] = 1'b0;
  assign \A[13][8] [2] = 1'b0;
  assign \A[13][8] [1] = 1'b0;
  assign \A[13][9] [4] = 1'b0;
  assign \A[13][9] [3] = 1'b0;
  assign \A[13][9] [2] = 1'b0;
  assign \A[13][9] [1] = 1'b0;
  assign \A[13][10] [4] = 1'b0;
  assign \A[13][10] [3] = 1'b0;
  assign \A[13][10] [2] = 1'b0;
  assign \A[13][10] [1] = 1'b0;
  assign \A[13][10] [0] = 1'b0;
  assign \A[13][12] [4] = 1'b0;
  assign \A[13][12] [3] = 1'b0;
  assign \A[13][12] [2] = 1'b0;
  assign \A[13][12] [1] = 1'b0;
  assign \A[13][14] [4] = 1'b0;
  assign \A[13][14] [3] = 1'b0;
  assign \A[13][14] [2] = 1'b0;
  assign \A[13][14] [1] = 1'b0;
  assign \A[13][15] [4] = 1'b0;
  assign \A[13][15] [3] = 1'b0;
  assign \A[13][15] [2] = 1'b0;
  assign \A[13][15] [1] = 1'b0;
  assign \A[13][16] [0] = 1'b0;
  assign \A[13][17] [0] = 1'b0;
  assign \A[13][18] [4] = 1'b0;
  assign \A[13][18] [3] = 1'b0;
  assign \A[13][18] [2] = 1'b0;
  assign \A[13][18] [1] = 1'b0;
  assign \A[13][18] [0] = 1'b0;
  assign \A[13][20] [0] = 1'b0;
  assign \A[13][21] [4] = 1'b0;
  assign \A[13][21] [3] = 1'b0;
  assign \A[13][21] [2] = 1'b0;
  assign \A[13][21] [1] = 1'b0;
  assign \A[13][22] [4] = 1'b0;
  assign \A[13][22] [3] = 1'b0;
  assign \A[13][22] [2] = 1'b0;
  assign \A[13][22] [1] = 1'b0;
  assign \A[13][23] [4] = 1'b0;
  assign \A[13][23] [3] = 1'b0;
  assign \A[13][23] [2] = 1'b0;
  assign \A[13][23] [1] = 1'b0;
  assign \A[13][23] [0] = 1'b0;
  assign \A[13][24] [4] = 1'b0;
  assign \A[13][24] [3] = 1'b0;
  assign \A[13][24] [2] = 1'b0;
  assign \A[13][24] [1] = 1'b0;
  assign \A[13][24] [0] = 1'b0;
  assign \A[13][25] [4] = 1'b0;
  assign \A[13][25] [3] = 1'b0;
  assign \A[13][25] [2] = 1'b0;
  assign \A[13][25] [1] = 1'b0;
  assign \A[13][25] [0] = 1'b0;
  assign \A[13][26] [0] = 1'b0;
  assign \A[13][28] [4] = 1'b0;
  assign \A[13][28] [3] = 1'b0;
  assign \A[13][28] [2] = 1'b0;
  assign \A[13][28] [0] = 1'b0;
  assign \A[13][29] [4] = 1'b0;
  assign \A[13][29] [3] = 1'b0;
  assign \A[13][29] [2] = 1'b0;
  assign \A[13][29] [1] = 1'b0;
  assign \A[13][29] [0] = 1'b0;
  assign \A[13][30] [4] = 1'b0;
  assign \A[13][30] [3] = 1'b0;
  assign \A[13][30] [2] = 1'b0;
  assign \A[13][30] [1] = 1'b0;
  assign \A[13][31] [4] = 1'b0;
  assign \A[13][31] [3] = 1'b0;
  assign \A[13][31] [2] = 1'b0;
  assign \A[13][31] [1] = 1'b0;
  assign \A[13][32] [4] = 1'b0;
  assign \A[13][32] [3] = 1'b0;
  assign \A[13][32] [2] = 1'b0;
  assign \A[13][33] [4] = 1'b0;
  assign \A[13][33] [3] = 1'b0;
  assign \A[13][33] [2] = 1'b0;
  assign \A[13][33] [1] = 1'b0;
  assign \A[13][34] [4] = 1'b0;
  assign \A[13][34] [3] = 1'b0;
  assign \A[13][34] [2] = 1'b0;
  assign \A[13][34] [1] = 1'b0;
  assign \A[13][34] [0] = 1'b0;
  assign \A[13][35] [4] = 1'b0;
  assign \A[13][35] [3] = 1'b0;
  assign \A[13][35] [2] = 1'b0;
  assign \A[13][35] [1] = 1'b0;
  assign \A[13][35] [0] = 1'b0;
  assign \A[13][36] [1] = 1'b0;
  assign \A[13][36] [0] = 1'b0;
  assign \A[13][38] [4] = 1'b0;
  assign \A[13][38] [3] = 1'b0;
  assign \A[13][38] [2] = 1'b0;
  assign \A[13][38] [1] = 1'b0;
  assign \A[13][38] [0] = 1'b0;
  assign \A[13][39] [4] = 1'b0;
  assign \A[13][39] [3] = 1'b0;
  assign \A[13][39] [2] = 1'b0;
  assign \A[13][39] [1] = 1'b0;
  assign \A[13][39] [0] = 1'b0;
  assign \A[13][40] [4] = 1'b0;
  assign \A[13][40] [3] = 1'b0;
  assign \A[13][40] [2] = 1'b0;
  assign \A[13][40] [1] = 1'b0;
  assign \A[13][40] [0] = 1'b0;
  assign \A[13][41] [4] = 1'b0;
  assign \A[13][41] [3] = 1'b0;
  assign \A[13][41] [2] = 1'b0;
  assign \A[13][41] [1] = 1'b0;
  assign \A[13][42] [4] = 1'b0;
  assign \A[13][42] [3] = 1'b0;
  assign \A[13][42] [2] = 1'b0;
  assign \A[13][42] [1] = 1'b0;
  assign \A[13][43] [4] = 1'b0;
  assign \A[13][43] [3] = 1'b0;
  assign \A[13][43] [2] = 1'b0;
  assign \A[13][43] [1] = 1'b0;
  assign \A[13][44] [4] = 1'b0;
  assign \A[13][44] [3] = 1'b0;
  assign \A[13][44] [2] = 1'b0;
  assign \A[13][44] [1] = 1'b0;
  assign \A[13][45] [4] = 1'b0;
  assign \A[13][45] [3] = 1'b0;
  assign \A[13][45] [2] = 1'b0;
  assign \A[13][45] [1] = 1'b0;
  assign \A[13][45] [0] = 1'b0;
  assign \A[13][47] [4] = 1'b0;
  assign \A[13][47] [3] = 1'b0;
  assign \A[13][47] [2] = 1'b0;
  assign \A[13][47] [1] = 1'b0;
  assign \A[13][47] [0] = 1'b0;
  assign \A[13][48] [4] = 1'b0;
  assign \A[13][48] [3] = 1'b0;
  assign \A[13][48] [2] = 1'b0;
  assign \A[13][48] [0] = 1'b0;
  assign \A[13][49] [4] = 1'b0;
  assign \A[13][49] [3] = 1'b0;
  assign \A[13][49] [2] = 1'b0;
  assign \A[13][49] [1] = 1'b0;
  assign \A[13][49] [0] = 1'b0;
  assign \A[13][50] [4] = 1'b0;
  assign \A[13][50] [3] = 1'b0;
  assign \A[13][50] [2] = 1'b0;
  assign \A[13][50] [1] = 1'b0;
  assign \A[13][51] [4] = 1'b0;
  assign \A[13][51] [3] = 1'b0;
  assign \A[13][51] [2] = 1'b0;
  assign \A[13][52] [4] = 1'b0;
  assign \A[13][52] [3] = 1'b0;
  assign \A[13][52] [2] = 1'b0;
  assign \A[13][52] [0] = 1'b0;
  assign \A[13][53] [4] = 1'b0;
  assign \A[13][53] [3] = 1'b0;
  assign \A[13][53] [2] = 1'b0;
  assign \A[13][53] [1] = 1'b0;
  assign \A[13][53] [0] = 1'b0;
  assign \A[13][54] [0] = 1'b0;
  assign \A[13][55] [4] = 1'b0;
  assign \A[13][55] [3] = 1'b0;
  assign \A[13][55] [2] = 1'b0;
  assign \A[13][55] [1] = 1'b0;
  assign \A[13][55] [0] = 1'b0;
  assign \A[13][58] [4] = 1'b0;
  assign \A[13][58] [3] = 1'b0;
  assign \A[13][58] [2] = 1'b0;
  assign \A[13][58] [1] = 1'b0;
  assign \A[13][58] [0] = 1'b0;
  assign \A[13][59] [0] = 1'b0;
  assign \A[13][60] [1] = 1'b0;
  assign \A[13][61] [4] = 1'b0;
  assign \A[13][61] [3] = 1'b0;
  assign \A[13][61] [2] = 1'b0;
  assign \A[13][61] [1] = 1'b0;
  assign \A[13][62] [4] = 1'b0;
  assign \A[13][62] [3] = 1'b0;
  assign \A[13][62] [2] = 1'b0;
  assign \A[13][62] [1] = 1'b0;
  assign \A[13][63] [4] = 1'b0;
  assign \A[13][63] [3] = 1'b0;
  assign \A[13][63] [2] = 1'b0;
  assign \A[13][64] [4] = 1'b0;
  assign \A[13][64] [3] = 1'b0;
  assign \A[13][64] [2] = 1'b0;
  assign \A[13][64] [1] = 1'b0;
  assign \A[13][65] [4] = 1'b0;
  assign \A[13][65] [3] = 1'b0;
  assign \A[13][65] [2] = 1'b0;
  assign \A[13][65] [1] = 1'b0;
  assign \A[13][66] [4] = 1'b0;
  assign \A[13][66] [3] = 1'b0;
  assign \A[13][66] [2] = 1'b0;
  assign \A[13][66] [1] = 1'b0;
  assign \A[13][66] [0] = 1'b0;
  assign \A[13][67] [0] = 1'b0;
  assign \A[13][68] [4] = 1'b0;
  assign \A[13][68] [3] = 1'b0;
  assign \A[13][68] [2] = 1'b0;
  assign \A[13][68] [1] = 1'b0;
  assign \A[13][69] [4] = 1'b0;
  assign \A[13][69] [3] = 1'b0;
  assign \A[13][69] [2] = 1'b0;
  assign \A[13][69] [1] = 1'b0;
  assign \A[13][70] [1] = 1'b0;
  assign \A[13][71] [4] = 1'b0;
  assign \A[13][71] [3] = 1'b0;
  assign \A[13][71] [2] = 1'b0;
  assign \A[13][71] [1] = 1'b0;
  assign \A[13][71] [0] = 1'b0;
  assign \A[13][72] [4] = 1'b0;
  assign \A[13][72] [3] = 1'b0;
  assign \A[13][72] [2] = 1'b0;
  assign \A[13][74] [4] = 1'b0;
  assign \A[13][74] [3] = 1'b0;
  assign \A[13][74] [2] = 1'b0;
  assign \A[13][74] [1] = 1'b0;
  assign \A[13][74] [0] = 1'b0;
  assign \A[13][75] [4] = 1'b0;
  assign \A[13][75] [3] = 1'b0;
  assign \A[13][75] [2] = 1'b0;
  assign \A[13][75] [1] = 1'b0;
  assign \A[13][76] [4] = 1'b0;
  assign \A[13][76] [3] = 1'b0;
  assign \A[13][76] [2] = 1'b0;
  assign \A[13][76] [1] = 1'b0;
  assign \A[13][76] [0] = 1'b0;
  assign \A[13][77] [4] = 1'b0;
  assign \A[13][77] [3] = 1'b0;
  assign \A[13][77] [2] = 1'b0;
  assign \A[13][77] [1] = 1'b0;
  assign \A[13][78] [4] = 1'b0;
  assign \A[13][78] [3] = 1'b0;
  assign \A[13][78] [2] = 1'b0;
  assign \A[13][78] [1] = 1'b0;
  assign \A[13][78] [0] = 1'b0;
  assign \A[13][79] [0] = 1'b0;
  assign \A[13][80] [4] = 1'b0;
  assign \A[13][80] [3] = 1'b0;
  assign \A[13][80] [2] = 1'b0;
  assign \A[13][80] [1] = 1'b0;
  assign \A[13][80] [0] = 1'b0;
  assign \A[13][82] [4] = 1'b0;
  assign \A[13][82] [3] = 1'b0;
  assign \A[13][82] [2] = 1'b0;
  assign \A[13][83] [4] = 1'b0;
  assign \A[13][83] [3] = 1'b0;
  assign \A[13][83] [2] = 1'b0;
  assign \A[13][83] [1] = 1'b0;
  assign \A[13][84] [0] = 1'b0;
  assign \A[13][85] [0] = 1'b0;
  assign \A[13][86] [4] = 1'b0;
  assign \A[13][86] [3] = 1'b0;
  assign \A[13][86] [2] = 1'b0;
  assign \A[13][86] [1] = 1'b0;
  assign \A[13][86] [0] = 1'b0;
  assign \A[13][87] [0] = 1'b0;
  assign \A[13][88] [4] = 1'b0;
  assign \A[13][88] [3] = 1'b0;
  assign \A[13][88] [2] = 1'b0;
  assign \A[13][88] [1] = 1'b0;
  assign \A[13][89] [4] = 1'b0;
  assign \A[13][89] [3] = 1'b0;
  assign \A[13][89] [2] = 1'b0;
  assign \A[13][89] [1] = 1'b0;
  assign \A[13][90] [0] = 1'b0;
  assign \A[13][92] [4] = 1'b0;
  assign \A[13][92] [3] = 1'b0;
  assign \A[13][92] [2] = 1'b0;
  assign \A[13][92] [0] = 1'b0;
  assign \A[13][93] [4] = 1'b0;
  assign \A[13][93] [3] = 1'b0;
  assign \A[13][93] [2] = 1'b0;
  assign \A[13][93] [0] = 1'b0;
  assign \A[13][94] [4] = 1'b0;
  assign \A[13][94] [3] = 1'b0;
  assign \A[13][94] [2] = 1'b0;
  assign \A[13][94] [1] = 1'b0;
  assign \A[13][95] [4] = 1'b0;
  assign \A[13][95] [3] = 1'b0;
  assign \A[13][95] [2] = 1'b0;
  assign \A[13][95] [1] = 1'b0;
  assign \A[13][96] [4] = 1'b0;
  assign \A[13][96] [3] = 1'b0;
  assign \A[13][96] [2] = 1'b0;
  assign \A[13][96] [1] = 1'b0;
  assign \A[13][96] [0] = 1'b0;
  assign \A[13][97] [1] = 1'b0;
  assign \A[13][98] [4] = 1'b0;
  assign \A[13][98] [3] = 1'b0;
  assign \A[13][98] [2] = 1'b0;
  assign \A[13][98] [1] = 1'b0;
  assign \A[13][99] [4] = 1'b0;
  assign \A[13][99] [3] = 1'b0;
  assign \A[13][99] [2] = 1'b0;
  assign \A[13][99] [0] = 1'b0;
  assign \A[13][100] [4] = 1'b0;
  assign \A[13][100] [3] = 1'b0;
  assign \A[13][100] [2] = 1'b0;
  assign \A[13][100] [1] = 1'b0;
  assign \A[13][100] [0] = 1'b0;
  assign \A[13][101] [4] = 1'b0;
  assign \A[13][101] [3] = 1'b0;
  assign \A[13][101] [2] = 1'b0;
  assign \A[13][101] [1] = 1'b0;
  assign \A[13][102] [4] = 1'b0;
  assign \A[13][102] [3] = 1'b0;
  assign \A[13][102] [2] = 1'b0;
  assign \A[13][102] [1] = 1'b0;
  assign \A[13][103] [0] = 1'b0;
  assign \A[13][105] [4] = 1'b0;
  assign \A[13][105] [3] = 1'b0;
  assign \A[13][105] [2] = 1'b0;
  assign \A[13][105] [1] = 1'b0;
  assign \A[13][105] [0] = 1'b0;
  assign \A[13][107] [4] = 1'b0;
  assign \A[13][107] [3] = 1'b0;
  assign \A[13][107] [2] = 1'b0;
  assign \A[13][107] [1] = 1'b0;
  assign \A[13][108] [4] = 1'b0;
  assign \A[13][108] [3] = 1'b0;
  assign \A[13][108] [2] = 1'b0;
  assign \A[13][108] [1] = 1'b0;
  assign \A[13][110] [4] = 1'b0;
  assign \A[13][110] [3] = 1'b0;
  assign \A[13][110] [2] = 1'b0;
  assign \A[13][110] [1] = 1'b0;
  assign \A[13][110] [0] = 1'b0;
  assign \A[13][111] [4] = 1'b0;
  assign \A[13][111] [3] = 1'b0;
  assign \A[13][111] [2] = 1'b0;
  assign \A[13][111] [1] = 1'b0;
  assign \A[13][111] [0] = 1'b0;
  assign \A[13][112] [4] = 1'b0;
  assign \A[13][112] [3] = 1'b0;
  assign \A[13][112] [2] = 1'b0;
  assign \A[13][112] [1] = 1'b0;
  assign \A[13][115] [4] = 1'b0;
  assign \A[13][115] [3] = 1'b0;
  assign \A[13][115] [2] = 1'b0;
  assign \A[13][115] [1] = 1'b0;
  assign \A[13][115] [0] = 1'b0;
  assign \A[13][116] [4] = 1'b0;
  assign \A[13][116] [3] = 1'b0;
  assign \A[13][116] [2] = 1'b0;
  assign \A[13][116] [1] = 1'b0;
  assign \A[13][116] [0] = 1'b0;
  assign \A[13][119] [4] = 1'b0;
  assign \A[13][119] [3] = 1'b0;
  assign \A[13][119] [2] = 1'b0;
  assign \A[13][119] [1] = 1'b0;
  assign \A[13][121] [4] = 1'b0;
  assign \A[13][121] [3] = 1'b0;
  assign \A[13][121] [2] = 1'b0;
  assign \A[13][121] [1] = 1'b0;
  assign \A[13][122] [4] = 1'b0;
  assign \A[13][122] [3] = 1'b0;
  assign \A[13][122] [2] = 1'b0;
  assign \A[13][122] [1] = 1'b0;
  assign \A[13][122] [0] = 1'b0;
  assign \A[13][123] [4] = 1'b0;
  assign \A[13][123] [3] = 1'b0;
  assign \A[13][123] [2] = 1'b0;
  assign \A[13][123] [1] = 1'b0;
  assign \A[13][124] [4] = 1'b0;
  assign \A[13][124] [3] = 1'b0;
  assign \A[13][124] [2] = 1'b0;
  assign \A[13][124] [1] = 1'b0;
  assign \A[13][124] [0] = 1'b0;
  assign \A[13][125] [4] = 1'b0;
  assign \A[13][125] [3] = 1'b0;
  assign \A[13][125] [2] = 1'b0;
  assign \A[13][125] [1] = 1'b0;
  assign \A[13][127] [4] = 1'b0;
  assign \A[13][127] [3] = 1'b0;
  assign \A[13][127] [2] = 1'b0;
  assign \A[13][127] [1] = 1'b0;
  assign \A[13][128] [4] = 1'b0;
  assign \A[13][128] [3] = 1'b0;
  assign \A[13][128] [2] = 1'b0;
  assign \A[13][128] [0] = 1'b0;
  assign \A[13][129] [4] = 1'b0;
  assign \A[13][129] [3] = 1'b0;
  assign \A[13][129] [2] = 1'b0;
  assign \A[13][129] [1] = 1'b0;
  assign \A[13][129] [0] = 1'b0;
  assign \A[13][130] [0] = 1'b0;
  assign \A[13][131] [4] = 1'b0;
  assign \A[13][131] [3] = 1'b0;
  assign \A[13][131] [2] = 1'b0;
  assign \A[13][131] [0] = 1'b0;
  assign \A[13][132] [4] = 1'b0;
  assign \A[13][132] [3] = 1'b0;
  assign \A[13][132] [2] = 1'b0;
  assign \A[13][132] [1] = 1'b0;
  assign \A[13][132] [0] = 1'b0;
  assign \A[13][133] [4] = 1'b0;
  assign \A[13][133] [3] = 1'b0;
  assign \A[13][133] [2] = 1'b0;
  assign \A[13][133] [1] = 1'b0;
  assign \A[13][134] [0] = 1'b0;
  assign \A[13][136] [4] = 1'b0;
  assign \A[13][136] [3] = 1'b0;
  assign \A[13][136] [2] = 1'b0;
  assign \A[13][136] [1] = 1'b0;
  assign \A[13][136] [0] = 1'b0;
  assign \A[13][138] [4] = 1'b0;
  assign \A[13][138] [3] = 1'b0;
  assign \A[13][138] [2] = 1'b0;
  assign \A[13][138] [1] = 1'b0;
  assign \A[13][138] [0] = 1'b0;
  assign \A[13][139] [0] = 1'b0;
  assign \A[13][141] [0] = 1'b0;
  assign \A[13][142] [4] = 1'b0;
  assign \A[13][142] [3] = 1'b0;
  assign \A[13][142] [2] = 1'b0;
  assign \A[13][142] [1] = 1'b0;
  assign \A[13][142] [0] = 1'b0;
  assign \A[13][143] [2] = 1'b0;
  assign \A[13][144] [4] = 1'b0;
  assign \A[13][144] [3] = 1'b0;
  assign \A[13][144] [2] = 1'b0;
  assign \A[13][144] [1] = 1'b0;
  assign \A[13][145] [4] = 1'b0;
  assign \A[13][145] [3] = 1'b0;
  assign \A[13][145] [2] = 1'b0;
  assign \A[13][145] [1] = 1'b0;
  assign \A[13][145] [0] = 1'b0;
  assign \A[13][147] [4] = 1'b0;
  assign \A[13][147] [3] = 1'b0;
  assign \A[13][147] [2] = 1'b0;
  assign \A[13][147] [1] = 1'b0;
  assign \A[13][147] [0] = 1'b0;
  assign \A[13][148] [0] = 1'b0;
  assign \A[13][149] [4] = 1'b0;
  assign \A[13][149] [3] = 1'b0;
  assign \A[13][149] [2] = 1'b0;
  assign \A[13][149] [1] = 1'b0;
  assign \A[13][149] [0] = 1'b0;
  assign \A[13][150] [4] = 1'b0;
  assign \A[13][150] [3] = 1'b0;
  assign \A[13][150] [2] = 1'b0;
  assign \A[13][150] [0] = 1'b0;
  assign \A[13][151] [4] = 1'b0;
  assign \A[13][151] [3] = 1'b0;
  assign \A[13][151] [2] = 1'b0;
  assign \A[13][151] [1] = 1'b0;
  assign \A[13][151] [0] = 1'b0;
  assign \A[13][152] [4] = 1'b0;
  assign \A[13][152] [3] = 1'b0;
  assign \A[13][152] [2] = 1'b0;
  assign \A[13][152] [0] = 1'b0;
  assign \A[13][153] [4] = 1'b0;
  assign \A[13][153] [3] = 1'b0;
  assign \A[13][153] [2] = 1'b0;
  assign \A[13][153] [0] = 1'b0;
  assign \A[13][154] [4] = 1'b0;
  assign \A[13][154] [3] = 1'b0;
  assign \A[13][154] [2] = 1'b0;
  assign \A[13][154] [1] = 1'b0;
  assign \A[13][154] [0] = 1'b0;
  assign \A[13][155] [4] = 1'b0;
  assign \A[13][155] [3] = 1'b0;
  assign \A[13][155] [2] = 1'b0;
  assign \A[13][155] [1] = 1'b0;
  assign \A[13][155] [0] = 1'b0;
  assign \A[13][156] [4] = 1'b0;
  assign \A[13][156] [3] = 1'b0;
  assign \A[13][156] [2] = 1'b0;
  assign \A[13][156] [1] = 1'b0;
  assign \A[13][157] [4] = 1'b0;
  assign \A[13][157] [3] = 1'b0;
  assign \A[13][157] [2] = 1'b0;
  assign \A[13][157] [0] = 1'b0;
  assign \A[13][158] [4] = 1'b0;
  assign \A[13][158] [3] = 1'b0;
  assign \A[13][158] [2] = 1'b0;
  assign \A[13][158] [1] = 1'b0;
  assign \A[13][159] [0] = 1'b0;
  assign \A[13][160] [4] = 1'b0;
  assign \A[13][160] [3] = 1'b0;
  assign \A[13][160] [2] = 1'b0;
  assign \A[13][160] [1] = 1'b0;
  assign \A[13][161] [4] = 1'b0;
  assign \A[13][161] [3] = 1'b0;
  assign \A[13][161] [2] = 1'b0;
  assign \A[13][161] [0] = 1'b0;
  assign \A[13][163] [4] = 1'b0;
  assign \A[13][163] [3] = 1'b0;
  assign \A[13][163] [2] = 1'b0;
  assign \A[13][163] [1] = 1'b0;
  assign \A[13][163] [0] = 1'b0;
  assign \A[13][164] [4] = 1'b0;
  assign \A[13][164] [3] = 1'b0;
  assign \A[13][164] [2] = 1'b0;
  assign \A[13][164] [1] = 1'b0;
  assign \A[13][164] [0] = 1'b0;
  assign \A[13][165] [4] = 1'b0;
  assign \A[13][165] [3] = 1'b0;
  assign \A[13][165] [2] = 1'b0;
  assign \A[13][165] [1] = 1'b0;
  assign \A[13][167] [4] = 1'b0;
  assign \A[13][167] [3] = 1'b0;
  assign \A[13][167] [2] = 1'b0;
  assign \A[13][170] [4] = 1'b0;
  assign \A[13][170] [3] = 1'b0;
  assign \A[13][170] [2] = 1'b0;
  assign \A[13][170] [1] = 1'b0;
  assign \A[13][170] [0] = 1'b0;
  assign \A[13][172] [0] = 1'b0;
  assign \A[13][173] [4] = 1'b0;
  assign \A[13][173] [3] = 1'b0;
  assign \A[13][173] [2] = 1'b0;
  assign \A[13][173] [1] = 1'b0;
  assign \A[13][175] [4] = 1'b0;
  assign \A[13][175] [3] = 1'b0;
  assign \A[13][175] [2] = 1'b0;
  assign \A[13][175] [0] = 1'b0;
  assign \A[13][176] [4] = 1'b0;
  assign \A[13][176] [3] = 1'b0;
  assign \A[13][176] [2] = 1'b0;
  assign \A[13][176] [0] = 1'b0;
  assign \A[13][177] [4] = 1'b0;
  assign \A[13][177] [3] = 1'b0;
  assign \A[13][177] [2] = 1'b0;
  assign \A[13][177] [1] = 1'b0;
  assign \A[13][177] [0] = 1'b0;
  assign \A[13][178] [4] = 1'b0;
  assign \A[13][178] [3] = 1'b0;
  assign \A[13][178] [2] = 1'b0;
  assign \A[13][178] [1] = 1'b0;
  assign \A[13][178] [0] = 1'b0;
  assign \A[13][179] [4] = 1'b0;
  assign \A[13][179] [3] = 1'b0;
  assign \A[13][179] [2] = 1'b0;
  assign \A[13][179] [1] = 1'b0;
  assign \A[13][180] [4] = 1'b0;
  assign \A[13][180] [3] = 1'b0;
  assign \A[13][180] [2] = 1'b0;
  assign \A[13][180] [1] = 1'b0;
  assign \A[13][181] [4] = 1'b0;
  assign \A[13][181] [3] = 1'b0;
  assign \A[13][181] [2] = 1'b0;
  assign \A[13][181] [0] = 1'b0;
  assign \A[13][182] [4] = 1'b0;
  assign \A[13][182] [3] = 1'b0;
  assign \A[13][182] [2] = 1'b0;
  assign \A[13][182] [1] = 1'b0;
  assign \A[13][183] [4] = 1'b0;
  assign \A[13][183] [3] = 1'b0;
  assign \A[13][183] [2] = 1'b0;
  assign \A[13][183] [1] = 1'b0;
  assign \A[13][183] [0] = 1'b0;
  assign \A[13][184] [4] = 1'b0;
  assign \A[13][184] [3] = 1'b0;
  assign \A[13][184] [2] = 1'b0;
  assign \A[13][184] [0] = 1'b0;
  assign \A[13][185] [4] = 1'b0;
  assign \A[13][185] [3] = 1'b0;
  assign \A[13][185] [2] = 1'b0;
  assign \A[13][185] [1] = 1'b0;
  assign \A[13][185] [0] = 1'b0;
  assign \A[13][187] [0] = 1'b0;
  assign \A[13][188] [4] = 1'b0;
  assign \A[13][188] [3] = 1'b0;
  assign \A[13][188] [2] = 1'b0;
  assign \A[13][188] [1] = 1'b0;
  assign \A[13][188] [0] = 1'b0;
  assign \A[13][190] [4] = 1'b0;
  assign \A[13][190] [3] = 1'b0;
  assign \A[13][190] [2] = 1'b0;
  assign \A[13][190] [1] = 1'b0;
  assign \A[13][190] [0] = 1'b0;
  assign \A[13][191] [4] = 1'b0;
  assign \A[13][191] [3] = 1'b0;
  assign \A[13][191] [2] = 1'b0;
  assign \A[13][191] [0] = 1'b0;
  assign \A[13][192] [4] = 1'b0;
  assign \A[13][192] [3] = 1'b0;
  assign \A[13][192] [2] = 1'b0;
  assign \A[13][193] [0] = 1'b0;
  assign \A[13][194] [4] = 1'b0;
  assign \A[13][194] [3] = 1'b0;
  assign \A[13][194] [2] = 1'b0;
  assign \A[13][194] [1] = 1'b0;
  assign \A[13][195] [4] = 1'b0;
  assign \A[13][195] [3] = 1'b0;
  assign \A[13][195] [2] = 1'b0;
  assign \A[13][195] [0] = 1'b0;
  assign \A[13][196] [4] = 1'b0;
  assign \A[13][196] [3] = 1'b0;
  assign \A[13][196] [2] = 1'b0;
  assign \A[13][196] [1] = 1'b0;
  assign \A[13][196] [0] = 1'b0;
  assign \A[13][197] [4] = 1'b0;
  assign \A[13][197] [3] = 1'b0;
  assign \A[13][197] [2] = 1'b0;
  assign \A[13][197] [1] = 1'b0;
  assign \A[13][197] [0] = 1'b0;
  assign \A[13][198] [4] = 1'b0;
  assign \A[13][198] [3] = 1'b0;
  assign \A[13][198] [2] = 1'b0;
  assign \A[13][198] [1] = 1'b0;
  assign \A[13][199] [4] = 1'b0;
  assign \A[13][199] [3] = 1'b0;
  assign \A[13][199] [2] = 1'b0;
  assign \A[13][199] [1] = 1'b0;
  assign \A[13][200] [4] = 1'b0;
  assign \A[13][200] [3] = 1'b0;
  assign \A[13][200] [2] = 1'b0;
  assign \A[13][200] [1] = 1'b0;
  assign \A[13][200] [0] = 1'b0;
  assign \A[13][201] [4] = 1'b0;
  assign \A[13][201] [3] = 1'b0;
  assign \A[13][201] [2] = 1'b0;
  assign \A[13][201] [1] = 1'b0;
  assign \A[13][202] [4] = 1'b0;
  assign \A[13][202] [3] = 1'b0;
  assign \A[13][202] [2] = 1'b0;
  assign \A[13][202] [1] = 1'b0;
  assign \A[13][204] [4] = 1'b0;
  assign \A[13][204] [3] = 1'b0;
  assign \A[13][204] [2] = 1'b0;
  assign \A[13][204] [1] = 1'b0;
  assign \A[13][205] [4] = 1'b0;
  assign \A[13][205] [3] = 1'b0;
  assign \A[13][205] [2] = 1'b0;
  assign \A[13][206] [4] = 1'b0;
  assign \A[13][206] [3] = 1'b0;
  assign \A[13][206] [2] = 1'b0;
  assign \A[13][206] [1] = 1'b0;
  assign \A[13][206] [0] = 1'b0;
  assign \A[13][208] [4] = 1'b0;
  assign \A[13][208] [3] = 1'b0;
  assign \A[13][208] [2] = 1'b0;
  assign \A[13][208] [0] = 1'b0;
  assign \A[13][209] [4] = 1'b0;
  assign \A[13][209] [3] = 1'b0;
  assign \A[13][209] [2] = 1'b0;
  assign \A[13][209] [1] = 1'b0;
  assign \A[13][209] [0] = 1'b0;
  assign \A[13][210] [4] = 1'b0;
  assign \A[13][210] [3] = 1'b0;
  assign \A[13][210] [2] = 1'b0;
  assign \A[13][210] [0] = 1'b0;
  assign \A[13][212] [4] = 1'b0;
  assign \A[13][212] [3] = 1'b0;
  assign \A[13][212] [2] = 1'b0;
  assign \A[13][212] [1] = 1'b0;
  assign \A[13][212] [0] = 1'b0;
  assign \A[13][213] [4] = 1'b0;
  assign \A[13][213] [3] = 1'b0;
  assign \A[13][213] [2] = 1'b0;
  assign \A[13][213] [0] = 1'b0;
  assign \A[13][214] [4] = 1'b0;
  assign \A[13][214] [3] = 1'b0;
  assign \A[13][214] [2] = 1'b0;
  assign \A[13][214] [1] = 1'b0;
  assign \A[13][214] [0] = 1'b0;
  assign \A[13][217] [4] = 1'b0;
  assign \A[13][217] [3] = 1'b0;
  assign \A[13][217] [2] = 1'b0;
  assign \A[13][218] [4] = 1'b0;
  assign \A[13][218] [3] = 1'b0;
  assign \A[13][218] [2] = 1'b0;
  assign \A[13][218] [1] = 1'b0;
  assign \A[13][218] [0] = 1'b0;
  assign \A[13][219] [4] = 1'b0;
  assign \A[13][219] [3] = 1'b0;
  assign \A[13][219] [2] = 1'b0;
  assign \A[13][219] [1] = 1'b0;
  assign \A[13][219] [0] = 1'b0;
  assign \A[13][220] [4] = 1'b0;
  assign \A[13][220] [3] = 1'b0;
  assign \A[13][220] [2] = 1'b0;
  assign \A[13][221] [4] = 1'b0;
  assign \A[13][221] [3] = 1'b0;
  assign \A[13][221] [2] = 1'b0;
  assign \A[13][221] [1] = 1'b0;
  assign \A[13][221] [0] = 1'b0;
  assign \A[13][224] [4] = 1'b0;
  assign \A[13][224] [3] = 1'b0;
  assign \A[13][224] [2] = 1'b0;
  assign \A[13][224] [0] = 1'b0;
  assign \A[13][226] [0] = 1'b0;
  assign \A[13][227] [4] = 1'b0;
  assign \A[13][227] [3] = 1'b0;
  assign \A[13][227] [2] = 1'b0;
  assign \A[13][227] [1] = 1'b0;
  assign \A[13][227] [0] = 1'b0;
  assign \A[13][229] [4] = 1'b0;
  assign \A[13][229] [3] = 1'b0;
  assign \A[13][229] [2] = 1'b0;
  assign \A[13][229] [0] = 1'b0;
  assign \A[13][230] [4] = 1'b0;
  assign \A[13][230] [3] = 1'b0;
  assign \A[13][230] [2] = 1'b0;
  assign \A[13][230] [0] = 1'b0;
  assign \A[13][231] [4] = 1'b0;
  assign \A[13][231] [3] = 1'b0;
  assign \A[13][231] [2] = 1'b0;
  assign \A[13][232] [4] = 1'b0;
  assign \A[13][232] [3] = 1'b0;
  assign \A[13][232] [2] = 1'b0;
  assign \A[13][232] [1] = 1'b0;
  assign \A[13][232] [0] = 1'b0;
  assign \A[13][233] [4] = 1'b0;
  assign \A[13][233] [3] = 1'b0;
  assign \A[13][233] [2] = 1'b0;
  assign \A[13][234] [4] = 1'b0;
  assign \A[13][234] [3] = 1'b0;
  assign \A[13][234] [2] = 1'b0;
  assign \A[13][234] [1] = 1'b0;
  assign \A[13][234] [0] = 1'b0;
  assign \A[13][235] [4] = 1'b0;
  assign \A[13][235] [3] = 1'b0;
  assign \A[13][235] [2] = 1'b0;
  assign \A[13][235] [1] = 1'b0;
  assign \A[13][238] [4] = 1'b0;
  assign \A[13][238] [3] = 1'b0;
  assign \A[13][238] [2] = 1'b0;
  assign \A[13][238] [1] = 1'b0;
  assign \A[13][238] [0] = 1'b0;
  assign \A[13][239] [0] = 1'b0;
  assign \A[13][240] [4] = 1'b0;
  assign \A[13][240] [3] = 1'b0;
  assign \A[13][240] [2] = 1'b0;
  assign \A[13][240] [1] = 1'b0;
  assign \A[13][240] [0] = 1'b0;
  assign \A[13][242] [0] = 1'b0;
  assign \A[13][243] [4] = 1'b0;
  assign \A[13][243] [3] = 1'b0;
  assign \A[13][243] [2] = 1'b0;
  assign \A[13][243] [1] = 1'b0;
  assign \A[13][243] [0] = 1'b0;
  assign \A[13][244] [4] = 1'b0;
  assign \A[13][244] [3] = 1'b0;
  assign \A[13][244] [2] = 1'b0;
  assign \A[13][244] [0] = 1'b0;
  assign \A[13][245] [4] = 1'b0;
  assign \A[13][245] [3] = 1'b0;
  assign \A[13][245] [2] = 1'b0;
  assign \A[13][245] [1] = 1'b0;
  assign \A[13][246] [4] = 1'b0;
  assign \A[13][246] [3] = 1'b0;
  assign \A[13][246] [2] = 1'b0;
  assign \A[13][246] [0] = 1'b0;
  assign \A[13][247] [0] = 1'b0;
  assign \A[13][248] [4] = 1'b0;
  assign \A[13][248] [3] = 1'b0;
  assign \A[13][248] [2] = 1'b0;
  assign \A[13][248] [1] = 1'b0;
  assign \A[13][250] [4] = 1'b0;
  assign \A[13][250] [3] = 1'b0;
  assign \A[13][250] [2] = 1'b0;
  assign \A[13][250] [1] = 1'b0;
  assign \A[13][251] [4] = 1'b0;
  assign \A[13][251] [3] = 1'b0;
  assign \A[13][251] [2] = 1'b0;
  assign \A[13][251] [1] = 1'b0;
  assign \A[13][252] [0] = 1'b0;
  assign \A[13][254] [4] = 1'b0;
  assign \A[13][254] [3] = 1'b0;
  assign \A[13][254] [2] = 1'b0;
  assign \A[13][254] [1] = 1'b0;
  assign \A[13][255] [4] = 1'b0;
  assign \A[13][255] [3] = 1'b0;
  assign \A[13][255] [2] = 1'b0;
  assign \A[13][255] [1] = 1'b0;
  assign \A[13][255] [0] = 1'b0;
  assign \A[14][0] [4] = 1'b0;
  assign \A[14][0] [3] = 1'b0;
  assign \A[14][0] [2] = 1'b0;
  assign \A[14][0] [1] = 1'b0;
  assign \A[14][1] [1] = 1'b0;
  assign \A[14][1] [0] = 1'b0;
  assign \A[14][2] [4] = 1'b0;
  assign \A[14][2] [3] = 1'b0;
  assign \A[14][2] [2] = 1'b0;
  assign \A[14][2] [1] = 1'b0;
  assign \A[14][2] [0] = 1'b0;
  assign \A[14][5] [4] = 1'b0;
  assign \A[14][5] [3] = 1'b0;
  assign \A[14][5] [2] = 1'b0;
  assign \A[14][5] [0] = 1'b0;
  assign \A[14][6] [4] = 1'b0;
  assign \A[14][6] [3] = 1'b0;
  assign \A[14][6] [2] = 1'b0;
  assign \A[14][6] [1] = 1'b0;
  assign \A[14][7] [4] = 1'b0;
  assign \A[14][7] [3] = 1'b0;
  assign \A[14][7] [2] = 1'b0;
  assign \A[14][7] [0] = 1'b0;
  assign \A[14][8] [4] = 1'b0;
  assign \A[14][8] [3] = 1'b0;
  assign \A[14][8] [2] = 1'b0;
  assign \A[14][8] [1] = 1'b0;
  assign \A[14][9] [4] = 1'b0;
  assign \A[14][9] [3] = 1'b0;
  assign \A[14][9] [2] = 1'b0;
  assign \A[14][9] [1] = 1'b0;
  assign \A[14][9] [0] = 1'b0;
  assign \A[14][13] [4] = 1'b0;
  assign \A[14][13] [3] = 1'b0;
  assign \A[14][13] [2] = 1'b0;
  assign \A[14][13] [1] = 1'b0;
  assign \A[14][13] [0] = 1'b0;
  assign \A[14][14] [4] = 1'b0;
  assign \A[14][14] [3] = 1'b0;
  assign \A[14][14] [2] = 1'b0;
  assign \A[14][14] [1] = 1'b0;
  assign \A[14][14] [0] = 1'b0;
  assign \A[14][15] [1] = 1'b0;
  assign \A[14][16] [4] = 1'b0;
  assign \A[14][16] [3] = 1'b0;
  assign \A[14][16] [2] = 1'b0;
  assign \A[14][16] [1] = 1'b0;
  assign \A[14][16] [0] = 1'b0;
  assign \A[14][17] [4] = 1'b0;
  assign \A[14][17] [3] = 1'b0;
  assign \A[14][17] [2] = 1'b0;
  assign \A[14][18] [4] = 1'b0;
  assign \A[14][18] [3] = 1'b0;
  assign \A[14][18] [2] = 1'b0;
  assign \A[14][18] [1] = 1'b0;
  assign \A[14][20] [4] = 1'b0;
  assign \A[14][20] [3] = 1'b0;
  assign \A[14][20] [2] = 1'b0;
  assign \A[14][20] [1] = 1'b0;
  assign \A[14][20] [0] = 1'b0;
  assign \A[14][21] [1] = 1'b0;
  assign \A[14][22] [4] = 1'b0;
  assign \A[14][22] [3] = 1'b0;
  assign \A[14][22] [2] = 1'b0;
  assign \A[14][22] [1] = 1'b0;
  assign \A[14][22] [0] = 1'b0;
  assign \A[14][23] [4] = 1'b0;
  assign \A[14][23] [3] = 1'b0;
  assign \A[14][23] [2] = 1'b0;
  assign \A[14][23] [1] = 1'b0;
  assign \A[14][24] [4] = 1'b0;
  assign \A[14][24] [3] = 1'b0;
  assign \A[14][24] [2] = 1'b0;
  assign \A[14][25] [4] = 1'b0;
  assign \A[14][25] [3] = 1'b0;
  assign \A[14][25] [2] = 1'b0;
  assign \A[14][25] [1] = 1'b0;
  assign \A[14][25] [0] = 1'b0;
  assign \A[14][26] [4] = 1'b0;
  assign \A[14][26] [3] = 1'b0;
  assign \A[14][26] [2] = 1'b0;
  assign \A[14][26] [1] = 1'b0;
  assign \A[14][26] [0] = 1'b0;
  assign \A[14][27] [4] = 1'b0;
  assign \A[14][27] [3] = 1'b0;
  assign \A[14][27] [2] = 1'b0;
  assign \A[14][27] [0] = 1'b0;
  assign \A[14][28] [4] = 1'b0;
  assign \A[14][28] [3] = 1'b0;
  assign \A[14][28] [2] = 1'b0;
  assign \A[14][28] [1] = 1'b0;
  assign \A[14][28] [0] = 1'b0;
  assign \A[14][29] [4] = 1'b0;
  assign \A[14][29] [3] = 1'b0;
  assign \A[14][29] [2] = 1'b0;
  assign \A[14][29] [1] = 1'b0;
  assign \A[14][29] [0] = 1'b0;
  assign \A[14][30] [0] = 1'b0;
  assign \A[14][31] [4] = 1'b0;
  assign \A[14][31] [3] = 1'b0;
  assign \A[14][31] [2] = 1'b0;
  assign \A[14][31] [1] = 1'b0;
  assign \A[14][31] [0] = 1'b0;
  assign \A[14][33] [4] = 1'b0;
  assign \A[14][33] [3] = 1'b0;
  assign \A[14][33] [1] = 1'b0;
  assign \A[14][33] [0] = 1'b0;
  assign \A[14][35] [0] = 1'b0;
  assign \A[14][37] [4] = 1'b0;
  assign \A[14][37] [3] = 1'b0;
  assign \A[14][37] [2] = 1'b0;
  assign \A[14][37] [0] = 1'b0;
  assign \A[14][39] [4] = 1'b0;
  assign \A[14][39] [3] = 1'b0;
  assign \A[14][39] [2] = 1'b0;
  assign \A[14][39] [0] = 1'b0;
  assign \A[14][41] [4] = 1'b0;
  assign \A[14][41] [3] = 1'b0;
  assign \A[14][41] [2] = 1'b0;
  assign \A[14][41] [1] = 1'b0;
  assign \A[14][41] [0] = 1'b0;
  assign \A[14][42] [0] = 1'b0;
  assign \A[14][43] [4] = 1'b0;
  assign \A[14][43] [3] = 1'b0;
  assign \A[14][43] [2] = 1'b0;
  assign \A[14][43] [1] = 1'b0;
  assign \A[14][43] [0] = 1'b0;
  assign \A[14][44] [0] = 1'b0;
  assign \A[14][45] [1] = 1'b0;
  assign \A[14][46] [0] = 1'b0;
  assign \A[14][47] [4] = 1'b0;
  assign \A[14][47] [3] = 1'b0;
  assign \A[14][47] [2] = 1'b0;
  assign \A[14][47] [1] = 1'b0;
  assign \A[14][48] [4] = 1'b0;
  assign \A[14][48] [3] = 1'b0;
  assign \A[14][48] [2] = 1'b0;
  assign \A[14][48] [1] = 1'b0;
  assign \A[14][49] [4] = 1'b0;
  assign \A[14][49] [3] = 1'b0;
  assign \A[14][49] [2] = 1'b0;
  assign \A[14][50] [4] = 1'b0;
  assign \A[14][50] [3] = 1'b0;
  assign \A[14][50] [2] = 1'b0;
  assign \A[14][51] [0] = 1'b0;
  assign \A[14][52] [4] = 1'b0;
  assign \A[14][52] [3] = 1'b0;
  assign \A[14][52] [2] = 1'b0;
  assign \A[14][52] [1] = 1'b0;
  assign \A[14][53] [4] = 1'b0;
  assign \A[14][53] [3] = 1'b0;
  assign \A[14][53] [2] = 1'b0;
  assign \A[14][53] [1] = 1'b0;
  assign \A[14][53] [0] = 1'b0;
  assign \A[14][54] [4] = 1'b0;
  assign \A[14][54] [3] = 1'b0;
  assign \A[14][54] [2] = 1'b0;
  assign \A[14][54] [1] = 1'b0;
  assign \A[14][55] [1] = 1'b0;
  assign \A[14][56] [4] = 1'b0;
  assign \A[14][56] [3] = 1'b0;
  assign \A[14][56] [2] = 1'b0;
  assign \A[14][56] [1] = 1'b0;
  assign \A[14][57] [0] = 1'b0;
  assign \A[14][58] [4] = 1'b0;
  assign \A[14][58] [3] = 1'b0;
  assign \A[14][58] [2] = 1'b0;
  assign \A[14][58] [1] = 1'b0;
  assign \A[14][58] [0] = 1'b0;
  assign \A[14][62] [4] = 1'b0;
  assign \A[14][62] [3] = 1'b0;
  assign \A[14][62] [2] = 1'b0;
  assign \A[14][62] [1] = 1'b0;
  assign \A[14][63] [4] = 1'b0;
  assign \A[14][63] [3] = 1'b0;
  assign \A[14][63] [2] = 1'b0;
  assign \A[14][63] [0] = 1'b0;
  assign \A[14][64] [4] = 1'b0;
  assign \A[14][64] [3] = 1'b0;
  assign \A[14][64] [2] = 1'b0;
  assign \A[14][64] [1] = 1'b0;
  assign \A[14][65] [4] = 1'b0;
  assign \A[14][65] [3] = 1'b0;
  assign \A[14][65] [2] = 1'b0;
  assign \A[14][65] [0] = 1'b0;
  assign \A[14][66] [4] = 1'b0;
  assign \A[14][66] [3] = 1'b0;
  assign \A[14][66] [2] = 1'b0;
  assign \A[14][66] [1] = 1'b0;
  assign \A[14][67] [4] = 1'b0;
  assign \A[14][67] [3] = 1'b0;
  assign \A[14][67] [2] = 1'b0;
  assign \A[14][67] [1] = 1'b0;
  assign \A[14][67] [0] = 1'b0;
  assign \A[14][68] [4] = 1'b0;
  assign \A[14][68] [3] = 1'b0;
  assign \A[14][68] [2] = 1'b0;
  assign \A[14][68] [1] = 1'b0;
  assign \A[14][69] [4] = 1'b0;
  assign \A[14][69] [3] = 1'b0;
  assign \A[14][69] [2] = 1'b0;
  assign \A[14][69] [1] = 1'b0;
  assign \A[14][70] [4] = 1'b0;
  assign \A[14][70] [3] = 1'b0;
  assign \A[14][70] [2] = 1'b0;
  assign \A[14][70] [1] = 1'b0;
  assign \A[14][70] [0] = 1'b0;
  assign \A[14][71] [4] = 1'b0;
  assign \A[14][71] [3] = 1'b0;
  assign \A[14][71] [2] = 1'b0;
  assign \A[14][71] [1] = 1'b0;
  assign \A[14][71] [0] = 1'b0;
  assign \A[14][73] [4] = 1'b0;
  assign \A[14][73] [3] = 1'b0;
  assign \A[14][73] [2] = 1'b0;
  assign \A[14][73] [1] = 1'b0;
  assign \A[14][74] [0] = 1'b0;
  assign \A[14][75] [4] = 1'b0;
  assign \A[14][75] [3] = 1'b0;
  assign \A[14][75] [2] = 1'b0;
  assign \A[14][75] [0] = 1'b0;
  assign \A[14][77] [0] = 1'b0;
  assign \A[14][78] [4] = 1'b0;
  assign \A[14][78] [3] = 1'b0;
  assign \A[14][78] [2] = 1'b0;
  assign \A[14][78] [1] = 1'b0;
  assign \A[14][78] [0] = 1'b0;
  assign \A[14][80] [0] = 1'b0;
  assign \A[14][81] [4] = 1'b0;
  assign \A[14][81] [3] = 1'b0;
  assign \A[14][81] [2] = 1'b0;
  assign \A[14][81] [1] = 1'b0;
  assign \A[14][81] [0] = 1'b0;
  assign \A[14][82] [4] = 1'b0;
  assign \A[14][82] [3] = 1'b0;
  assign \A[14][82] [1] = 1'b0;
  assign \A[14][82] [0] = 1'b0;
  assign \A[14][83] [4] = 1'b0;
  assign \A[14][83] [3] = 1'b0;
  assign \A[14][83] [2] = 1'b0;
  assign \A[14][83] [1] = 1'b0;
  assign \A[14][83] [0] = 1'b0;
  assign \A[14][84] [4] = 1'b0;
  assign \A[14][84] [3] = 1'b0;
  assign \A[14][84] [2] = 1'b0;
  assign \A[14][84] [1] = 1'b0;
  assign \A[14][84] [0] = 1'b0;
  assign \A[14][85] [4] = 1'b0;
  assign \A[14][85] [3] = 1'b0;
  assign \A[14][85] [2] = 1'b0;
  assign \A[14][85] [1] = 1'b0;
  assign \A[14][85] [0] = 1'b0;
  assign \A[14][86] [4] = 1'b0;
  assign \A[14][86] [3] = 1'b0;
  assign \A[14][86] [1] = 1'b0;
  assign \A[14][86] [0] = 1'b0;
  assign \A[14][87] [1] = 1'b0;
  assign \A[14][88] [4] = 1'b0;
  assign \A[14][88] [3] = 1'b0;
  assign \A[14][88] [2] = 1'b0;
  assign \A[14][88] [1] = 1'b0;
  assign \A[14][89] [4] = 1'b0;
  assign \A[14][89] [3] = 1'b0;
  assign \A[14][89] [2] = 1'b0;
  assign \A[14][89] [1] = 1'b0;
  assign \A[14][89] [0] = 1'b0;
  assign \A[14][90] [4] = 1'b0;
  assign \A[14][90] [3] = 1'b0;
  assign \A[14][90] [2] = 1'b0;
  assign \A[14][90] [1] = 1'b0;
  assign \A[14][90] [0] = 1'b0;
  assign \A[14][91] [4] = 1'b0;
  assign \A[14][91] [3] = 1'b0;
  assign \A[14][91] [2] = 1'b0;
  assign \A[14][91] [1] = 1'b0;
  assign \A[14][91] [0] = 1'b0;
  assign \A[14][92] [4] = 1'b0;
  assign \A[14][92] [3] = 1'b0;
  assign \A[14][92] [2] = 1'b0;
  assign \A[14][92] [1] = 1'b0;
  assign \A[14][92] [0] = 1'b0;
  assign \A[14][93] [4] = 1'b0;
  assign \A[14][93] [3] = 1'b0;
  assign \A[14][93] [2] = 1'b0;
  assign \A[14][93] [1] = 1'b0;
  assign \A[14][93] [0] = 1'b0;
  assign \A[14][94] [4] = 1'b0;
  assign \A[14][94] [3] = 1'b0;
  assign \A[14][94] [2] = 1'b0;
  assign \A[14][94] [1] = 1'b0;
  assign \A[14][97] [4] = 1'b0;
  assign \A[14][97] [3] = 1'b0;
  assign \A[14][97] [2] = 1'b0;
  assign \A[14][97] [1] = 1'b0;
  assign \A[14][97] [0] = 1'b0;
  assign \A[14][98] [4] = 1'b0;
  assign \A[14][98] [3] = 1'b0;
  assign \A[14][98] [2] = 1'b0;
  assign \A[14][98] [1] = 1'b0;
  assign \A[14][99] [1] = 1'b0;
  assign \A[14][100] [4] = 1'b0;
  assign \A[14][100] [3] = 1'b0;
  assign \A[14][100] [2] = 1'b0;
  assign \A[14][100] [1] = 1'b0;
  assign \A[14][100] [0] = 1'b0;
  assign \A[14][102] [4] = 1'b0;
  assign \A[14][102] [3] = 1'b0;
  assign \A[14][102] [2] = 1'b0;
  assign \A[14][102] [0] = 1'b0;
  assign \A[14][103] [1] = 1'b0;
  assign \A[14][104] [4] = 1'b0;
  assign \A[14][104] [3] = 1'b0;
  assign \A[14][104] [2] = 1'b0;
  assign \A[14][104] [1] = 1'b0;
  assign \A[14][104] [0] = 1'b0;
  assign \A[14][107] [4] = 1'b0;
  assign \A[14][107] [3] = 1'b0;
  assign \A[14][107] [2] = 1'b0;
  assign \A[14][107] [1] = 1'b0;
  assign \A[14][108] [4] = 1'b0;
  assign \A[14][108] [3] = 1'b0;
  assign \A[14][108] [2] = 1'b0;
  assign \A[14][108] [1] = 1'b0;
  assign \A[14][108] [0] = 1'b0;
  assign \A[14][109] [4] = 1'b0;
  assign \A[14][109] [3] = 1'b0;
  assign \A[14][109] [2] = 1'b0;
  assign \A[14][109] [1] = 1'b0;
  assign \A[14][110] [4] = 1'b0;
  assign \A[14][110] [3] = 1'b0;
  assign \A[14][110] [2] = 1'b0;
  assign \A[14][110] [1] = 1'b0;
  assign \A[14][111] [0] = 1'b0;
  assign \A[14][112] [0] = 1'b0;
  assign \A[14][113] [4] = 1'b0;
  assign \A[14][113] [3] = 1'b0;
  assign \A[14][113] [2] = 1'b0;
  assign \A[14][113] [1] = 1'b0;
  assign \A[14][114] [1] = 1'b0;
  assign \A[14][115] [4] = 1'b0;
  assign \A[14][115] [3] = 1'b0;
  assign \A[14][115] [2] = 1'b0;
  assign \A[14][115] [1] = 1'b0;
  assign \A[14][117] [4] = 1'b0;
  assign \A[14][117] [3] = 1'b0;
  assign \A[14][117] [2] = 1'b0;
  assign \A[14][117] [1] = 1'b0;
  assign \A[14][119] [4] = 1'b0;
  assign \A[14][119] [3] = 1'b0;
  assign \A[14][119] [2] = 1'b0;
  assign \A[14][119] [1] = 1'b0;
  assign \A[14][119] [0] = 1'b0;
  assign \A[14][120] [4] = 1'b0;
  assign \A[14][120] [3] = 1'b0;
  assign \A[14][120] [2] = 1'b0;
  assign \A[14][120] [1] = 1'b0;
  assign \A[14][120] [0] = 1'b0;
  assign \A[14][121] [4] = 1'b0;
  assign \A[14][121] [3] = 1'b0;
  assign \A[14][121] [2] = 1'b0;
  assign \A[14][121] [1] = 1'b0;
  assign \A[14][121] [0] = 1'b0;
  assign \A[14][122] [4] = 1'b0;
  assign \A[14][122] [3] = 1'b0;
  assign \A[14][122] [2] = 1'b0;
  assign \A[14][122] [1] = 1'b0;
  assign \A[14][122] [0] = 1'b0;
  assign \A[14][123] [4] = 1'b0;
  assign \A[14][123] [3] = 1'b0;
  assign \A[14][123] [2] = 1'b0;
  assign \A[14][123] [1] = 1'b0;
  assign \A[14][124] [4] = 1'b0;
  assign \A[14][124] [3] = 1'b0;
  assign \A[14][124] [2] = 1'b0;
  assign \A[14][124] [1] = 1'b0;
  assign \A[14][125] [0] = 1'b0;
  assign \A[14][126] [4] = 1'b0;
  assign \A[14][126] [3] = 1'b0;
  assign \A[14][126] [2] = 1'b0;
  assign \A[14][126] [0] = 1'b0;
  assign \A[14][127] [4] = 1'b0;
  assign \A[14][127] [3] = 1'b0;
  assign \A[14][127] [2] = 1'b0;
  assign \A[14][127] [1] = 1'b0;
  assign \A[14][127] [0] = 1'b0;
  assign \A[14][128] [4] = 1'b0;
  assign \A[14][128] [3] = 1'b0;
  assign \A[14][128] [2] = 1'b0;
  assign \A[14][128] [1] = 1'b0;
  assign \A[14][130] [4] = 1'b0;
  assign \A[14][130] [3] = 1'b0;
  assign \A[14][130] [2] = 1'b0;
  assign \A[14][130] [1] = 1'b0;
  assign \A[14][130] [0] = 1'b0;
  assign \A[14][131] [1] = 1'b0;
  assign \A[14][132] [4] = 1'b0;
  assign \A[14][132] [3] = 1'b0;
  assign \A[14][132] [2] = 1'b0;
  assign \A[14][132] [1] = 1'b0;
  assign \A[14][136] [4] = 1'b0;
  assign \A[14][136] [3] = 1'b0;
  assign \A[14][136] [2] = 1'b0;
  assign \A[14][136] [1] = 1'b0;
  assign \A[14][136] [0] = 1'b0;
  assign \A[14][137] [0] = 1'b0;
  assign \A[14][138] [4] = 1'b0;
  assign \A[14][138] [3] = 1'b0;
  assign \A[14][138] [1] = 1'b0;
  assign \A[14][138] [0] = 1'b0;
  assign \A[14][139] [4] = 1'b0;
  assign \A[14][139] [3] = 1'b0;
  assign \A[14][139] [2] = 1'b0;
  assign \A[14][139] [1] = 1'b0;
  assign \A[14][140] [4] = 1'b0;
  assign \A[14][140] [3] = 1'b0;
  assign \A[14][140] [2] = 1'b0;
  assign \A[14][140] [1] = 1'b0;
  assign \A[14][140] [0] = 1'b0;
  assign \A[14][143] [4] = 1'b0;
  assign \A[14][143] [3] = 1'b0;
  assign \A[14][143] [2] = 1'b0;
  assign \A[14][143] [1] = 1'b0;
  assign \A[14][143] [0] = 1'b0;
  assign \A[14][144] [4] = 1'b0;
  assign \A[14][144] [3] = 1'b0;
  assign \A[14][144] [2] = 1'b0;
  assign \A[14][144] [1] = 1'b0;
  assign \A[14][144] [0] = 1'b0;
  assign \A[14][148] [4] = 1'b0;
  assign \A[14][148] [3] = 1'b0;
  assign \A[14][148] [2] = 1'b0;
  assign \A[14][148] [1] = 1'b0;
  assign \A[14][148] [0] = 1'b0;
  assign \A[14][152] [4] = 1'b0;
  assign \A[14][152] [3] = 1'b0;
  assign \A[14][152] [2] = 1'b0;
  assign \A[14][152] [1] = 1'b0;
  assign \A[14][152] [0] = 1'b0;
  assign \A[14][153] [4] = 1'b0;
  assign \A[14][153] [3] = 1'b0;
  assign \A[14][153] [2] = 1'b0;
  assign \A[14][153] [1] = 1'b0;
  assign \A[14][155] [4] = 1'b0;
  assign \A[14][155] [3] = 1'b0;
  assign \A[14][155] [2] = 1'b0;
  assign \A[14][155] [0] = 1'b0;
  assign \A[14][156] [4] = 1'b0;
  assign \A[14][156] [3] = 1'b0;
  assign \A[14][156] [2] = 1'b0;
  assign \A[14][156] [1] = 1'b0;
  assign \A[14][157] [0] = 1'b0;
  assign \A[14][158] [4] = 1'b0;
  assign \A[14][158] [3] = 1'b0;
  assign \A[14][158] [2] = 1'b0;
  assign \A[14][158] [1] = 1'b0;
  assign \A[14][158] [0] = 1'b0;
  assign \A[14][160] [4] = 1'b0;
  assign \A[14][160] [3] = 1'b0;
  assign \A[14][160] [2] = 1'b0;
  assign \A[14][160] [1] = 1'b0;
  assign \A[14][161] [4] = 1'b0;
  assign \A[14][161] [3] = 1'b0;
  assign \A[14][161] [2] = 1'b0;
  assign \A[14][161] [0] = 1'b0;
  assign \A[14][162] [4] = 1'b0;
  assign \A[14][162] [3] = 1'b0;
  assign \A[14][162] [2] = 1'b0;
  assign \A[14][162] [1] = 1'b0;
  assign \A[14][162] [0] = 1'b0;
  assign \A[14][163] [4] = 1'b0;
  assign \A[14][163] [3] = 1'b0;
  assign \A[14][163] [2] = 1'b0;
  assign \A[14][163] [1] = 1'b0;
  assign \A[14][163] [0] = 1'b0;
  assign \A[14][164] [0] = 1'b0;
  assign \A[14][165] [4] = 1'b0;
  assign \A[14][165] [3] = 1'b0;
  assign \A[14][165] [2] = 1'b0;
  assign \A[14][165] [1] = 1'b0;
  assign \A[14][166] [4] = 1'b0;
  assign \A[14][166] [3] = 1'b0;
  assign \A[14][166] [2] = 1'b0;
  assign \A[14][166] [1] = 1'b0;
  assign \A[14][166] [0] = 1'b0;
  assign \A[14][167] [4] = 1'b0;
  assign \A[14][167] [3] = 1'b0;
  assign \A[14][167] [2] = 1'b0;
  assign \A[14][167] [1] = 1'b0;
  assign \A[14][167] [0] = 1'b0;
  assign \A[14][168] [4] = 1'b0;
  assign \A[14][168] [3] = 1'b0;
  assign \A[14][168] [2] = 1'b0;
  assign \A[14][168] [1] = 1'b0;
  assign \A[14][168] [0] = 1'b0;
  assign \A[14][169] [4] = 1'b0;
  assign \A[14][169] [3] = 1'b0;
  assign \A[14][169] [2] = 1'b0;
  assign \A[14][169] [1] = 1'b0;
  assign \A[14][170] [4] = 1'b0;
  assign \A[14][170] [3] = 1'b0;
  assign \A[14][170] [2] = 1'b0;
  assign \A[14][170] [1] = 1'b0;
  assign \A[14][170] [0] = 1'b0;
  assign \A[14][172] [4] = 1'b0;
  assign \A[14][172] [3] = 1'b0;
  assign \A[14][172] [2] = 1'b0;
  assign \A[14][172] [1] = 1'b0;
  assign \A[14][172] [0] = 1'b0;
  assign \A[14][173] [4] = 1'b0;
  assign \A[14][173] [3] = 1'b0;
  assign \A[14][173] [2] = 1'b0;
  assign \A[14][174] [4] = 1'b0;
  assign \A[14][174] [3] = 1'b0;
  assign \A[14][174] [2] = 1'b0;
  assign \A[14][174] [1] = 1'b0;
  assign \A[14][175] [4] = 1'b0;
  assign \A[14][175] [3] = 1'b0;
  assign \A[14][175] [2] = 1'b0;
  assign \A[14][175] [1] = 1'b0;
  assign \A[14][176] [4] = 1'b0;
  assign \A[14][176] [3] = 1'b0;
  assign \A[14][176] [2] = 1'b0;
  assign \A[14][176] [1] = 1'b0;
  assign \A[14][176] [0] = 1'b0;
  assign \A[14][177] [4] = 1'b0;
  assign \A[14][177] [3] = 1'b0;
  assign \A[14][177] [2] = 1'b0;
  assign \A[14][177] [1] = 1'b0;
  assign \A[14][179] [4] = 1'b0;
  assign \A[14][179] [3] = 1'b0;
  assign \A[14][179] [2] = 1'b0;
  assign \A[14][179] [1] = 1'b0;
  assign \A[14][179] [0] = 1'b0;
  assign \A[14][180] [4] = 1'b0;
  assign \A[14][180] [3] = 1'b0;
  assign \A[14][180] [2] = 1'b0;
  assign \A[14][180] [0] = 1'b0;
  assign \A[14][181] [4] = 1'b0;
  assign \A[14][181] [3] = 1'b0;
  assign \A[14][181] [2] = 1'b0;
  assign \A[14][181] [1] = 1'b0;
  assign \A[14][183] [1] = 1'b0;
  assign \A[14][183] [0] = 1'b0;
  assign \A[14][184] [4] = 1'b0;
  assign \A[14][184] [3] = 1'b0;
  assign \A[14][184] [2] = 1'b0;
  assign \A[14][184] [1] = 1'b0;
  assign \A[14][184] [0] = 1'b0;
  assign \A[14][186] [4] = 1'b0;
  assign \A[14][186] [3] = 1'b0;
  assign \A[14][186] [2] = 1'b0;
  assign \A[14][186] [1] = 1'b0;
  assign \A[14][186] [0] = 1'b0;
  assign \A[14][187] [4] = 1'b0;
  assign \A[14][187] [3] = 1'b0;
  assign \A[14][187] [2] = 1'b0;
  assign \A[14][187] [0] = 1'b0;
  assign \A[14][188] [4] = 1'b0;
  assign \A[14][188] [3] = 1'b0;
  assign \A[14][188] [2] = 1'b0;
  assign \A[14][188] [1] = 1'b0;
  assign \A[14][188] [0] = 1'b0;
  assign \A[14][190] [4] = 1'b0;
  assign \A[14][190] [3] = 1'b0;
  assign \A[14][190] [2] = 1'b0;
  assign \A[14][190] [0] = 1'b0;
  assign \A[14][191] [4] = 1'b0;
  assign \A[14][191] [3] = 1'b0;
  assign \A[14][191] [2] = 1'b0;
  assign \A[14][191] [1] = 1'b0;
  assign \A[14][192] [4] = 1'b0;
  assign \A[14][192] [3] = 1'b0;
  assign \A[14][192] [2] = 1'b0;
  assign \A[14][192] [1] = 1'b0;
  assign \A[14][192] [0] = 1'b0;
  assign \A[14][193] [0] = 1'b0;
  assign \A[14][195] [4] = 1'b0;
  assign \A[14][195] [3] = 1'b0;
  assign \A[14][195] [2] = 1'b0;
  assign \A[14][196] [4] = 1'b0;
  assign \A[14][196] [3] = 1'b0;
  assign \A[14][196] [2] = 1'b0;
  assign \A[14][196] [1] = 1'b0;
  assign \A[14][197] [4] = 1'b0;
  assign \A[14][197] [3] = 1'b0;
  assign \A[14][197] [2] = 1'b0;
  assign \A[14][197] [1] = 1'b0;
  assign \A[14][197] [0] = 1'b0;
  assign \A[14][198] [4] = 1'b0;
  assign \A[14][198] [3] = 1'b0;
  assign \A[14][198] [2] = 1'b0;
  assign \A[14][199] [4] = 1'b0;
  assign \A[14][199] [3] = 1'b0;
  assign \A[14][199] [2] = 1'b0;
  assign \A[14][199] [1] = 1'b0;
  assign \A[14][199] [0] = 1'b0;
  assign \A[14][200] [0] = 1'b0;
  assign \A[14][202] [4] = 1'b0;
  assign \A[14][202] [3] = 1'b0;
  assign \A[14][202] [2] = 1'b0;
  assign \A[14][202] [1] = 1'b0;
  assign \A[14][203] [4] = 1'b0;
  assign \A[14][203] [3] = 1'b0;
  assign \A[14][203] [2] = 1'b0;
  assign \A[14][204] [4] = 1'b0;
  assign \A[14][204] [3] = 1'b0;
  assign \A[14][204] [2] = 1'b0;
  assign \A[14][204] [1] = 1'b0;
  assign \A[14][205] [4] = 1'b0;
  assign \A[14][205] [3] = 1'b0;
  assign \A[14][205] [2] = 1'b0;
  assign \A[14][205] [1] = 1'b0;
  assign \A[14][208] [4] = 1'b0;
  assign \A[14][208] [3] = 1'b0;
  assign \A[14][208] [2] = 1'b0;
  assign \A[14][210] [1] = 1'b0;
  assign \A[14][211] [4] = 1'b0;
  assign \A[14][211] [3] = 1'b0;
  assign \A[14][211] [2] = 1'b0;
  assign \A[14][211] [1] = 1'b0;
  assign \A[14][211] [0] = 1'b0;
  assign \A[14][212] [4] = 1'b0;
  assign \A[14][212] [3] = 1'b0;
  assign \A[14][212] [2] = 1'b0;
  assign \A[14][212] [1] = 1'b0;
  assign \A[14][212] [0] = 1'b0;
  assign \A[14][213] [1] = 1'b0;
  assign \A[14][215] [4] = 1'b0;
  assign \A[14][215] [3] = 1'b0;
  assign \A[14][215] [2] = 1'b0;
  assign \A[14][215] [1] = 1'b0;
  assign \A[14][215] [0] = 1'b0;
  assign \A[14][216] [4] = 1'b0;
  assign \A[14][216] [3] = 1'b0;
  assign \A[14][216] [2] = 1'b0;
  assign \A[14][216] [1] = 1'b0;
  assign \A[14][217] [4] = 1'b0;
  assign \A[14][217] [3] = 1'b0;
  assign \A[14][217] [2] = 1'b0;
  assign \A[14][217] [1] = 1'b0;
  assign \A[14][217] [0] = 1'b0;
  assign \A[14][218] [4] = 1'b0;
  assign \A[14][218] [3] = 1'b0;
  assign \A[14][218] [2] = 1'b0;
  assign \A[14][218] [0] = 1'b0;
  assign \A[14][219] [4] = 1'b0;
  assign \A[14][219] [3] = 1'b0;
  assign \A[14][219] [2] = 1'b0;
  assign \A[14][219] [1] = 1'b0;
  assign \A[14][222] [4] = 1'b0;
  assign \A[14][222] [3] = 1'b0;
  assign \A[14][222] [2] = 1'b0;
  assign \A[14][222] [1] = 1'b0;
  assign \A[14][222] [0] = 1'b0;
  assign \A[14][223] [4] = 1'b0;
  assign \A[14][223] [3] = 1'b0;
  assign \A[14][223] [2] = 1'b0;
  assign \A[14][223] [1] = 1'b0;
  assign \A[14][224] [1] = 1'b0;
  assign \A[14][226] [4] = 1'b0;
  assign \A[14][226] [3] = 1'b0;
  assign \A[14][226] [2] = 1'b0;
  assign \A[14][226] [1] = 1'b0;
  assign \A[14][226] [0] = 1'b0;
  assign \A[14][228] [4] = 1'b0;
  assign \A[14][228] [3] = 1'b0;
  assign \A[14][228] [2] = 1'b0;
  assign \A[14][228] [1] = 1'b0;
  assign \A[14][229] [4] = 1'b0;
  assign \A[14][229] [3] = 1'b0;
  assign \A[14][229] [2] = 1'b0;
  assign \A[14][229] [1] = 1'b0;
  assign \A[14][233] [4] = 1'b0;
  assign \A[14][233] [3] = 1'b0;
  assign \A[14][233] [2] = 1'b0;
  assign \A[14][233] [1] = 1'b0;
  assign \A[14][234] [4] = 1'b0;
  assign \A[14][234] [3] = 1'b0;
  assign \A[14][234] [2] = 1'b0;
  assign \A[14][234] [1] = 1'b0;
  assign \A[14][237] [4] = 1'b0;
  assign \A[14][237] [3] = 1'b0;
  assign \A[14][237] [2] = 1'b0;
  assign \A[14][237] [1] = 1'b0;
  assign \A[14][237] [0] = 1'b0;
  assign \A[14][240] [4] = 1'b0;
  assign \A[14][240] [3] = 1'b0;
  assign \A[14][240] [2] = 1'b0;
  assign \A[14][240] [1] = 1'b0;
  assign \A[14][241] [0] = 1'b0;
  assign \A[14][242] [4] = 1'b0;
  assign \A[14][242] [3] = 1'b0;
  assign \A[14][242] [2] = 1'b0;
  assign \A[14][242] [1] = 1'b0;
  assign \A[14][242] [0] = 1'b0;
  assign \A[14][243] [4] = 1'b0;
  assign \A[14][243] [3] = 1'b0;
  assign \A[14][243] [2] = 1'b0;
  assign \A[14][243] [0] = 1'b0;
  assign \A[14][244] [4] = 1'b0;
  assign \A[14][244] [3] = 1'b0;
  assign \A[14][244] [2] = 1'b0;
  assign \A[14][244] [1] = 1'b0;
  assign \A[14][244] [0] = 1'b0;
  assign \A[14][245] [4] = 1'b0;
  assign \A[14][245] [3] = 1'b0;
  assign \A[14][245] [2] = 1'b0;
  assign \A[14][245] [1] = 1'b0;
  assign \A[14][245] [0] = 1'b0;
  assign \A[14][247] [4] = 1'b0;
  assign \A[14][247] [3] = 1'b0;
  assign \A[14][247] [2] = 1'b0;
  assign \A[14][247] [1] = 1'b0;
  assign \A[14][247] [0] = 1'b0;
  assign \A[14][248] [0] = 1'b0;
  assign \A[14][249] [2] = 1'b0;
  assign \A[14][250] [4] = 1'b0;
  assign \A[14][250] [3] = 1'b0;
  assign \A[14][250] [2] = 1'b0;
  assign \A[14][250] [1] = 1'b0;
  assign \A[14][253] [4] = 1'b0;
  assign \A[14][253] [3] = 1'b0;
  assign \A[14][253] [2] = 1'b0;
  assign \A[14][253] [0] = 1'b0;
  assign \A[14][254] [4] = 1'b0;
  assign \A[14][254] [3] = 1'b0;
  assign \A[14][254] [2] = 1'b0;
  assign \A[14][255] [4] = 1'b0;
  assign \A[14][255] [3] = 1'b0;
  assign \A[14][255] [2] = 1'b0;
  assign \A[15][0] [4] = 1'b0;
  assign \A[15][0] [3] = 1'b0;
  assign \A[15][0] [2] = 1'b0;
  assign \A[15][0] [1] = 1'b0;
  assign \A[15][0] [0] = 1'b0;
  assign \A[15][1] [4] = 1'b0;
  assign \A[15][1] [3] = 1'b0;
  assign \A[15][1] [2] = 1'b0;
  assign \A[15][1] [0] = 1'b0;
  assign \A[15][2] [4] = 1'b0;
  assign \A[15][2] [3] = 1'b0;
  assign \A[15][2] [2] = 1'b0;
  assign \A[15][2] [0] = 1'b0;
  assign \A[15][3] [0] = 1'b0;
  assign \A[15][4] [4] = 1'b0;
  assign \A[15][4] [3] = 1'b0;
  assign \A[15][4] [2] = 1'b0;
  assign \A[15][4] [1] = 1'b0;
  assign \A[15][4] [0] = 1'b0;
  assign \A[15][5] [4] = 1'b0;
  assign \A[15][5] [3] = 1'b0;
  assign \A[15][5] [2] = 1'b0;
  assign \A[15][5] [1] = 1'b0;
  assign \A[15][5] [0] = 1'b0;
  assign \A[15][6] [4] = 1'b0;
  assign \A[15][6] [3] = 1'b0;
  assign \A[15][6] [2] = 1'b0;
  assign \A[15][6] [1] = 1'b0;
  assign \A[15][6] [0] = 1'b0;
  assign \A[15][8] [4] = 1'b0;
  assign \A[15][8] [3] = 1'b0;
  assign \A[15][8] [2] = 1'b0;
  assign \A[15][8] [1] = 1'b0;
  assign \A[15][8] [0] = 1'b0;
  assign \A[15][9] [4] = 1'b0;
  assign \A[15][9] [3] = 1'b0;
  assign \A[15][9] [2] = 1'b0;
  assign \A[15][9] [1] = 1'b0;
  assign \A[15][10] [0] = 1'b0;
  assign \A[15][13] [0] = 1'b0;
  assign \A[15][14] [4] = 1'b0;
  assign \A[15][14] [3] = 1'b0;
  assign \A[15][14] [2] = 1'b0;
  assign \A[15][14] [1] = 1'b0;
  assign \A[15][14] [0] = 1'b0;
  assign \A[15][20] [4] = 1'b0;
  assign \A[15][20] [3] = 1'b0;
  assign \A[15][20] [2] = 1'b0;
  assign \A[15][20] [1] = 1'b0;
  assign \A[15][21] [0] = 1'b0;
  assign \A[15][22] [0] = 1'b0;
  assign \A[15][23] [4] = 1'b0;
  assign \A[15][23] [3] = 1'b0;
  assign \A[15][23] [2] = 1'b0;
  assign \A[15][23] [1] = 1'b0;
  assign \A[15][23] [0] = 1'b0;
  assign \A[15][25] [4] = 1'b0;
  assign \A[15][25] [3] = 1'b0;
  assign \A[15][25] [2] = 1'b0;
  assign \A[15][25] [1] = 1'b0;
  assign \A[15][25] [0] = 1'b0;
  assign \A[15][26] [0] = 1'b0;
  assign \A[15][28] [0] = 1'b0;
  assign \A[15][29] [4] = 1'b0;
  assign \A[15][29] [3] = 1'b0;
  assign \A[15][29] [2] = 1'b0;
  assign \A[15][29] [1] = 1'b0;
  assign \A[15][30] [4] = 1'b0;
  assign \A[15][30] [3] = 1'b0;
  assign \A[15][30] [2] = 1'b0;
  assign \A[15][30] [1] = 1'b0;
  assign \A[15][30] [0] = 1'b0;
  assign \A[15][32] [0] = 1'b0;
  assign \A[15][33] [4] = 1'b0;
  assign \A[15][33] [3] = 1'b0;
  assign \A[15][33] [2] = 1'b0;
  assign \A[15][33] [1] = 1'b0;
  assign \A[15][34] [0] = 1'b0;
  assign \A[15][35] [4] = 1'b0;
  assign \A[15][35] [3] = 1'b0;
  assign \A[15][35] [2] = 1'b0;
  assign \A[15][35] [1] = 1'b0;
  assign \A[15][36] [0] = 1'b0;
  assign \A[15][38] [0] = 1'b0;
  assign \A[15][39] [4] = 1'b0;
  assign \A[15][39] [3] = 1'b0;
  assign \A[15][39] [2] = 1'b0;
  assign \A[15][39] [1] = 1'b0;
  assign \A[15][39] [0] = 1'b0;
  assign \A[15][40] [4] = 1'b0;
  assign \A[15][40] [3] = 1'b0;
  assign \A[15][40] [2] = 1'b0;
  assign \A[15][40] [1] = 1'b0;
  assign \A[15][41] [4] = 1'b0;
  assign \A[15][41] [3] = 1'b0;
  assign \A[15][41] [2] = 1'b0;
  assign \A[15][41] [1] = 1'b0;
  assign \A[15][42] [1] = 1'b0;
  assign \A[15][43] [0] = 1'b0;
  assign \A[15][46] [4] = 1'b0;
  assign \A[15][46] [3] = 1'b0;
  assign \A[15][46] [2] = 1'b0;
  assign \A[15][46] [1] = 1'b0;
  assign \A[15][46] [0] = 1'b0;
  assign \A[15][47] [4] = 1'b0;
  assign \A[15][47] [3] = 1'b0;
  assign \A[15][47] [2] = 1'b0;
  assign \A[15][47] [0] = 1'b0;
  assign \A[15][48] [4] = 1'b0;
  assign \A[15][48] [3] = 1'b0;
  assign \A[15][48] [2] = 1'b0;
  assign \A[15][48] [1] = 1'b0;
  assign \A[15][48] [0] = 1'b0;
  assign \A[15][49] [4] = 1'b0;
  assign \A[15][49] [3] = 1'b0;
  assign \A[15][49] [2] = 1'b0;
  assign \A[15][49] [0] = 1'b0;
  assign \A[15][50] [4] = 1'b0;
  assign \A[15][50] [3] = 1'b0;
  assign \A[15][50] [2] = 1'b0;
  assign \A[15][50] [0] = 1'b0;
  assign \A[15][51] [4] = 1'b0;
  assign \A[15][51] [3] = 1'b0;
  assign \A[15][51] [2] = 1'b0;
  assign \A[15][51] [1] = 1'b0;
  assign \A[15][51] [0] = 1'b0;
  assign \A[15][54] [4] = 1'b0;
  assign \A[15][54] [3] = 1'b0;
  assign \A[15][54] [2] = 1'b0;
  assign \A[15][54] [0] = 1'b0;
  assign \A[15][56] [4] = 1'b0;
  assign \A[15][56] [3] = 1'b0;
  assign \A[15][56] [2] = 1'b0;
  assign \A[15][56] [1] = 1'b0;
  assign \A[15][57] [4] = 1'b0;
  assign \A[15][57] [3] = 1'b0;
  assign \A[15][57] [2] = 1'b0;
  assign \A[15][57] [1] = 1'b0;
  assign \A[15][58] [4] = 1'b0;
  assign \A[15][58] [3] = 1'b0;
  assign \A[15][58] [1] = 1'b0;
  assign \A[15][58] [0] = 1'b0;
  assign \A[15][60] [4] = 1'b0;
  assign \A[15][60] [3] = 1'b0;
  assign \A[15][60] [2] = 1'b0;
  assign \A[15][60] [1] = 1'b0;
  assign \A[15][61] [0] = 1'b0;
  assign \A[15][62] [4] = 1'b0;
  assign \A[15][62] [3] = 1'b0;
  assign \A[15][62] [2] = 1'b0;
  assign \A[15][62] [1] = 1'b0;
  assign \A[15][62] [0] = 1'b0;
  assign \A[15][63] [4] = 1'b0;
  assign \A[15][63] [3] = 1'b0;
  assign \A[15][63] [2] = 1'b0;
  assign \A[15][63] [1] = 1'b0;
  assign \A[15][63] [0] = 1'b0;
  assign \A[15][65] [4] = 1'b0;
  assign \A[15][65] [3] = 1'b0;
  assign \A[15][65] [2] = 1'b0;
  assign \A[15][65] [1] = 1'b0;
  assign \A[15][66] [4] = 1'b0;
  assign \A[15][66] [3] = 1'b0;
  assign \A[15][66] [2] = 1'b0;
  assign \A[15][66] [1] = 1'b0;
  assign \A[15][66] [0] = 1'b0;
  assign \A[15][67] [4] = 1'b0;
  assign \A[15][67] [3] = 1'b0;
  assign \A[15][67] [2] = 1'b0;
  assign \A[15][67] [1] = 1'b0;
  assign \A[15][68] [4] = 1'b0;
  assign \A[15][68] [3] = 1'b0;
  assign \A[15][68] [2] = 1'b0;
  assign \A[15][68] [1] = 1'b0;
  assign \A[15][68] [0] = 1'b0;
  assign \A[15][70] [4] = 1'b0;
  assign \A[15][70] [3] = 1'b0;
  assign \A[15][70] [2] = 1'b0;
  assign \A[15][70] [0] = 1'b0;
  assign \A[15][71] [4] = 1'b0;
  assign \A[15][71] [3] = 1'b0;
  assign \A[15][71] [2] = 1'b0;
  assign \A[15][71] [0] = 1'b0;
  assign \A[15][73] [0] = 1'b0;
  assign \A[15][74] [1] = 1'b0;
  assign \A[15][75] [4] = 1'b0;
  assign \A[15][75] [3] = 1'b0;
  assign \A[15][75] [2] = 1'b0;
  assign \A[15][75] [1] = 1'b0;
  assign \A[15][77] [4] = 1'b0;
  assign \A[15][77] [3] = 1'b0;
  assign \A[15][77] [2] = 1'b0;
  assign \A[15][77] [1] = 1'b0;
  assign \A[15][77] [0] = 1'b0;
  assign \A[15][78] [4] = 1'b0;
  assign \A[15][78] [3] = 1'b0;
  assign \A[15][78] [2] = 1'b0;
  assign \A[15][78] [1] = 1'b0;
  assign \A[15][79] [4] = 1'b0;
  assign \A[15][79] [3] = 1'b0;
  assign \A[15][79] [2] = 1'b0;
  assign \A[15][79] [1] = 1'b0;
  assign \A[15][79] [0] = 1'b0;
  assign \A[15][80] [4] = 1'b0;
  assign \A[15][80] [3] = 1'b0;
  assign \A[15][80] [2] = 1'b0;
  assign \A[15][80] [1] = 1'b0;
  assign \A[15][81] [1] = 1'b0;
  assign \A[15][82] [4] = 1'b0;
  assign \A[15][82] [3] = 1'b0;
  assign \A[15][82] [2] = 1'b0;
  assign \A[15][82] [1] = 1'b0;
  assign \A[15][82] [0] = 1'b0;
  assign \A[15][83] [0] = 1'b0;
  assign \A[15][84] [4] = 1'b0;
  assign \A[15][84] [3] = 1'b0;
  assign \A[15][84] [2] = 1'b0;
  assign \A[15][84] [1] = 1'b0;
  assign \A[15][84] [0] = 1'b0;
  assign \A[15][85] [4] = 1'b0;
  assign \A[15][85] [3] = 1'b0;
  assign \A[15][85] [2] = 1'b0;
  assign \A[15][85] [0] = 1'b0;
  assign \A[15][86] [0] = 1'b0;
  assign \A[15][87] [4] = 1'b0;
  assign \A[15][87] [3] = 1'b0;
  assign \A[15][87] [2] = 1'b0;
  assign \A[15][87] [1] = 1'b0;
  assign \A[15][87] [0] = 1'b0;
  assign \A[15][88] [4] = 1'b0;
  assign \A[15][88] [3] = 1'b0;
  assign \A[15][88] [2] = 1'b0;
  assign \A[15][88] [1] = 1'b0;
  assign \A[15][88] [0] = 1'b0;
  assign \A[15][89] [4] = 1'b0;
  assign \A[15][89] [3] = 1'b0;
  assign \A[15][89] [2] = 1'b0;
  assign \A[15][89] [1] = 1'b0;
  assign \A[15][89] [0] = 1'b0;
  assign \A[15][90] [4] = 1'b0;
  assign \A[15][90] [3] = 1'b0;
  assign \A[15][90] [2] = 1'b0;
  assign \A[15][90] [1] = 1'b0;
  assign \A[15][90] [0] = 1'b0;
  assign \A[15][91] [4] = 1'b0;
  assign \A[15][91] [3] = 1'b0;
  assign \A[15][91] [2] = 1'b0;
  assign \A[15][91] [1] = 1'b0;
  assign \A[15][92] [4] = 1'b0;
  assign \A[15][92] [3] = 1'b0;
  assign \A[15][92] [2] = 1'b0;
  assign \A[15][92] [1] = 1'b0;
  assign \A[15][93] [0] = 1'b0;
  assign \A[15][94] [4] = 1'b0;
  assign \A[15][94] [3] = 1'b0;
  assign \A[15][94] [2] = 1'b0;
  assign \A[15][94] [1] = 1'b0;
  assign \A[15][95] [4] = 1'b0;
  assign \A[15][95] [3] = 1'b0;
  assign \A[15][95] [2] = 1'b0;
  assign \A[15][95] [1] = 1'b0;
  assign \A[15][95] [0] = 1'b0;
  assign \A[15][96] [4] = 1'b0;
  assign \A[15][96] [3] = 1'b0;
  assign \A[15][96] [2] = 1'b0;
  assign \A[15][96] [1] = 1'b0;
  assign \A[15][98] [4] = 1'b0;
  assign \A[15][98] [3] = 1'b0;
  assign \A[15][98] [2] = 1'b0;
  assign \A[15][98] [1] = 1'b0;
  assign \A[15][99] [4] = 1'b0;
  assign \A[15][99] [3] = 1'b0;
  assign \A[15][99] [2] = 1'b0;
  assign \A[15][100] [1] = 1'b0;
  assign \A[15][101] [4] = 1'b0;
  assign \A[15][101] [3] = 1'b0;
  assign \A[15][101] [2] = 1'b0;
  assign \A[15][102] [4] = 1'b0;
  assign \A[15][102] [3] = 1'b0;
  assign \A[15][102] [2] = 1'b0;
  assign \A[15][102] [1] = 1'b0;
  assign \A[15][104] [4] = 1'b0;
  assign \A[15][104] [3] = 1'b0;
  assign \A[15][104] [2] = 1'b0;
  assign \A[15][104] [1] = 1'b0;
  assign \A[15][105] [0] = 1'b0;
  assign \A[15][106] [4] = 1'b0;
  assign \A[15][106] [3] = 1'b0;
  assign \A[15][106] [2] = 1'b0;
  assign \A[15][106] [1] = 1'b0;
  assign \A[15][109] [4] = 1'b0;
  assign \A[15][109] [3] = 1'b0;
  assign \A[15][109] [2] = 1'b0;
  assign \A[15][109] [1] = 1'b0;
  assign \A[15][110] [4] = 1'b0;
  assign \A[15][110] [3] = 1'b0;
  assign \A[15][110] [2] = 1'b0;
  assign \A[15][110] [1] = 1'b0;
  assign \A[15][110] [0] = 1'b0;
  assign \A[15][111] [0] = 1'b0;
  assign \A[15][112] [4] = 1'b0;
  assign \A[15][112] [3] = 1'b0;
  assign \A[15][112] [2] = 1'b0;
  assign \A[15][112] [1] = 1'b0;
  assign \A[15][112] [0] = 1'b0;
  assign \A[15][115] [4] = 1'b0;
  assign \A[15][115] [3] = 1'b0;
  assign \A[15][115] [2] = 1'b0;
  assign \A[15][115] [0] = 1'b0;
  assign \A[15][116] [4] = 1'b0;
  assign \A[15][116] [3] = 1'b0;
  assign \A[15][116] [2] = 1'b0;
  assign \A[15][116] [1] = 1'b0;
  assign \A[15][116] [0] = 1'b0;
  assign \A[15][118] [4] = 1'b0;
  assign \A[15][118] [3] = 1'b0;
  assign \A[15][118] [2] = 1'b0;
  assign \A[15][118] [1] = 1'b0;
  assign \A[15][120] [4] = 1'b0;
  assign \A[15][120] [3] = 1'b0;
  assign \A[15][120] [2] = 1'b0;
  assign \A[15][120] [1] = 1'b0;
  assign \A[15][120] [0] = 1'b0;
  assign \A[15][121] [4] = 1'b0;
  assign \A[15][121] [3] = 1'b0;
  assign \A[15][121] [2] = 1'b0;
  assign \A[15][121] [1] = 1'b0;
  assign \A[15][121] [0] = 1'b0;
  assign \A[15][122] [4] = 1'b0;
  assign \A[15][122] [3] = 1'b0;
  assign \A[15][122] [2] = 1'b0;
  assign \A[15][122] [1] = 1'b0;
  assign \A[15][122] [0] = 1'b0;
  assign \A[15][123] [4] = 1'b0;
  assign \A[15][123] [3] = 1'b0;
  assign \A[15][123] [2] = 1'b0;
  assign \A[15][123] [1] = 1'b0;
  assign \A[15][123] [0] = 1'b0;
  assign \A[15][124] [4] = 1'b0;
  assign \A[15][124] [3] = 1'b0;
  assign \A[15][124] [2] = 1'b0;
  assign \A[15][124] [1] = 1'b0;
  assign \A[15][124] [0] = 1'b0;
  assign \A[15][125] [1] = 1'b0;
  assign \A[15][126] [4] = 1'b0;
  assign \A[15][126] [3] = 1'b0;
  assign \A[15][126] [2] = 1'b0;
  assign \A[15][126] [0] = 1'b0;
  assign \A[15][127] [4] = 1'b0;
  assign \A[15][127] [3] = 1'b0;
  assign \A[15][127] [2] = 1'b0;
  assign \A[15][127] [1] = 1'b0;
  assign \A[15][129] [4] = 1'b0;
  assign \A[15][129] [3] = 1'b0;
  assign \A[15][129] [2] = 1'b0;
  assign \A[15][129] [1] = 1'b0;
  assign \A[15][129] [0] = 1'b0;
  assign \A[15][132] [0] = 1'b0;
  assign \A[15][134] [0] = 1'b0;
  assign \A[15][135] [0] = 1'b0;
  assign \A[15][136] [4] = 1'b0;
  assign \A[15][136] [3] = 1'b0;
  assign \A[15][136] [2] = 1'b0;
  assign \A[15][136] [1] = 1'b0;
  assign \A[15][136] [0] = 1'b0;
  assign \A[15][137] [4] = 1'b0;
  assign \A[15][137] [3] = 1'b0;
  assign \A[15][137] [2] = 1'b0;
  assign \A[15][137] [1] = 1'b0;
  assign \A[15][138] [4] = 1'b0;
  assign \A[15][138] [3] = 1'b0;
  assign \A[15][138] [2] = 1'b0;
  assign \A[15][138] [1] = 1'b0;
  assign \A[15][138] [0] = 1'b0;
  assign \A[15][139] [0] = 1'b0;
  assign \A[15][140] [4] = 1'b0;
  assign \A[15][140] [3] = 1'b0;
  assign \A[15][140] [2] = 1'b0;
  assign \A[15][141] [4] = 1'b0;
  assign \A[15][141] [3] = 1'b0;
  assign \A[15][141] [2] = 1'b0;
  assign \A[15][141] [1] = 1'b0;
  assign \A[15][142] [4] = 1'b0;
  assign \A[15][142] [3] = 1'b0;
  assign \A[15][142] [2] = 1'b0;
  assign \A[15][142] [1] = 1'b0;
  assign \A[15][142] [0] = 1'b0;
  assign \A[15][143] [0] = 1'b0;
  assign \A[15][145] [0] = 1'b0;
  assign \A[15][146] [4] = 1'b0;
  assign \A[15][146] [3] = 1'b0;
  assign \A[15][146] [2] = 1'b0;
  assign \A[15][146] [1] = 1'b0;
  assign \A[15][147] [4] = 1'b0;
  assign \A[15][147] [3] = 1'b0;
  assign \A[15][147] [2] = 1'b0;
  assign \A[15][147] [1] = 1'b0;
  assign \A[15][147] [0] = 1'b0;
  assign \A[15][149] [4] = 1'b0;
  assign \A[15][149] [3] = 1'b0;
  assign \A[15][149] [2] = 1'b0;
  assign \A[15][149] [1] = 1'b0;
  assign \A[15][149] [0] = 1'b0;
  assign \A[15][150] [4] = 1'b0;
  assign \A[15][150] [3] = 1'b0;
  assign \A[15][150] [2] = 1'b0;
  assign \A[15][150] [1] = 1'b0;
  assign \A[15][150] [0] = 1'b0;
  assign \A[15][152] [0] = 1'b0;
  assign \A[15][154] [1] = 1'b0;
  assign \A[15][155] [4] = 1'b0;
  assign \A[15][155] [3] = 1'b0;
  assign \A[15][155] [2] = 1'b0;
  assign \A[15][155] [1] = 1'b0;
  assign \A[15][155] [0] = 1'b0;
  assign \A[15][156] [4] = 1'b0;
  assign \A[15][156] [3] = 1'b0;
  assign \A[15][156] [1] = 1'b0;
  assign \A[15][156] [0] = 1'b0;
  assign \A[15][157] [4] = 1'b0;
  assign \A[15][157] [3] = 1'b0;
  assign \A[15][157] [2] = 1'b0;
  assign \A[15][157] [1] = 1'b0;
  assign \A[15][157] [0] = 1'b0;
  assign \A[15][159] [4] = 1'b0;
  assign \A[15][159] [3] = 1'b0;
  assign \A[15][159] [2] = 1'b0;
  assign \A[15][159] [1] = 1'b0;
  assign \A[15][160] [4] = 1'b0;
  assign \A[15][160] [3] = 1'b0;
  assign \A[15][160] [2] = 1'b0;
  assign \A[15][160] [1] = 1'b0;
  assign \A[15][161] [4] = 1'b0;
  assign \A[15][161] [3] = 1'b0;
  assign \A[15][161] [2] = 1'b0;
  assign \A[15][161] [1] = 1'b0;
  assign \A[15][161] [0] = 1'b0;
  assign \A[15][164] [4] = 1'b0;
  assign \A[15][164] [3] = 1'b0;
  assign \A[15][164] [2] = 1'b0;
  assign \A[15][164] [1] = 1'b0;
  assign \A[15][164] [0] = 1'b0;
  assign \A[15][165] [4] = 1'b0;
  assign \A[15][165] [3] = 1'b0;
  assign \A[15][165] [2] = 1'b0;
  assign \A[15][165] [1] = 1'b0;
  assign \A[15][166] [4] = 1'b0;
  assign \A[15][166] [3] = 1'b0;
  assign \A[15][166] [2] = 1'b0;
  assign \A[15][166] [1] = 1'b0;
  assign \A[15][167] [4] = 1'b0;
  assign \A[15][167] [3] = 1'b0;
  assign \A[15][167] [2] = 1'b0;
  assign \A[15][167] [1] = 1'b0;
  assign \A[15][167] [0] = 1'b0;
  assign \A[15][168] [4] = 1'b0;
  assign \A[15][168] [3] = 1'b0;
  assign \A[15][168] [2] = 1'b0;
  assign \A[15][168] [1] = 1'b0;
  assign \A[15][168] [0] = 1'b0;
  assign \A[15][169] [1] = 1'b0;
  assign \A[15][170] [4] = 1'b0;
  assign \A[15][170] [3] = 1'b0;
  assign \A[15][170] [2] = 1'b0;
  assign \A[15][170] [0] = 1'b0;
  assign \A[15][171] [4] = 1'b0;
  assign \A[15][171] [3] = 1'b0;
  assign \A[15][171] [2] = 1'b0;
  assign \A[15][171] [1] = 1'b0;
  assign \A[15][171] [0] = 1'b0;
  assign \A[15][172] [0] = 1'b0;
  assign \A[15][173] [1] = 1'b0;
  assign \A[15][175] [4] = 1'b0;
  assign \A[15][175] [3] = 1'b0;
  assign \A[15][175] [2] = 1'b0;
  assign \A[15][175] [1] = 1'b0;
  assign \A[15][177] [0] = 1'b0;
  assign \A[15][178] [0] = 1'b0;
  assign \A[15][180] [4] = 1'b0;
  assign \A[15][180] [3] = 1'b0;
  assign \A[15][180] [2] = 1'b0;
  assign \A[15][180] [1] = 1'b0;
  assign \A[15][181] [0] = 1'b0;
  assign \A[15][183] [4] = 1'b0;
  assign \A[15][183] [3] = 1'b0;
  assign \A[15][183] [2] = 1'b0;
  assign \A[15][183] [1] = 1'b0;
  assign \A[15][183] [0] = 1'b0;
  assign \A[15][184] [4] = 1'b0;
  assign \A[15][184] [3] = 1'b0;
  assign \A[15][184] [2] = 1'b0;
  assign \A[15][184] [1] = 1'b0;
  assign \A[15][185] [4] = 1'b0;
  assign \A[15][185] [3] = 1'b0;
  assign \A[15][185] [2] = 1'b0;
  assign \A[15][185] [1] = 1'b0;
  assign \A[15][187] [4] = 1'b0;
  assign \A[15][187] [3] = 1'b0;
  assign \A[15][187] [2] = 1'b0;
  assign \A[15][187] [1] = 1'b0;
  assign \A[15][187] [0] = 1'b0;
  assign \A[15][188] [4] = 1'b0;
  assign \A[15][188] [3] = 1'b0;
  assign \A[15][188] [2] = 1'b0;
  assign \A[15][188] [1] = 1'b0;
  assign \A[15][189] [1] = 1'b0;
  assign \A[15][190] [4] = 1'b0;
  assign \A[15][190] [3] = 1'b0;
  assign \A[15][190] [2] = 1'b0;
  assign \A[15][190] [0] = 1'b0;
  assign \A[15][191] [4] = 1'b0;
  assign \A[15][191] [3] = 1'b0;
  assign \A[15][191] [2] = 1'b0;
  assign \A[15][191] [1] = 1'b0;
  assign \A[15][191] [0] = 1'b0;
  assign \A[15][192] [4] = 1'b0;
  assign \A[15][192] [3] = 1'b0;
  assign \A[15][192] [2] = 1'b0;
  assign \A[15][192] [1] = 1'b0;
  assign \A[15][193] [4] = 1'b0;
  assign \A[15][193] [3] = 1'b0;
  assign \A[15][193] [2] = 1'b0;
  assign \A[15][193] [1] = 1'b0;
  assign \A[15][194] [4] = 1'b0;
  assign \A[15][194] [3] = 1'b0;
  assign \A[15][194] [2] = 1'b0;
  assign \A[15][194] [1] = 1'b0;
  assign \A[15][194] [0] = 1'b0;
  assign \A[15][197] [4] = 1'b0;
  assign \A[15][197] [3] = 1'b0;
  assign \A[15][197] [2] = 1'b0;
  assign \A[15][197] [1] = 1'b0;
  assign \A[15][197] [0] = 1'b0;
  assign \A[15][198] [0] = 1'b0;
  assign \A[15][201] [4] = 1'b0;
  assign \A[15][201] [3] = 1'b0;
  assign \A[15][201] [2] = 1'b0;
  assign \A[15][201] [1] = 1'b0;
  assign \A[15][201] [0] = 1'b0;
  assign \A[15][202] [4] = 1'b0;
  assign \A[15][202] [3] = 1'b0;
  assign \A[15][202] [2] = 1'b0;
  assign \A[15][202] [0] = 1'b0;
  assign \A[15][203] [4] = 1'b0;
  assign \A[15][203] [3] = 1'b0;
  assign \A[15][203] [2] = 1'b0;
  assign \A[15][203] [1] = 1'b0;
  assign \A[15][203] [0] = 1'b0;
  assign \A[15][207] [4] = 1'b0;
  assign \A[15][207] [3] = 1'b0;
  assign \A[15][207] [2] = 1'b0;
  assign \A[15][207] [1] = 1'b0;
  assign \A[15][207] [0] = 1'b0;
  assign \A[15][208] [4] = 1'b0;
  assign \A[15][208] [3] = 1'b0;
  assign \A[15][208] [2] = 1'b0;
  assign \A[15][208] [1] = 1'b0;
  assign \A[15][208] [0] = 1'b0;
  assign \A[15][209] [4] = 1'b0;
  assign \A[15][209] [3] = 1'b0;
  assign \A[15][209] [2] = 1'b0;
  assign \A[15][209] [1] = 1'b0;
  assign \A[15][210] [4] = 1'b0;
  assign \A[15][210] [3] = 1'b0;
  assign \A[15][210] [2] = 1'b0;
  assign \A[15][210] [1] = 1'b0;
  assign \A[15][211] [4] = 1'b0;
  assign \A[15][211] [3] = 1'b0;
  assign \A[15][211] [2] = 1'b0;
  assign \A[15][211] [1] = 1'b0;
  assign \A[15][211] [0] = 1'b0;
  assign \A[15][213] [0] = 1'b0;
  assign \A[15][214] [4] = 1'b0;
  assign \A[15][214] [3] = 1'b0;
  assign \A[15][214] [2] = 1'b0;
  assign \A[15][214] [0] = 1'b0;
  assign \A[15][216] [4] = 1'b0;
  assign \A[15][216] [3] = 1'b0;
  assign \A[15][216] [2] = 1'b0;
  assign \A[15][216] [1] = 1'b0;
  assign \A[15][217] [4] = 1'b0;
  assign \A[15][217] [3] = 1'b0;
  assign \A[15][217] [2] = 1'b0;
  assign \A[15][217] [1] = 1'b0;
  assign \A[15][219] [4] = 1'b0;
  assign \A[15][219] [3] = 1'b0;
  assign \A[15][219] [2] = 1'b0;
  assign \A[15][219] [1] = 1'b0;
  assign \A[15][220] [0] = 1'b0;
  assign \A[15][222] [0] = 1'b0;
  assign \A[15][224] [4] = 1'b0;
  assign \A[15][224] [3] = 1'b0;
  assign \A[15][224] [2] = 1'b0;
  assign \A[15][224] [1] = 1'b0;
  assign \A[15][224] [0] = 1'b0;
  assign \A[15][225] [4] = 1'b0;
  assign \A[15][225] [3] = 1'b0;
  assign \A[15][225] [2] = 1'b0;
  assign \A[15][226] [4] = 1'b0;
  assign \A[15][226] [3] = 1'b0;
  assign \A[15][226] [2] = 1'b0;
  assign \A[15][226] [1] = 1'b0;
  assign \A[15][226] [0] = 1'b0;
  assign \A[15][227] [4] = 1'b0;
  assign \A[15][227] [3] = 1'b0;
  assign \A[15][227] [2] = 1'b0;
  assign \A[15][227] [0] = 1'b0;
  assign \A[15][228] [4] = 1'b0;
  assign \A[15][228] [3] = 1'b0;
  assign \A[15][228] [2] = 1'b0;
  assign \A[15][228] [1] = 1'b0;
  assign \A[15][228] [0] = 1'b0;
  assign \A[15][230] [4] = 1'b0;
  assign \A[15][230] [3] = 1'b0;
  assign \A[15][230] [2] = 1'b0;
  assign \A[15][230] [1] = 1'b0;
  assign \A[15][230] [0] = 1'b0;
  assign \A[15][231] [4] = 1'b0;
  assign \A[15][231] [3] = 1'b0;
  assign \A[15][231] [2] = 1'b0;
  assign \A[15][231] [1] = 1'b0;
  assign \A[15][231] [0] = 1'b0;
  assign \A[15][233] [4] = 1'b0;
  assign \A[15][233] [3] = 1'b0;
  assign \A[15][233] [2] = 1'b0;
  assign \A[15][233] [1] = 1'b0;
  assign \A[15][235] [4] = 1'b0;
  assign \A[15][235] [3] = 1'b0;
  assign \A[15][235] [2] = 1'b0;
  assign \A[15][235] [1] = 1'b0;
  assign \A[15][235] [0] = 1'b0;
  assign \A[15][236] [4] = 1'b0;
  assign \A[15][236] [3] = 1'b0;
  assign \A[15][236] [2] = 1'b0;
  assign \A[15][236] [1] = 1'b0;
  assign \A[15][236] [0] = 1'b0;
  assign \A[15][237] [4] = 1'b0;
  assign \A[15][237] [3] = 1'b0;
  assign \A[15][237] [2] = 1'b0;
  assign \A[15][237] [0] = 1'b0;
  assign \A[15][239] [4] = 1'b0;
  assign \A[15][239] [3] = 1'b0;
  assign \A[15][239] [2] = 1'b0;
  assign \A[15][239] [1] = 1'b0;
  assign \A[15][239] [0] = 1'b0;
  assign \A[15][240] [4] = 1'b0;
  assign \A[15][240] [3] = 1'b0;
  assign \A[15][240] [2] = 1'b0;
  assign \A[15][240] [0] = 1'b0;
  assign \A[15][241] [4] = 1'b0;
  assign \A[15][241] [3] = 1'b0;
  assign \A[15][241] [2] = 1'b0;
  assign \A[15][241] [1] = 1'b0;
  assign \A[15][242] [4] = 1'b0;
  assign \A[15][242] [3] = 1'b0;
  assign \A[15][242] [2] = 1'b0;
  assign \A[15][242] [0] = 1'b0;
  assign \A[15][243] [0] = 1'b0;
  assign \A[15][244] [4] = 1'b0;
  assign \A[15][244] [3] = 1'b0;
  assign \A[15][244] [2] = 1'b0;
  assign \A[15][244] [1] = 1'b0;
  assign \A[15][244] [0] = 1'b0;
  assign \A[15][246] [4] = 1'b0;
  assign \A[15][246] [3] = 1'b0;
  assign \A[15][246] [2] = 1'b0;
  assign \A[15][246] [1] = 1'b0;
  assign \A[15][247] [4] = 1'b0;
  assign \A[15][247] [3] = 1'b0;
  assign \A[15][247] [2] = 1'b0;
  assign \A[15][247] [1] = 1'b0;
  assign \A[15][247] [0] = 1'b0;
  assign \A[15][248] [1] = 1'b0;
  assign \A[15][249] [4] = 1'b0;
  assign \A[15][249] [3] = 1'b0;
  assign \A[15][249] [2] = 1'b0;
  assign \A[15][249] [1] = 1'b0;
  assign \A[15][249] [0] = 1'b0;
  assign \A[15][250] [4] = 1'b0;
  assign \A[15][250] [3] = 1'b0;
  assign \A[15][250] [2] = 1'b0;
  assign \A[15][250] [0] = 1'b0;
  assign \A[15][251] [4] = 1'b0;
  assign \A[15][251] [3] = 1'b0;
  assign \A[15][251] [2] = 1'b0;
  assign \A[15][251] [1] = 1'b0;
  assign \A[15][252] [4] = 1'b0;
  assign \A[15][252] [3] = 1'b0;
  assign \A[15][252] [2] = 1'b0;
  assign \A[15][252] [1] = 1'b0;
  assign \A[15][253] [4] = 1'b0;
  assign \A[15][253] [3] = 1'b0;
  assign \A[15][253] [2] = 1'b0;
  assign \A[15][253] [1] = 1'b0;
  assign \A[15][253] [0] = 1'b0;
  assign \A[15][254] [4] = 1'b0;
  assign \A[15][254] [3] = 1'b0;
  assign \A[15][254] [2] = 1'b0;
  assign \A[15][254] [1] = 1'b0;
  assign \A[16][0] [4] = 1'b0;
  assign \A[16][0] [3] = 1'b0;
  assign \A[16][0] [2] = 1'b0;
  assign \A[16][0] [1] = 1'b0;
  assign \A[16][0] [0] = 1'b0;
  assign \A[16][1] [4] = 1'b0;
  assign \A[16][1] [3] = 1'b0;
  assign \A[16][1] [2] = 1'b0;
  assign \A[16][1] [1] = 1'b0;
  assign \A[16][1] [0] = 1'b0;
  assign \A[16][3] [0] = 1'b0;
  assign \A[16][4] [4] = 1'b0;
  assign \A[16][4] [3] = 1'b0;
  assign \A[16][4] [2] = 1'b0;
  assign \A[16][4] [1] = 1'b0;
  assign \A[16][4] [0] = 1'b0;
  assign \A[16][5] [4] = 1'b0;
  assign \A[16][5] [3] = 1'b0;
  assign \A[16][5] [2] = 1'b0;
  assign \A[16][5] [0] = 1'b0;
  assign \A[16][6] [0] = 1'b0;
  assign \A[16][9] [4] = 1'b0;
  assign \A[16][9] [3] = 1'b0;
  assign \A[16][9] [2] = 1'b0;
  assign \A[16][9] [0] = 1'b0;
  assign \A[16][11] [4] = 1'b0;
  assign \A[16][11] [3] = 1'b0;
  assign \A[16][11] [2] = 1'b0;
  assign \A[16][11] [1] = 1'b0;
  assign \A[16][11] [0] = 1'b0;
  assign \A[16][12] [4] = 1'b0;
  assign \A[16][12] [3] = 1'b0;
  assign \A[16][12] [2] = 1'b0;
  assign \A[16][13] [0] = 1'b0;
  assign \A[16][14] [1] = 1'b0;
  assign \A[16][14] [0] = 1'b0;
  assign \A[16][15] [0] = 1'b0;
  assign \A[16][16] [4] = 1'b0;
  assign \A[16][16] [3] = 1'b0;
  assign \A[16][16] [2] = 1'b0;
  assign \A[16][17] [4] = 1'b0;
  assign \A[16][17] [3] = 1'b0;
  assign \A[16][17] [2] = 1'b0;
  assign \A[16][17] [1] = 1'b0;
  assign \A[16][17] [0] = 1'b0;
  assign \A[16][19] [1] = 1'b0;
  assign \A[16][21] [0] = 1'b0;
  assign \A[16][23] [0] = 1'b0;
  assign \A[16][25] [4] = 1'b0;
  assign \A[16][25] [3] = 1'b0;
  assign \A[16][25] [2] = 1'b0;
  assign \A[16][25] [1] = 1'b0;
  assign \A[16][25] [0] = 1'b0;
  assign \A[16][27] [4] = 1'b0;
  assign \A[16][27] [3] = 1'b0;
  assign \A[16][27] [2] = 1'b0;
  assign \A[16][27] [1] = 1'b0;
  assign \A[16][28] [1] = 1'b0;
  assign \A[16][29] [4] = 1'b0;
  assign \A[16][29] [3] = 1'b0;
  assign \A[16][29] [2] = 1'b0;
  assign \A[16][29] [1] = 1'b0;
  assign \A[16][29] [0] = 1'b0;
  assign \A[16][30] [4] = 1'b0;
  assign \A[16][30] [3] = 1'b0;
  assign \A[16][30] [2] = 1'b0;
  assign \A[16][30] [1] = 1'b0;
  assign \A[16][31] [4] = 1'b0;
  assign \A[16][31] [3] = 1'b0;
  assign \A[16][31] [2] = 1'b0;
  assign \A[16][31] [1] = 1'b0;
  assign \A[16][31] [0] = 1'b0;
  assign \A[16][32] [4] = 1'b0;
  assign \A[16][32] [3] = 1'b0;
  assign \A[16][32] [2] = 1'b0;
  assign \A[16][32] [1] = 1'b0;
  assign \A[16][32] [0] = 1'b0;
  assign \A[16][33] [4] = 1'b0;
  assign \A[16][33] [3] = 1'b0;
  assign \A[16][33] [2] = 1'b0;
  assign \A[16][33] [1] = 1'b0;
  assign \A[16][34] [4] = 1'b0;
  assign \A[16][34] [3] = 1'b0;
  assign \A[16][34] [2] = 1'b0;
  assign \A[16][34] [1] = 1'b0;
  assign \A[16][34] [0] = 1'b0;
  assign \A[16][35] [4] = 1'b0;
  assign \A[16][35] [3] = 1'b0;
  assign \A[16][35] [2] = 1'b0;
  assign \A[16][35] [1] = 1'b0;
  assign \A[16][35] [0] = 1'b0;
  assign \A[16][36] [0] = 1'b0;
  assign \A[16][38] [4] = 1'b0;
  assign \A[16][38] [3] = 1'b0;
  assign \A[16][38] [2] = 1'b0;
  assign \A[16][38] [1] = 1'b0;
  assign \A[16][38] [0] = 1'b0;
  assign \A[16][39] [4] = 1'b0;
  assign \A[16][39] [3] = 1'b0;
  assign \A[16][39] [2] = 1'b0;
  assign \A[16][39] [1] = 1'b0;
  assign \A[16][40] [4] = 1'b0;
  assign \A[16][40] [3] = 1'b0;
  assign \A[16][40] [2] = 1'b0;
  assign \A[16][40] [1] = 1'b0;
  assign \A[16][40] [0] = 1'b0;
  assign \A[16][41] [0] = 1'b0;
  assign \A[16][43] [0] = 1'b0;
  assign \A[16][44] [0] = 1'b0;
  assign \A[16][45] [0] = 1'b0;
  assign \A[16][46] [4] = 1'b0;
  assign \A[16][46] [3] = 1'b0;
  assign \A[16][46] [2] = 1'b0;
  assign \A[16][46] [0] = 1'b0;
  assign \A[16][47] [0] = 1'b0;
  assign \A[16][48] [4] = 1'b0;
  assign \A[16][48] [3] = 1'b0;
  assign \A[16][48] [2] = 1'b0;
  assign \A[16][48] [1] = 1'b0;
  assign \A[16][48] [0] = 1'b0;
  assign \A[16][49] [4] = 1'b0;
  assign \A[16][49] [3] = 1'b0;
  assign \A[16][49] [2] = 1'b0;
  assign \A[16][49] [1] = 1'b0;
  assign \A[16][49] [0] = 1'b0;
  assign \A[16][50] [4] = 1'b0;
  assign \A[16][50] [3] = 1'b0;
  assign \A[16][50] [2] = 1'b0;
  assign \A[16][50] [1] = 1'b0;
  assign \A[16][51] [4] = 1'b0;
  assign \A[16][51] [3] = 1'b0;
  assign \A[16][51] [2] = 1'b0;
  assign \A[16][51] [0] = 1'b0;
  assign \A[16][52] [4] = 1'b0;
  assign \A[16][52] [3] = 1'b0;
  assign \A[16][52] [2] = 1'b0;
  assign \A[16][52] [1] = 1'b0;
  assign \A[16][54] [4] = 1'b0;
  assign \A[16][54] [3] = 1'b0;
  assign \A[16][54] [2] = 1'b0;
  assign \A[16][54] [0] = 1'b0;
  assign \A[16][57] [4] = 1'b0;
  assign \A[16][57] [3] = 1'b0;
  assign \A[16][57] [2] = 1'b0;
  assign \A[16][57] [1] = 1'b0;
  assign \A[16][60] [4] = 1'b0;
  assign \A[16][60] [3] = 1'b0;
  assign \A[16][60] [2] = 1'b0;
  assign \A[16][60] [1] = 1'b0;
  assign \A[16][63] [4] = 1'b0;
  assign \A[16][63] [3] = 1'b0;
  assign \A[16][63] [2] = 1'b0;
  assign \A[16][63] [1] = 1'b0;
  assign \A[16][64] [4] = 1'b0;
  assign \A[16][64] [3] = 1'b0;
  assign \A[16][64] [2] = 1'b0;
  assign \A[16][64] [1] = 1'b0;
  assign \A[16][65] [0] = 1'b0;
  assign \A[16][66] [0] = 1'b0;
  assign \A[16][68] [4] = 1'b0;
  assign \A[16][68] [3] = 1'b0;
  assign \A[16][68] [2] = 1'b0;
  assign \A[16][68] [1] = 1'b0;
  assign \A[16][68] [0] = 1'b0;
  assign \A[16][70] [4] = 1'b0;
  assign \A[16][70] [3] = 1'b0;
  assign \A[16][70] [2] = 1'b0;
  assign \A[16][70] [1] = 1'b0;
  assign \A[16][70] [0] = 1'b0;
  assign \A[16][72] [4] = 1'b0;
  assign \A[16][72] [3] = 1'b0;
  assign \A[16][72] [2] = 1'b0;
  assign \A[16][72] [1] = 1'b0;
  assign \A[16][72] [0] = 1'b0;
  assign \A[16][74] [4] = 1'b0;
  assign \A[16][74] [3] = 1'b0;
  assign \A[16][74] [2] = 1'b0;
  assign \A[16][75] [4] = 1'b0;
  assign \A[16][75] [3] = 1'b0;
  assign \A[16][75] [2] = 1'b0;
  assign \A[16][75] [1] = 1'b0;
  assign \A[16][75] [0] = 1'b0;
  assign \A[16][76] [4] = 1'b0;
  assign \A[16][76] [3] = 1'b0;
  assign \A[16][76] [1] = 1'b0;
  assign \A[16][78] [4] = 1'b0;
  assign \A[16][78] [3] = 1'b0;
  assign \A[16][78] [2] = 1'b0;
  assign \A[16][78] [1] = 1'b0;
  assign \A[16][80] [0] = 1'b0;
  assign \A[16][81] [4] = 1'b0;
  assign \A[16][81] [3] = 1'b0;
  assign \A[16][81] [2] = 1'b0;
  assign \A[16][81] [1] = 1'b0;
  assign \A[16][83] [1] = 1'b0;
  assign \A[16][85] [1] = 1'b0;
  assign \A[16][87] [4] = 1'b0;
  assign \A[16][87] [3] = 1'b0;
  assign \A[16][87] [2] = 1'b0;
  assign \A[16][87] [0] = 1'b0;
  assign \A[16][88] [4] = 1'b0;
  assign \A[16][88] [3] = 1'b0;
  assign \A[16][88] [2] = 1'b0;
  assign \A[16][88] [1] = 1'b0;
  assign \A[16][89] [0] = 1'b0;
  assign \A[16][90] [4] = 1'b0;
  assign \A[16][90] [3] = 1'b0;
  assign \A[16][90] [2] = 1'b0;
  assign \A[16][90] [1] = 1'b0;
  assign \A[16][90] [0] = 1'b0;
  assign \A[16][91] [0] = 1'b0;
  assign \A[16][92] [4] = 1'b0;
  assign \A[16][92] [3] = 1'b0;
  assign \A[16][92] [2] = 1'b0;
  assign \A[16][92] [0] = 1'b0;
  assign \A[16][93] [4] = 1'b0;
  assign \A[16][93] [3] = 1'b0;
  assign \A[16][93] [2] = 1'b0;
  assign \A[16][93] [1] = 1'b0;
  assign \A[16][95] [4] = 1'b0;
  assign \A[16][95] [3] = 1'b0;
  assign \A[16][95] [2] = 1'b0;
  assign \A[16][95] [1] = 1'b0;
  assign \A[16][95] [0] = 1'b0;
  assign \A[16][96] [4] = 1'b0;
  assign \A[16][96] [3] = 1'b0;
  assign \A[16][96] [2] = 1'b0;
  assign \A[16][96] [1] = 1'b0;
  assign \A[16][97] [4] = 1'b0;
  assign \A[16][97] [3] = 1'b0;
  assign \A[16][97] [2] = 1'b0;
  assign \A[16][97] [1] = 1'b0;
  assign \A[16][98] [4] = 1'b0;
  assign \A[16][98] [3] = 1'b0;
  assign \A[16][98] [2] = 1'b0;
  assign \A[16][98] [1] = 1'b0;
  assign \A[16][98] [0] = 1'b0;
  assign \A[16][99] [4] = 1'b0;
  assign \A[16][99] [3] = 1'b0;
  assign \A[16][99] [2] = 1'b0;
  assign \A[16][99] [1] = 1'b0;
  assign \A[16][100] [4] = 1'b0;
  assign \A[16][100] [3] = 1'b0;
  assign \A[16][100] [2] = 1'b0;
  assign \A[16][100] [1] = 1'b0;
  assign \A[16][101] [4] = 1'b0;
  assign \A[16][101] [3] = 1'b0;
  assign \A[16][101] [2] = 1'b0;
  assign \A[16][101] [0] = 1'b0;
  assign \A[16][102] [1] = 1'b0;
  assign \A[16][102] [0] = 1'b0;
  assign \A[16][104] [4] = 1'b0;
  assign \A[16][104] [3] = 1'b0;
  assign \A[16][104] [2] = 1'b0;
  assign \A[16][104] [1] = 1'b0;
  assign \A[16][104] [0] = 1'b0;
  assign \A[16][105] [4] = 1'b0;
  assign \A[16][105] [3] = 1'b0;
  assign \A[16][105] [2] = 1'b0;
  assign \A[16][105] [1] = 1'b0;
  assign \A[16][106] [0] = 1'b0;
  assign \A[16][107] [4] = 1'b0;
  assign \A[16][107] [3] = 1'b0;
  assign \A[16][107] [2] = 1'b0;
  assign \A[16][108] [4] = 1'b0;
  assign \A[16][108] [3] = 1'b0;
  assign \A[16][108] [2] = 1'b0;
  assign \A[16][108] [1] = 1'b0;
  assign \A[16][109] [4] = 1'b0;
  assign \A[16][109] [3] = 1'b0;
  assign \A[16][109] [2] = 1'b0;
  assign \A[16][109] [1] = 1'b0;
  assign \A[16][110] [4] = 1'b0;
  assign \A[16][110] [3] = 1'b0;
  assign \A[16][110] [2] = 1'b0;
  assign \A[16][110] [1] = 1'b0;
  assign \A[16][111] [0] = 1'b0;
  assign \A[16][112] [4] = 1'b0;
  assign \A[16][112] [3] = 1'b0;
  assign \A[16][112] [2] = 1'b0;
  assign \A[16][112] [1] = 1'b0;
  assign \A[16][112] [0] = 1'b0;
  assign \A[16][113] [4] = 1'b0;
  assign \A[16][113] [3] = 1'b0;
  assign \A[16][113] [2] = 1'b0;
  assign \A[16][113] [1] = 1'b0;
  assign \A[16][113] [0] = 1'b0;
  assign \A[16][116] [4] = 1'b0;
  assign \A[16][116] [3] = 1'b0;
  assign \A[16][116] [2] = 1'b0;
  assign \A[16][116] [1] = 1'b0;
  assign \A[16][116] [0] = 1'b0;
  assign \A[16][117] [4] = 1'b0;
  assign \A[16][117] [3] = 1'b0;
  assign \A[16][117] [2] = 1'b0;
  assign \A[16][117] [0] = 1'b0;
  assign \A[16][118] [0] = 1'b0;
  assign \A[16][119] [4] = 1'b0;
  assign \A[16][119] [3] = 1'b0;
  assign \A[16][119] [2] = 1'b0;
  assign \A[16][119] [1] = 1'b0;
  assign \A[16][119] [0] = 1'b0;
  assign \A[16][121] [4] = 1'b0;
  assign \A[16][121] [3] = 1'b0;
  assign \A[16][121] [2] = 1'b0;
  assign \A[16][121] [1] = 1'b0;
  assign \A[16][122] [4] = 1'b0;
  assign \A[16][122] [3] = 1'b0;
  assign \A[16][122] [2] = 1'b0;
  assign \A[16][122] [1] = 1'b0;
  assign \A[16][122] [0] = 1'b0;
  assign \A[16][124] [4] = 1'b0;
  assign \A[16][124] [3] = 1'b0;
  assign \A[16][124] [2] = 1'b0;
  assign \A[16][125] [4] = 1'b0;
  assign \A[16][125] [3] = 1'b0;
  assign \A[16][125] [2] = 1'b0;
  assign \A[16][125] [1] = 1'b0;
  assign \A[16][126] [0] = 1'b0;
  assign \A[16][128] [4] = 1'b0;
  assign \A[16][128] [3] = 1'b0;
  assign \A[16][128] [2] = 1'b0;
  assign \A[16][128] [1] = 1'b0;
  assign \A[16][128] [0] = 1'b0;
  assign \A[16][129] [4] = 1'b0;
  assign \A[16][129] [3] = 1'b0;
  assign \A[16][129] [2] = 1'b0;
  assign \A[16][129] [0] = 1'b0;
  assign \A[16][130] [4] = 1'b0;
  assign \A[16][130] [3] = 1'b0;
  assign \A[16][130] [2] = 1'b0;
  assign \A[16][130] [0] = 1'b0;
  assign \A[16][132] [4] = 1'b0;
  assign \A[16][132] [3] = 1'b0;
  assign \A[16][132] [2] = 1'b0;
  assign \A[16][132] [1] = 1'b0;
  assign \A[16][133] [4] = 1'b0;
  assign \A[16][133] [3] = 1'b0;
  assign \A[16][133] [2] = 1'b0;
  assign \A[16][133] [1] = 1'b0;
  assign \A[16][133] [0] = 1'b0;
  assign \A[16][134] [4] = 1'b0;
  assign \A[16][134] [3] = 1'b0;
  assign \A[16][134] [2] = 1'b0;
  assign \A[16][134] [1] = 1'b0;
  assign \A[16][135] [0] = 1'b0;
  assign \A[16][136] [4] = 1'b0;
  assign \A[16][136] [3] = 1'b0;
  assign \A[16][136] [2] = 1'b0;
  assign \A[16][136] [1] = 1'b0;
  assign \A[16][136] [0] = 1'b0;
  assign \A[16][137] [4] = 1'b0;
  assign \A[16][137] [3] = 1'b0;
  assign \A[16][137] [2] = 1'b0;
  assign \A[16][137] [1] = 1'b0;
  assign \A[16][137] [0] = 1'b0;
  assign \A[16][138] [4] = 1'b0;
  assign \A[16][138] [3] = 1'b0;
  assign \A[16][138] [2] = 1'b0;
  assign \A[16][138] [1] = 1'b0;
  assign \A[16][138] [0] = 1'b0;
  assign \A[16][139] [0] = 1'b0;
  assign \A[16][141] [0] = 1'b0;
  assign \A[16][144] [4] = 1'b0;
  assign \A[16][144] [3] = 1'b0;
  assign \A[16][144] [2] = 1'b0;
  assign \A[16][144] [1] = 1'b0;
  assign \A[16][144] [0] = 1'b0;
  assign \A[16][145] [4] = 1'b0;
  assign \A[16][145] [3] = 1'b0;
  assign \A[16][145] [2] = 1'b0;
  assign \A[16][145] [1] = 1'b0;
  assign \A[16][146] [4] = 1'b0;
  assign \A[16][146] [3] = 1'b0;
  assign \A[16][146] [2] = 1'b0;
  assign \A[16][146] [1] = 1'b0;
  assign \A[16][146] [0] = 1'b0;
  assign \A[16][147] [4] = 1'b0;
  assign \A[16][147] [3] = 1'b0;
  assign \A[16][147] [2] = 1'b0;
  assign \A[16][148] [4] = 1'b0;
  assign \A[16][148] [3] = 1'b0;
  assign \A[16][148] [2] = 1'b0;
  assign \A[16][148] [1] = 1'b0;
  assign \A[16][148] [0] = 1'b0;
  assign \A[16][149] [4] = 1'b0;
  assign \A[16][149] [3] = 1'b0;
  assign \A[16][149] [2] = 1'b0;
  assign \A[16][149] [1] = 1'b0;
  assign \A[16][149] [0] = 1'b0;
  assign \A[16][150] [4] = 1'b0;
  assign \A[16][150] [3] = 1'b0;
  assign \A[16][150] [2] = 1'b0;
  assign \A[16][150] [1] = 1'b0;
  assign \A[16][151] [1] = 1'b0;
  assign \A[16][152] [4] = 1'b0;
  assign \A[16][152] [3] = 1'b0;
  assign \A[16][152] [2] = 1'b0;
  assign \A[16][152] [1] = 1'b0;
  assign \A[16][153] [0] = 1'b0;
  assign \A[16][154] [4] = 1'b0;
  assign \A[16][154] [3] = 1'b0;
  assign \A[16][154] [2] = 1'b0;
  assign \A[16][154] [1] = 1'b0;
  assign \A[16][154] [0] = 1'b0;
  assign \A[16][155] [4] = 1'b0;
  assign \A[16][155] [3] = 1'b0;
  assign \A[16][155] [2] = 1'b0;
  assign \A[16][155] [1] = 1'b0;
  assign \A[16][157] [0] = 1'b0;
  assign \A[16][159] [0] = 1'b0;
  assign \A[16][160] [4] = 1'b0;
  assign \A[16][160] [3] = 1'b0;
  assign \A[16][160] [2] = 1'b0;
  assign \A[16][160] [0] = 1'b0;
  assign \A[16][161] [4] = 1'b0;
  assign \A[16][161] [3] = 1'b0;
  assign \A[16][161] [2] = 1'b0;
  assign \A[16][161] [1] = 1'b0;
  assign \A[16][161] [0] = 1'b0;
  assign \A[16][162] [4] = 1'b0;
  assign \A[16][162] [3] = 1'b0;
  assign \A[16][162] [2] = 1'b0;
  assign \A[16][162] [0] = 1'b0;
  assign \A[16][163] [4] = 1'b0;
  assign \A[16][163] [3] = 1'b0;
  assign \A[16][163] [2] = 1'b0;
  assign \A[16][163] [1] = 1'b0;
  assign \A[16][163] [0] = 1'b0;
  assign \A[16][164] [4] = 1'b0;
  assign \A[16][164] [3] = 1'b0;
  assign \A[16][164] [2] = 1'b0;
  assign \A[16][164] [0] = 1'b0;
  assign \A[16][166] [0] = 1'b0;
  assign \A[16][167] [4] = 1'b0;
  assign \A[16][167] [3] = 1'b0;
  assign \A[16][167] [2] = 1'b0;
  assign \A[16][167] [0] = 1'b0;
  assign \A[16][168] [4] = 1'b0;
  assign \A[16][168] [3] = 1'b0;
  assign \A[16][168] [2] = 1'b0;
  assign \A[16][168] [0] = 1'b0;
  assign \A[16][169] [4] = 1'b0;
  assign \A[16][169] [3] = 1'b0;
  assign \A[16][169] [2] = 1'b0;
  assign \A[16][169] [1] = 1'b0;
  assign \A[16][169] [0] = 1'b0;
  assign \A[16][170] [4] = 1'b0;
  assign \A[16][170] [3] = 1'b0;
  assign \A[16][170] [2] = 1'b0;
  assign \A[16][170] [0] = 1'b0;
  assign \A[16][172] [4] = 1'b0;
  assign \A[16][172] [3] = 1'b0;
  assign \A[16][172] [2] = 1'b0;
  assign \A[16][172] [1] = 1'b0;
  assign \A[16][172] [0] = 1'b0;
  assign \A[16][173] [0] = 1'b0;
  assign \A[16][175] [4] = 1'b0;
  assign \A[16][175] [3] = 1'b0;
  assign \A[16][175] [2] = 1'b0;
  assign \A[16][175] [0] = 1'b0;
  assign \A[16][176] [4] = 1'b0;
  assign \A[16][176] [3] = 1'b0;
  assign \A[16][176] [2] = 1'b0;
  assign \A[16][176] [1] = 1'b0;
  assign \A[16][177] [4] = 1'b0;
  assign \A[16][177] [3] = 1'b0;
  assign \A[16][177] [2] = 1'b0;
  assign \A[16][177] [0] = 1'b0;
  assign \A[16][178] [0] = 1'b0;
  assign \A[16][179] [4] = 1'b0;
  assign \A[16][179] [3] = 1'b0;
  assign \A[16][179] [2] = 1'b0;
  assign \A[16][179] [1] = 1'b0;
  assign \A[16][180] [4] = 1'b0;
  assign \A[16][180] [3] = 1'b0;
  assign \A[16][180] [2] = 1'b0;
  assign \A[16][180] [1] = 1'b0;
  assign \A[16][180] [0] = 1'b0;
  assign \A[16][181] [4] = 1'b0;
  assign \A[16][181] [3] = 1'b0;
  assign \A[16][181] [2] = 1'b0;
  assign \A[16][182] [4] = 1'b0;
  assign \A[16][182] [3] = 1'b0;
  assign \A[16][182] [2] = 1'b0;
  assign \A[16][182] [1] = 1'b0;
  assign \A[16][183] [4] = 1'b0;
  assign \A[16][183] [3] = 1'b0;
  assign \A[16][183] [2] = 1'b0;
  assign \A[16][183] [1] = 1'b0;
  assign \A[16][183] [0] = 1'b0;
  assign \A[16][184] [0] = 1'b0;
  assign \A[16][186] [4] = 1'b0;
  assign \A[16][186] [3] = 1'b0;
  assign \A[16][186] [2] = 1'b0;
  assign \A[16][186] [1] = 1'b0;
  assign \A[16][187] [4] = 1'b0;
  assign \A[16][187] [3] = 1'b0;
  assign \A[16][187] [2] = 1'b0;
  assign \A[16][187] [1] = 1'b0;
  assign \A[16][187] [0] = 1'b0;
  assign \A[16][188] [4] = 1'b0;
  assign \A[16][188] [3] = 1'b0;
  assign \A[16][188] [2] = 1'b0;
  assign \A[16][188] [1] = 1'b0;
  assign \A[16][188] [0] = 1'b0;
  assign \A[16][190] [0] = 1'b0;
  assign \A[16][191] [4] = 1'b0;
  assign \A[16][191] [3] = 1'b0;
  assign \A[16][191] [2] = 1'b0;
  assign \A[16][191] [1] = 1'b0;
  assign \A[16][193] [4] = 1'b0;
  assign \A[16][193] [3] = 1'b0;
  assign \A[16][193] [2] = 1'b0;
  assign \A[16][193] [1] = 1'b0;
  assign \A[16][193] [0] = 1'b0;
  assign \A[16][194] [0] = 1'b0;
  assign \A[16][195] [4] = 1'b0;
  assign \A[16][195] [3] = 1'b0;
  assign \A[16][195] [2] = 1'b0;
  assign \A[16][195] [0] = 1'b0;
  assign \A[16][196] [0] = 1'b0;
  assign \A[16][197] [4] = 1'b0;
  assign \A[16][197] [3] = 1'b0;
  assign \A[16][197] [2] = 1'b0;
  assign \A[16][197] [1] = 1'b0;
  assign \A[16][197] [0] = 1'b0;
  assign \A[16][199] [4] = 1'b0;
  assign \A[16][199] [3] = 1'b0;
  assign \A[16][199] [2] = 1'b0;
  assign \A[16][199] [1] = 1'b0;
  assign \A[16][200] [0] = 1'b0;
  assign \A[16][201] [4] = 1'b0;
  assign \A[16][201] [3] = 1'b0;
  assign \A[16][201] [2] = 1'b0;
  assign \A[16][201] [1] = 1'b0;
  assign \A[16][201] [0] = 1'b0;
  assign \A[16][202] [1] = 1'b0;
  assign \A[16][204] [0] = 1'b0;
  assign \A[16][207] [4] = 1'b0;
  assign \A[16][207] [3] = 1'b0;
  assign \A[16][207] [2] = 1'b0;
  assign \A[16][207] [1] = 1'b0;
  assign \A[16][207] [0] = 1'b0;
  assign \A[16][208] [4] = 1'b0;
  assign \A[16][208] [3] = 1'b0;
  assign \A[16][208] [2] = 1'b0;
  assign \A[16][208] [1] = 1'b0;
  assign \A[16][208] [0] = 1'b0;
  assign \A[16][209] [4] = 1'b0;
  assign \A[16][209] [3] = 1'b0;
  assign \A[16][209] [2] = 1'b0;
  assign \A[16][209] [1] = 1'b0;
  assign \A[16][210] [4] = 1'b0;
  assign \A[16][210] [3] = 1'b0;
  assign \A[16][210] [2] = 1'b0;
  assign \A[16][210] [1] = 1'b0;
  assign \A[16][210] [0] = 1'b0;
  assign \A[16][211] [4] = 1'b0;
  assign \A[16][211] [3] = 1'b0;
  assign \A[16][211] [2] = 1'b0;
  assign \A[16][211] [0] = 1'b0;
  assign \A[16][212] [4] = 1'b0;
  assign \A[16][212] [3] = 1'b0;
  assign \A[16][212] [2] = 1'b0;
  assign \A[16][212] [1] = 1'b0;
  assign \A[16][213] [1] = 1'b0;
  assign \A[16][214] [4] = 1'b0;
  assign \A[16][214] [3] = 1'b0;
  assign \A[16][214] [2] = 1'b0;
  assign \A[16][214] [0] = 1'b0;
  assign \A[16][215] [4] = 1'b0;
  assign \A[16][215] [3] = 1'b0;
  assign \A[16][215] [2] = 1'b0;
  assign \A[16][215] [1] = 1'b0;
  assign \A[16][216] [0] = 1'b0;
  assign \A[16][218] [0] = 1'b0;
  assign \A[16][219] [4] = 1'b0;
  assign \A[16][219] [3] = 1'b0;
  assign \A[16][219] [2] = 1'b0;
  assign \A[16][219] [1] = 1'b0;
  assign \A[16][219] [0] = 1'b0;
  assign \A[16][220] [4] = 1'b0;
  assign \A[16][220] [3] = 1'b0;
  assign \A[16][220] [2] = 1'b0;
  assign \A[16][220] [1] = 1'b0;
  assign \A[16][221] [4] = 1'b0;
  assign \A[16][221] [3] = 1'b0;
  assign \A[16][221] [2] = 1'b0;
  assign \A[16][221] [1] = 1'b0;
  assign \A[16][221] [0] = 1'b0;
  assign \A[16][223] [0] = 1'b0;
  assign \A[16][224] [4] = 1'b0;
  assign \A[16][224] [3] = 1'b0;
  assign \A[16][224] [2] = 1'b0;
  assign \A[16][224] [1] = 1'b0;
  assign \A[16][224] [0] = 1'b0;
  assign \A[16][225] [4] = 1'b0;
  assign \A[16][225] [3] = 1'b0;
  assign \A[16][225] [2] = 1'b0;
  assign \A[16][225] [1] = 1'b0;
  assign \A[16][225] [0] = 1'b0;
  assign \A[16][226] [4] = 1'b0;
  assign \A[16][226] [3] = 1'b0;
  assign \A[16][226] [2] = 1'b0;
  assign \A[16][226] [1] = 1'b0;
  assign \A[16][226] [0] = 1'b0;
  assign \A[16][227] [4] = 1'b0;
  assign \A[16][227] [3] = 1'b0;
  assign \A[16][227] [2] = 1'b0;
  assign \A[16][227] [1] = 1'b0;
  assign \A[16][227] [0] = 1'b0;
  assign \A[16][228] [4] = 1'b0;
  assign \A[16][228] [3] = 1'b0;
  assign \A[16][228] [2] = 1'b0;
  assign \A[16][228] [1] = 1'b0;
  assign \A[16][228] [0] = 1'b0;
  assign \A[16][229] [4] = 1'b0;
  assign \A[16][229] [3] = 1'b0;
  assign \A[16][229] [2] = 1'b0;
  assign \A[16][229] [1] = 1'b0;
  assign \A[16][229] [0] = 1'b0;
  assign \A[16][230] [4] = 1'b0;
  assign \A[16][230] [3] = 1'b0;
  assign \A[16][230] [2] = 1'b0;
  assign \A[16][230] [0] = 1'b0;
  assign \A[16][231] [4] = 1'b0;
  assign \A[16][231] [3] = 1'b0;
  assign \A[16][231] [2] = 1'b0;
  assign \A[16][231] [1] = 1'b0;
  assign \A[16][232] [4] = 1'b0;
  assign \A[16][232] [3] = 1'b0;
  assign \A[16][232] [2] = 1'b0;
  assign \A[16][232] [1] = 1'b0;
  assign \A[16][232] [0] = 1'b0;
  assign \A[16][233] [0] = 1'b0;
  assign \A[16][234] [4] = 1'b0;
  assign \A[16][234] [3] = 1'b0;
  assign \A[16][234] [2] = 1'b0;
  assign \A[16][234] [0] = 1'b0;
  assign \A[16][237] [4] = 1'b0;
  assign \A[16][237] [3] = 1'b0;
  assign \A[16][237] [2] = 1'b0;
  assign \A[16][237] [1] = 1'b0;
  assign \A[16][237] [0] = 1'b0;
  assign \A[16][238] [4] = 1'b0;
  assign \A[16][238] [3] = 1'b0;
  assign \A[16][238] [2] = 1'b0;
  assign \A[16][238] [1] = 1'b0;
  assign \A[16][238] [0] = 1'b0;
  assign \A[16][239] [1] = 1'b0;
  assign \A[16][240] [4] = 1'b0;
  assign \A[16][240] [3] = 1'b0;
  assign \A[16][240] [2] = 1'b0;
  assign \A[16][240] [1] = 1'b0;
  assign \A[16][240] [0] = 1'b0;
  assign \A[16][241] [0] = 1'b0;
  assign \A[16][242] [0] = 1'b0;
  assign \A[16][245] [0] = 1'b0;
  assign \A[16][246] [4] = 1'b0;
  assign \A[16][246] [3] = 1'b0;
  assign \A[16][246] [2] = 1'b0;
  assign \A[16][246] [1] = 1'b0;
  assign \A[16][247] [4] = 1'b0;
  assign \A[16][247] [3] = 1'b0;
  assign \A[16][247] [2] = 1'b0;
  assign \A[16][247] [1] = 1'b0;
  assign \A[16][248] [4] = 1'b0;
  assign \A[16][248] [3] = 1'b0;
  assign \A[16][248] [2] = 1'b0;
  assign \A[16][248] [1] = 1'b0;
  assign \A[16][248] [0] = 1'b0;
  assign \A[16][249] [4] = 1'b0;
  assign \A[16][249] [3] = 1'b0;
  assign \A[16][249] [2] = 1'b0;
  assign \A[16][249] [0] = 1'b0;
  assign \A[16][250] [4] = 1'b0;
  assign \A[16][250] [3] = 1'b0;
  assign \A[16][250] [2] = 1'b0;
  assign \A[16][250] [1] = 1'b0;
  assign \A[16][250] [0] = 1'b0;
  assign \A[16][251] [4] = 1'b0;
  assign \A[16][251] [3] = 1'b0;
  assign \A[16][251] [2] = 1'b0;
  assign \A[16][251] [0] = 1'b0;
  assign \A[16][252] [4] = 1'b0;
  assign \A[16][252] [3] = 1'b0;
  assign \A[16][252] [2] = 1'b0;
  assign \A[16][252] [0] = 1'b0;
  assign \A[16][253] [4] = 1'b0;
  assign \A[16][253] [3] = 1'b0;
  assign \A[16][253] [2] = 1'b0;
  assign \A[16][253] [1] = 1'b0;
  assign \A[16][254] [4] = 1'b0;
  assign \A[16][254] [3] = 1'b0;
  assign \A[16][254] [2] = 1'b0;
  assign \A[16][254] [1] = 1'b0;
  assign \A[16][255] [4] = 1'b0;
  assign \A[16][255] [3] = 1'b0;
  assign \A[16][255] [2] = 1'b0;
  assign \A[16][255] [1] = 1'b0;
  assign \A[16][255] [0] = 1'b0;
  assign \A[17][1] [1] = 1'b0;
  assign \A[17][2] [4] = 1'b0;
  assign \A[17][2] [3] = 1'b0;
  assign \A[17][2] [2] = 1'b0;
  assign \A[17][2] [0] = 1'b0;
  assign \A[17][3] [4] = 1'b0;
  assign \A[17][3] [3] = 1'b0;
  assign \A[17][3] [2] = 1'b0;
  assign \A[17][3] [1] = 1'b0;
  assign \A[17][4] [1] = 1'b0;
  assign \A[17][5] [1] = 1'b0;
  assign \A[17][5] [0] = 1'b0;
  assign \A[17][6] [4] = 1'b0;
  assign \A[17][6] [3] = 1'b0;
  assign \A[17][6] [2] = 1'b0;
  assign \A[17][6] [0] = 1'b0;
  assign \A[17][7] [4] = 1'b0;
  assign \A[17][7] [3] = 1'b0;
  assign \A[17][7] [0] = 1'b0;
  assign \A[17][8] [4] = 1'b0;
  assign \A[17][8] [3] = 1'b0;
  assign \A[17][8] [2] = 1'b0;
  assign \A[17][8] [1] = 1'b0;
  assign \A[17][8] [0] = 1'b0;
  assign \A[17][9] [0] = 1'b0;
  assign \A[17][10] [4] = 1'b0;
  assign \A[17][10] [3] = 1'b0;
  assign \A[17][10] [2] = 1'b0;
  assign \A[17][10] [1] = 1'b0;
  assign \A[17][10] [0] = 1'b0;
  assign \A[17][11] [1] = 1'b0;
  assign \A[17][12] [1] = 1'b0;
  assign \A[17][14] [0] = 1'b0;
  assign \A[17][15] [2] = 1'b0;
  assign \A[17][16] [4] = 1'b0;
  assign \A[17][16] [3] = 1'b0;
  assign \A[17][16] [2] = 1'b0;
  assign \A[17][16] [1] = 1'b0;
  assign \A[17][16] [0] = 1'b0;
  assign \A[17][17] [4] = 1'b0;
  assign \A[17][17] [3] = 1'b0;
  assign \A[17][17] [2] = 1'b0;
  assign \A[17][17] [1] = 1'b0;
  assign \A[17][17] [0] = 1'b0;
  assign \A[17][18] [4] = 1'b0;
  assign \A[17][18] [3] = 1'b0;
  assign \A[17][18] [2] = 1'b0;
  assign \A[17][18] [0] = 1'b0;
  assign \A[17][20] [4] = 1'b0;
  assign \A[17][20] [3] = 1'b0;
  assign \A[17][20] [2] = 1'b0;
  assign \A[17][20] [1] = 1'b0;
  assign \A[17][20] [0] = 1'b0;
  assign \A[17][21] [4] = 1'b0;
  assign \A[17][21] [3] = 1'b0;
  assign \A[17][21] [2] = 1'b0;
  assign \A[17][21] [1] = 1'b0;
  assign \A[17][22] [4] = 1'b0;
  assign \A[17][22] [3] = 1'b0;
  assign \A[17][22] [2] = 1'b0;
  assign \A[17][22] [0] = 1'b0;
  assign \A[17][23] [4] = 1'b0;
  assign \A[17][23] [3] = 1'b0;
  assign \A[17][23] [2] = 1'b0;
  assign \A[17][23] [1] = 1'b0;
  assign \A[17][24] [0] = 1'b0;
  assign \A[17][25] [4] = 1'b0;
  assign \A[17][25] [3] = 1'b0;
  assign \A[17][25] [2] = 1'b0;
  assign \A[17][25] [1] = 1'b0;
  assign \A[17][26] [4] = 1'b0;
  assign \A[17][26] [3] = 1'b0;
  assign \A[17][26] [2] = 1'b0;
  assign \A[17][26] [1] = 1'b0;
  assign \A[17][27] [4] = 1'b0;
  assign \A[17][27] [3] = 1'b0;
  assign \A[17][27] [2] = 1'b0;
  assign \A[17][27] [0] = 1'b0;
  assign \A[17][28] [0] = 1'b0;
  assign \A[17][29] [4] = 1'b0;
  assign \A[17][29] [3] = 1'b0;
  assign \A[17][29] [2] = 1'b0;
  assign \A[17][29] [1] = 1'b0;
  assign \A[17][30] [4] = 1'b0;
  assign \A[17][30] [3] = 1'b0;
  assign \A[17][30] [2] = 1'b0;
  assign \A[17][30] [0] = 1'b0;
  assign \A[17][34] [4] = 1'b0;
  assign \A[17][34] [3] = 1'b0;
  assign \A[17][34] [2] = 1'b0;
  assign \A[17][34] [1] = 1'b0;
  assign \A[17][34] [0] = 1'b0;
  assign \A[17][36] [0] = 1'b0;
  assign \A[17][38] [4] = 1'b0;
  assign \A[17][38] [3] = 1'b0;
  assign \A[17][38] [2] = 1'b0;
  assign \A[17][38] [1] = 1'b0;
  assign \A[17][38] [0] = 1'b0;
  assign \A[17][40] [4] = 1'b0;
  assign \A[17][40] [3] = 1'b0;
  assign \A[17][40] [2] = 1'b0;
  assign \A[17][40] [1] = 1'b0;
  assign \A[17][40] [0] = 1'b0;
  assign \A[17][42] [4] = 1'b0;
  assign \A[17][42] [3] = 1'b0;
  assign \A[17][42] [2] = 1'b0;
  assign \A[17][42] [0] = 1'b0;
  assign \A[17][43] [0] = 1'b0;
  assign \A[17][44] [4] = 1'b0;
  assign \A[17][44] [3] = 1'b0;
  assign \A[17][44] [2] = 1'b0;
  assign \A[17][44] [1] = 1'b0;
  assign \A[17][45] [1] = 1'b0;
  assign \A[17][46] [4] = 1'b0;
  assign \A[17][46] [3] = 1'b0;
  assign \A[17][46] [2] = 1'b0;
  assign \A[17][46] [1] = 1'b0;
  assign \A[17][47] [4] = 1'b0;
  assign \A[17][47] [3] = 1'b0;
  assign \A[17][47] [1] = 1'b0;
  assign \A[17][49] [1] = 1'b0;
  assign \A[17][50] [4] = 1'b0;
  assign \A[17][50] [3] = 1'b0;
  assign \A[17][50] [2] = 1'b0;
  assign \A[17][50] [1] = 1'b0;
  assign \A[17][51] [0] = 1'b0;
  assign \A[17][52] [0] = 1'b0;
  assign \A[17][53] [0] = 1'b0;
  assign \A[17][55] [4] = 1'b0;
  assign \A[17][55] [3] = 1'b0;
  assign \A[17][55] [1] = 1'b0;
  assign \A[17][55] [0] = 1'b0;
  assign \A[17][56] [4] = 1'b0;
  assign \A[17][56] [3] = 1'b0;
  assign \A[17][56] [2] = 1'b0;
  assign \A[17][56] [1] = 1'b0;
  assign \A[17][56] [0] = 1'b0;
  assign \A[17][57] [4] = 1'b0;
  assign \A[17][57] [3] = 1'b0;
  assign \A[17][57] [2] = 1'b0;
  assign \A[17][57] [0] = 1'b0;
  assign \A[17][59] [4] = 1'b0;
  assign \A[17][59] [3] = 1'b0;
  assign \A[17][59] [2] = 1'b0;
  assign \A[17][59] [1] = 1'b0;
  assign \A[17][60] [4] = 1'b0;
  assign \A[17][60] [3] = 1'b0;
  assign \A[17][60] [2] = 1'b0;
  assign \A[17][60] [1] = 1'b0;
  assign \A[17][62] [4] = 1'b0;
  assign \A[17][62] [3] = 1'b0;
  assign \A[17][62] [2] = 1'b0;
  assign \A[17][62] [0] = 1'b0;
  assign \A[17][63] [4] = 1'b0;
  assign \A[17][63] [3] = 1'b0;
  assign \A[17][63] [2] = 1'b0;
  assign \A[17][64] [4] = 1'b0;
  assign \A[17][64] [3] = 1'b0;
  assign \A[17][64] [2] = 1'b0;
  assign \A[17][64] [1] = 1'b0;
  assign \A[17][64] [0] = 1'b0;
  assign \A[17][65] [1] = 1'b0;
  assign \A[17][65] [0] = 1'b0;
  assign \A[17][66] [1] = 1'b0;
  assign \A[17][67] [4] = 1'b0;
  assign \A[17][67] [3] = 1'b0;
  assign \A[17][67] [2] = 1'b0;
  assign \A[17][67] [0] = 1'b0;
  assign \A[17][68] [4] = 1'b0;
  assign \A[17][68] [3] = 1'b0;
  assign \A[17][68] [2] = 1'b0;
  assign \A[17][68] [1] = 1'b0;
  assign \A[17][68] [0] = 1'b0;
  assign \A[17][69] [4] = 1'b0;
  assign \A[17][69] [3] = 1'b0;
  assign \A[17][69] [2] = 1'b0;
  assign \A[17][69] [1] = 1'b0;
  assign \A[17][70] [4] = 1'b0;
  assign \A[17][70] [3] = 1'b0;
  assign \A[17][70] [2] = 1'b0;
  assign \A[17][70] [1] = 1'b0;
  assign \A[17][71] [4] = 1'b0;
  assign \A[17][71] [3] = 1'b0;
  assign \A[17][71] [2] = 1'b0;
  assign \A[17][71] [1] = 1'b0;
  assign \A[17][72] [0] = 1'b0;
  assign \A[17][74] [4] = 1'b0;
  assign \A[17][74] [3] = 1'b0;
  assign \A[17][74] [2] = 1'b0;
  assign \A[17][74] [0] = 1'b0;
  assign \A[17][75] [4] = 1'b0;
  assign \A[17][75] [3] = 1'b0;
  assign \A[17][75] [2] = 1'b0;
  assign \A[17][75] [1] = 1'b0;
  assign \A[17][75] [0] = 1'b0;
  assign \A[17][76] [4] = 1'b0;
  assign \A[17][76] [3] = 1'b0;
  assign \A[17][76] [1] = 1'b0;
  assign \A[17][78] [4] = 1'b0;
  assign \A[17][78] [3] = 1'b0;
  assign \A[17][78] [1] = 1'b0;
  assign \A[17][78] [0] = 1'b0;
  assign \A[17][79] [4] = 1'b0;
  assign \A[17][79] [3] = 1'b0;
  assign \A[17][79] [2] = 1'b0;
  assign \A[17][79] [1] = 1'b0;
  assign \A[17][79] [0] = 1'b0;
  assign \A[17][81] [0] = 1'b0;
  assign \A[17][82] [4] = 1'b0;
  assign \A[17][82] [3] = 1'b0;
  assign \A[17][82] [2] = 1'b0;
  assign \A[17][82] [1] = 1'b0;
  assign \A[17][82] [0] = 1'b0;
  assign \A[17][84] [0] = 1'b0;
  assign \A[17][85] [4] = 1'b0;
  assign \A[17][85] [3] = 1'b0;
  assign \A[17][85] [2] = 1'b0;
  assign \A[17][85] [1] = 1'b0;
  assign \A[17][86] [4] = 1'b0;
  assign \A[17][86] [3] = 1'b0;
  assign \A[17][86] [2] = 1'b0;
  assign \A[17][86] [1] = 1'b0;
  assign \A[17][88] [4] = 1'b0;
  assign \A[17][88] [3] = 1'b0;
  assign \A[17][88] [1] = 1'b0;
  assign \A[17][88] [0] = 1'b0;
  assign \A[17][89] [4] = 1'b0;
  assign \A[17][89] [3] = 1'b0;
  assign \A[17][89] [2] = 1'b0;
  assign \A[17][89] [1] = 1'b0;
  assign \A[17][90] [4] = 1'b0;
  assign \A[17][90] [3] = 1'b0;
  assign \A[17][90] [2] = 1'b0;
  assign \A[17][90] [1] = 1'b0;
  assign \A[17][90] [0] = 1'b0;
  assign \A[17][91] [4] = 1'b0;
  assign \A[17][91] [3] = 1'b0;
  assign \A[17][91] [2] = 1'b0;
  assign \A[17][91] [1] = 1'b0;
  assign \A[17][91] [0] = 1'b0;
  assign \A[17][92] [0] = 1'b0;
  assign \A[17][93] [4] = 1'b0;
  assign \A[17][93] [3] = 1'b0;
  assign \A[17][93] [2] = 1'b0;
  assign \A[17][93] [1] = 1'b0;
  assign \A[17][94] [0] = 1'b0;
  assign \A[17][95] [4] = 1'b0;
  assign \A[17][95] [3] = 1'b0;
  assign \A[17][95] [2] = 1'b0;
  assign \A[17][95] [1] = 1'b0;
  assign \A[17][95] [0] = 1'b0;
  assign \A[17][96] [4] = 1'b0;
  assign \A[17][96] [3] = 1'b0;
  assign \A[17][96] [2] = 1'b0;
  assign \A[17][96] [1] = 1'b0;
  assign \A[17][96] [0] = 1'b0;
  assign \A[17][97] [4] = 1'b0;
  assign \A[17][97] [3] = 1'b0;
  assign \A[17][97] [2] = 1'b0;
  assign \A[17][97] [1] = 1'b0;
  assign \A[17][97] [0] = 1'b0;
  assign \A[17][98] [4] = 1'b0;
  assign \A[17][98] [3] = 1'b0;
  assign \A[17][98] [2] = 1'b0;
  assign \A[17][98] [0] = 1'b0;
  assign \A[17][99] [0] = 1'b0;
  assign \A[17][100] [4] = 1'b0;
  assign \A[17][100] [3] = 1'b0;
  assign \A[17][100] [2] = 1'b0;
  assign \A[17][100] [0] = 1'b0;
  assign \A[17][101] [1] = 1'b0;
  assign \A[17][102] [1] = 1'b0;
  assign \A[17][103] [4] = 1'b0;
  assign \A[17][103] [3] = 1'b0;
  assign \A[17][103] [2] = 1'b0;
  assign \A[17][103] [1] = 1'b0;
  assign \A[17][103] [0] = 1'b0;
  assign \A[17][104] [4] = 1'b0;
  assign \A[17][104] [3] = 1'b0;
  assign \A[17][104] [2] = 1'b0;
  assign \A[17][104] [0] = 1'b0;
  assign \A[17][106] [4] = 1'b0;
  assign \A[17][106] [3] = 1'b0;
  assign \A[17][106] [2] = 1'b0;
  assign \A[17][106] [1] = 1'b0;
  assign \A[17][106] [0] = 1'b0;
  assign \A[17][107] [4] = 1'b0;
  assign \A[17][107] [3] = 1'b0;
  assign \A[17][107] [2] = 1'b0;
  assign \A[17][107] [1] = 1'b0;
  assign \A[17][107] [0] = 1'b0;
  assign \A[17][108] [4] = 1'b0;
  assign \A[17][108] [3] = 1'b0;
  assign \A[17][108] [2] = 1'b0;
  assign \A[17][108] [0] = 1'b0;
  assign \A[17][109] [0] = 1'b0;
  assign \A[17][110] [0] = 1'b0;
  assign \A[17][111] [4] = 1'b0;
  assign \A[17][111] [3] = 1'b0;
  assign \A[17][111] [2] = 1'b0;
  assign \A[17][111] [1] = 1'b0;
  assign \A[17][111] [0] = 1'b0;
  assign \A[17][112] [1] = 1'b0;
  assign \A[17][112] [0] = 1'b0;
  assign \A[17][113] [0] = 1'b0;
  assign \A[17][114] [4] = 1'b0;
  assign \A[17][114] [3] = 1'b0;
  assign \A[17][114] [2] = 1'b0;
  assign \A[17][114] [1] = 1'b0;
  assign \A[17][114] [0] = 1'b0;
  assign \A[17][116] [4] = 1'b0;
  assign \A[17][116] [3] = 1'b0;
  assign \A[17][116] [2] = 1'b0;
  assign \A[17][116] [1] = 1'b0;
  assign \A[17][116] [0] = 1'b0;
  assign \A[17][117] [0] = 1'b0;
  assign \A[17][119] [4] = 1'b0;
  assign \A[17][119] [3] = 1'b0;
  assign \A[17][119] [2] = 1'b0;
  assign \A[17][119] [0] = 1'b0;
  assign \A[17][120] [1] = 1'b0;
  assign \A[17][121] [4] = 1'b0;
  assign \A[17][121] [3] = 1'b0;
  assign \A[17][121] [2] = 1'b0;
  assign \A[17][121] [1] = 1'b0;
  assign \A[17][123] [4] = 1'b0;
  assign \A[17][123] [3] = 1'b0;
  assign \A[17][123] [2] = 1'b0;
  assign \A[17][123] [1] = 1'b0;
  assign \A[17][123] [0] = 1'b0;
  assign \A[17][125] [1] = 1'b0;
  assign \A[17][126] [0] = 1'b0;
  assign \A[17][127] [0] = 1'b0;
  assign \A[17][128] [0] = 1'b0;
  assign \A[17][130] [4] = 1'b0;
  assign \A[17][130] [3] = 1'b0;
  assign \A[17][130] [2] = 1'b0;
  assign \A[17][130] [1] = 1'b0;
  assign \A[17][131] [4] = 1'b0;
  assign \A[17][131] [3] = 1'b0;
  assign \A[17][131] [2] = 1'b0;
  assign \A[17][131] [1] = 1'b0;
  assign \A[17][132] [4] = 1'b0;
  assign \A[17][132] [3] = 1'b0;
  assign \A[17][132] [2] = 1'b0;
  assign \A[17][132] [0] = 1'b0;
  assign \A[17][133] [0] = 1'b0;
  assign \A[17][135] [4] = 1'b0;
  assign \A[17][135] [3] = 1'b0;
  assign \A[17][135] [2] = 1'b0;
  assign \A[17][135] [1] = 1'b0;
  assign \A[17][135] [0] = 1'b0;
  assign \A[17][137] [4] = 1'b0;
  assign \A[17][137] [3] = 1'b0;
  assign \A[17][137] [2] = 1'b0;
  assign \A[17][137] [0] = 1'b0;
  assign \A[17][138] [4] = 1'b0;
  assign \A[17][138] [3] = 1'b0;
  assign \A[17][138] [2] = 1'b0;
  assign \A[17][138] [1] = 1'b0;
  assign \A[17][138] [0] = 1'b0;
  assign \A[17][139] [0] = 1'b0;
  assign \A[17][140] [4] = 1'b0;
  assign \A[17][140] [3] = 1'b0;
  assign \A[17][140] [2] = 1'b0;
  assign \A[17][140] [1] = 1'b0;
  assign \A[17][141] [4] = 1'b0;
  assign \A[17][141] [3] = 1'b0;
  assign \A[17][141] [2] = 1'b0;
  assign \A[17][141] [1] = 1'b0;
  assign \A[17][141] [0] = 1'b0;
  assign \A[17][143] [0] = 1'b0;
  assign \A[17][144] [4] = 1'b0;
  assign \A[17][144] [3] = 1'b0;
  assign \A[17][144] [2] = 1'b0;
  assign \A[17][144] [1] = 1'b0;
  assign \A[17][144] [0] = 1'b0;
  assign \A[17][145] [0] = 1'b0;
  assign \A[17][147] [4] = 1'b0;
  assign \A[17][147] [3] = 1'b0;
  assign \A[17][147] [2] = 1'b0;
  assign \A[17][147] [1] = 1'b0;
  assign \A[17][147] [0] = 1'b0;
  assign \A[17][148] [2] = 1'b0;
  assign \A[17][150] [4] = 1'b0;
  assign \A[17][150] [3] = 1'b0;
  assign \A[17][150] [2] = 1'b0;
  assign \A[17][150] [1] = 1'b0;
  assign \A[17][151] [4] = 1'b0;
  assign \A[17][151] [3] = 1'b0;
  assign \A[17][151] [2] = 1'b0;
  assign \A[17][151] [0] = 1'b0;
  assign \A[17][152] [0] = 1'b0;
  assign \A[17][153] [4] = 1'b0;
  assign \A[17][153] [3] = 1'b0;
  assign \A[17][153] [2] = 1'b0;
  assign \A[17][153] [1] = 1'b0;
  assign \A[17][155] [4] = 1'b0;
  assign \A[17][155] [3] = 1'b0;
  assign \A[17][155] [2] = 1'b0;
  assign \A[17][155] [1] = 1'b0;
  assign \A[17][155] [0] = 1'b0;
  assign \A[17][156] [1] = 1'b0;
  assign \A[17][156] [0] = 1'b0;
  assign \A[17][157] [4] = 1'b0;
  assign \A[17][157] [3] = 1'b0;
  assign \A[17][157] [2] = 1'b0;
  assign \A[17][157] [1] = 1'b0;
  assign \A[17][158] [0] = 1'b0;
  assign \A[17][160] [4] = 1'b0;
  assign \A[17][160] [3] = 1'b0;
  assign \A[17][160] [2] = 1'b0;
  assign \A[17][160] [1] = 1'b0;
  assign \A[17][160] [0] = 1'b0;
  assign \A[17][161] [4] = 1'b0;
  assign \A[17][161] [3] = 1'b0;
  assign \A[17][161] [2] = 1'b0;
  assign \A[17][161] [1] = 1'b0;
  assign \A[17][162] [4] = 1'b0;
  assign \A[17][162] [3] = 1'b0;
  assign \A[17][162] [2] = 1'b0;
  assign \A[17][162] [0] = 1'b0;
  assign \A[17][163] [4] = 1'b0;
  assign \A[17][163] [3] = 1'b0;
  assign \A[17][163] [2] = 1'b0;
  assign \A[17][164] [4] = 1'b0;
  assign \A[17][164] [3] = 1'b0;
  assign \A[17][164] [2] = 1'b0;
  assign \A[17][164] [1] = 1'b0;
  assign \A[17][165] [4] = 1'b0;
  assign \A[17][165] [3] = 1'b0;
  assign \A[17][165] [2] = 1'b0;
  assign \A[17][165] [0] = 1'b0;
  assign \A[17][167] [4] = 1'b0;
  assign \A[17][167] [3] = 1'b0;
  assign \A[17][167] [2] = 1'b0;
  assign \A[17][167] [1] = 1'b0;
  assign \A[17][167] [0] = 1'b0;
  assign \A[17][168] [0] = 1'b0;
  assign \A[17][170] [4] = 1'b0;
  assign \A[17][170] [3] = 1'b0;
  assign \A[17][170] [2] = 1'b0;
  assign \A[17][170] [1] = 1'b0;
  assign \A[17][171] [1] = 1'b0;
  assign \A[17][171] [0] = 1'b0;
  assign \A[17][172] [0] = 1'b0;
  assign \A[17][173] [4] = 1'b0;
  assign \A[17][173] [3] = 1'b0;
  assign \A[17][173] [2] = 1'b0;
  assign \A[17][173] [1] = 1'b0;
  assign \A[17][173] [0] = 1'b0;
  assign \A[17][174] [4] = 1'b0;
  assign \A[17][174] [3] = 1'b0;
  assign \A[17][174] [2] = 1'b0;
  assign \A[17][174] [1] = 1'b0;
  assign \A[17][176] [4] = 1'b0;
  assign \A[17][176] [3] = 1'b0;
  assign \A[17][176] [2] = 1'b0;
  assign \A[17][176] [1] = 1'b0;
  assign \A[17][176] [0] = 1'b0;
  assign \A[17][177] [1] = 1'b0;
  assign \A[17][178] [4] = 1'b0;
  assign \A[17][178] [3] = 1'b0;
  assign \A[17][178] [2] = 1'b0;
  assign \A[17][178] [1] = 1'b0;
  assign \A[17][179] [4] = 1'b0;
  assign \A[17][179] [3] = 1'b0;
  assign \A[17][179] [2] = 1'b0;
  assign \A[17][179] [1] = 1'b0;
  assign \A[17][179] [0] = 1'b0;
  assign \A[17][181] [4] = 1'b0;
  assign \A[17][181] [3] = 1'b0;
  assign \A[17][181] [2] = 1'b0;
  assign \A[17][181] [1] = 1'b0;
  assign \A[17][182] [4] = 1'b0;
  assign \A[17][182] [3] = 1'b0;
  assign \A[17][182] [2] = 1'b0;
  assign \A[17][183] [4] = 1'b0;
  assign \A[17][183] [3] = 1'b0;
  assign \A[17][183] [2] = 1'b0;
  assign \A[17][183] [1] = 1'b0;
  assign \A[17][184] [4] = 1'b0;
  assign \A[17][184] [3] = 1'b0;
  assign \A[17][184] [2] = 1'b0;
  assign \A[17][184] [1] = 1'b0;
  assign \A[17][184] [0] = 1'b0;
  assign \A[17][186] [1] = 1'b0;
  assign \A[17][188] [0] = 1'b0;
  assign \A[17][189] [4] = 1'b0;
  assign \A[17][189] [3] = 1'b0;
  assign \A[17][189] [2] = 1'b0;
  assign \A[17][189] [1] = 1'b0;
  assign \A[17][190] [4] = 1'b0;
  assign \A[17][190] [3] = 1'b0;
  assign \A[17][190] [2] = 1'b0;
  assign \A[17][190] [1] = 1'b0;
  assign \A[17][190] [0] = 1'b0;
  assign \A[17][191] [4] = 1'b0;
  assign \A[17][191] [3] = 1'b0;
  assign \A[17][191] [2] = 1'b0;
  assign \A[17][191] [0] = 1'b0;
  assign \A[17][192] [4] = 1'b0;
  assign \A[17][192] [3] = 1'b0;
  assign \A[17][192] [2] = 1'b0;
  assign \A[17][192] [1] = 1'b0;
  assign \A[17][193] [4] = 1'b0;
  assign \A[17][193] [3] = 1'b0;
  assign \A[17][193] [2] = 1'b0;
  assign \A[17][193] [1] = 1'b0;
  assign \A[17][193] [0] = 1'b0;
  assign \A[17][195] [4] = 1'b0;
  assign \A[17][195] [3] = 1'b0;
  assign \A[17][195] [2] = 1'b0;
  assign \A[17][195] [1] = 1'b0;
  assign \A[17][197] [4] = 1'b0;
  assign \A[17][197] [3] = 1'b0;
  assign \A[17][197] [2] = 1'b0;
  assign \A[17][197] [1] = 1'b0;
  assign \A[17][197] [0] = 1'b0;
  assign \A[17][198] [4] = 1'b0;
  assign \A[17][198] [3] = 1'b0;
  assign \A[17][198] [2] = 1'b0;
  assign \A[17][198] [1] = 1'b0;
  assign \A[17][198] [0] = 1'b0;
  assign \A[17][199] [1] = 1'b0;
  assign \A[17][200] [0] = 1'b0;
  assign \A[17][202] [4] = 1'b0;
  assign \A[17][202] [3] = 1'b0;
  assign \A[17][202] [2] = 1'b0;
  assign \A[17][202] [1] = 1'b0;
  assign \A[17][202] [0] = 1'b0;
  assign \A[17][203] [4] = 1'b0;
  assign \A[17][203] [3] = 1'b0;
  assign \A[17][203] [2] = 1'b0;
  assign \A[17][203] [0] = 1'b0;
  assign \A[17][204] [4] = 1'b0;
  assign \A[17][204] [3] = 1'b0;
  assign \A[17][204] [2] = 1'b0;
  assign \A[17][204] [0] = 1'b0;
  assign \A[17][205] [4] = 1'b0;
  assign \A[17][205] [3] = 1'b0;
  assign \A[17][205] [2] = 1'b0;
  assign \A[17][205] [1] = 1'b0;
  assign \A[17][205] [0] = 1'b0;
  assign \A[17][206] [4] = 1'b0;
  assign \A[17][206] [3] = 1'b0;
  assign \A[17][206] [2] = 1'b0;
  assign \A[17][206] [1] = 1'b0;
  assign \A[17][206] [0] = 1'b0;
  assign \A[17][207] [4] = 1'b0;
  assign \A[17][207] [3] = 1'b0;
  assign \A[17][207] [2] = 1'b0;
  assign \A[17][207] [1] = 1'b0;
  assign \A[17][208] [4] = 1'b0;
  assign \A[17][208] [3] = 1'b0;
  assign \A[17][208] [1] = 1'b0;
  assign \A[17][210] [4] = 1'b0;
  assign \A[17][210] [3] = 1'b0;
  assign \A[17][210] [2] = 1'b0;
  assign \A[17][210] [1] = 1'b0;
  assign \A[17][210] [0] = 1'b0;
  assign \A[17][212] [4] = 1'b0;
  assign \A[17][212] [3] = 1'b0;
  assign \A[17][212] [2] = 1'b0;
  assign \A[17][212] [0] = 1'b0;
  assign \A[17][213] [0] = 1'b0;
  assign \A[17][214] [4] = 1'b0;
  assign \A[17][214] [3] = 1'b0;
  assign \A[17][214] [2] = 1'b0;
  assign \A[17][214] [1] = 1'b0;
  assign \A[17][214] [0] = 1'b0;
  assign \A[17][216] [4] = 1'b0;
  assign \A[17][216] [3] = 1'b0;
  assign \A[17][216] [2] = 1'b0;
  assign \A[17][216] [1] = 1'b0;
  assign \A[17][216] [0] = 1'b0;
  assign \A[17][217] [4] = 1'b0;
  assign \A[17][217] [3] = 1'b0;
  assign \A[17][217] [2] = 1'b0;
  assign \A[17][217] [1] = 1'b0;
  assign \A[17][217] [0] = 1'b0;
  assign \A[17][218] [4] = 1'b0;
  assign \A[17][218] [3] = 1'b0;
  assign \A[17][218] [2] = 1'b0;
  assign \A[17][218] [1] = 1'b0;
  assign \A[17][218] [0] = 1'b0;
  assign \A[17][219] [4] = 1'b0;
  assign \A[17][219] [3] = 1'b0;
  assign \A[17][219] [2] = 1'b0;
  assign \A[17][220] [0] = 1'b0;
  assign \A[17][221] [4] = 1'b0;
  assign \A[17][221] [3] = 1'b0;
  assign \A[17][221] [2] = 1'b0;
  assign \A[17][221] [1] = 1'b0;
  assign \A[17][222] [4] = 1'b0;
  assign \A[17][222] [3] = 1'b0;
  assign \A[17][222] [1] = 1'b0;
  assign \A[17][224] [4] = 1'b0;
  assign \A[17][224] [3] = 1'b0;
  assign \A[17][224] [2] = 1'b0;
  assign \A[17][224] [1] = 1'b0;
  assign \A[17][225] [0] = 1'b0;
  assign \A[17][226] [4] = 1'b0;
  assign \A[17][226] [3] = 1'b0;
  assign \A[17][226] [2] = 1'b0;
  assign \A[17][226] [1] = 1'b0;
  assign \A[17][226] [0] = 1'b0;
  assign \A[17][227] [4] = 1'b0;
  assign \A[17][227] [3] = 1'b0;
  assign \A[17][227] [2] = 1'b0;
  assign \A[17][227] [1] = 1'b0;
  assign \A[17][227] [0] = 1'b0;
  assign \A[17][228] [4] = 1'b0;
  assign \A[17][228] [3] = 1'b0;
  assign \A[17][228] [2] = 1'b0;
  assign \A[17][228] [1] = 1'b0;
  assign \A[17][228] [0] = 1'b0;
  assign \A[17][229] [4] = 1'b0;
  assign \A[17][229] [3] = 1'b0;
  assign \A[17][229] [2] = 1'b0;
  assign \A[17][229] [0] = 1'b0;
  assign \A[17][230] [1] = 1'b0;
  assign \A[17][231] [4] = 1'b0;
  assign \A[17][231] [3] = 1'b0;
  assign \A[17][231] [2] = 1'b0;
  assign \A[17][231] [1] = 1'b0;
  assign \A[17][232] [4] = 1'b0;
  assign \A[17][232] [3] = 1'b0;
  assign \A[17][232] [2] = 1'b0;
  assign \A[17][232] [1] = 1'b0;
  assign \A[17][233] [4] = 1'b0;
  assign \A[17][233] [3] = 1'b0;
  assign \A[17][233] [2] = 1'b0;
  assign \A[17][233] [0] = 1'b0;
  assign \A[17][234] [4] = 1'b0;
  assign \A[17][234] [3] = 1'b0;
  assign \A[17][234] [2] = 1'b0;
  assign \A[17][234] [1] = 1'b0;
  assign \A[17][235] [4] = 1'b0;
  assign \A[17][235] [3] = 1'b0;
  assign \A[17][235] [2] = 1'b0;
  assign \A[17][235] [0] = 1'b0;
  assign \A[17][236] [4] = 1'b0;
  assign \A[17][236] [3] = 1'b0;
  assign \A[17][236] [2] = 1'b0;
  assign \A[17][236] [1] = 1'b0;
  assign \A[17][237] [4] = 1'b0;
  assign \A[17][237] [3] = 1'b0;
  assign \A[17][237] [1] = 1'b0;
  assign \A[17][237] [0] = 1'b0;
  assign \A[17][238] [0] = 1'b0;
  assign \A[17][239] [4] = 1'b0;
  assign \A[17][239] [3] = 1'b0;
  assign \A[17][239] [2] = 1'b0;
  assign \A[17][239] [1] = 1'b0;
  assign \A[17][240] [4] = 1'b0;
  assign \A[17][240] [3] = 1'b0;
  assign \A[17][240] [2] = 1'b0;
  assign \A[17][240] [0] = 1'b0;
  assign \A[17][241] [4] = 1'b0;
  assign \A[17][241] [3] = 1'b0;
  assign \A[17][241] [2] = 1'b0;
  assign \A[17][241] [1] = 1'b0;
  assign \A[17][242] [4] = 1'b0;
  assign \A[17][242] [3] = 1'b0;
  assign \A[17][242] [2] = 1'b0;
  assign \A[17][242] [1] = 1'b0;
  assign \A[17][242] [0] = 1'b0;
  assign \A[17][243] [4] = 1'b0;
  assign \A[17][243] [3] = 1'b0;
  assign \A[17][243] [2] = 1'b0;
  assign \A[17][243] [1] = 1'b0;
  assign \A[17][243] [0] = 1'b0;
  assign \A[17][244] [4] = 1'b0;
  assign \A[17][244] [3] = 1'b0;
  assign \A[17][244] [2] = 1'b0;
  assign \A[17][244] [1] = 1'b0;
  assign \A[17][244] [0] = 1'b0;
  assign \A[17][246] [0] = 1'b0;
  assign \A[17][247] [4] = 1'b0;
  assign \A[17][247] [3] = 1'b0;
  assign \A[17][247] [2] = 1'b0;
  assign \A[17][247] [1] = 1'b0;
  assign \A[17][247] [0] = 1'b0;
  assign \A[17][248] [0] = 1'b0;
  assign \A[17][249] [1] = 1'b0;
  assign \A[17][249] [0] = 1'b0;
  assign \A[17][250] [4] = 1'b0;
  assign \A[17][250] [3] = 1'b0;
  assign \A[17][250] [2] = 1'b0;
  assign \A[17][250] [0] = 1'b0;
  assign \A[17][251] [4] = 1'b0;
  assign \A[17][251] [3] = 1'b0;
  assign \A[17][251] [2] = 1'b0;
  assign \A[17][252] [4] = 1'b0;
  assign \A[17][252] [3] = 1'b0;
  assign \A[17][252] [2] = 1'b0;
  assign \A[17][252] [1] = 1'b0;
  assign \A[17][253] [4] = 1'b0;
  assign \A[17][253] [3] = 1'b0;
  assign \A[17][253] [2] = 1'b0;
  assign \A[17][253] [0] = 1'b0;
  assign \A[17][254] [4] = 1'b0;
  assign \A[17][254] [3] = 1'b0;
  assign \A[17][254] [2] = 1'b0;
  assign \A[17][254] [1] = 1'b0;
  assign \A[18][0] [4] = 1'b0;
  assign \A[18][0] [3] = 1'b0;
  assign \A[18][0] [2] = 1'b0;
  assign \A[18][0] [1] = 1'b0;
  assign \A[18][1] [4] = 1'b0;
  assign \A[18][1] [3] = 1'b0;
  assign \A[18][1] [2] = 1'b0;
  assign \A[18][2] [4] = 1'b0;
  assign \A[18][2] [3] = 1'b0;
  assign \A[18][2] [2] = 1'b0;
  assign \A[18][2] [1] = 1'b0;
  assign \A[18][3] [4] = 1'b0;
  assign \A[18][3] [3] = 1'b0;
  assign \A[18][3] [2] = 1'b0;
  assign \A[18][3] [1] = 1'b0;
  assign \A[18][4] [4] = 1'b0;
  assign \A[18][4] [3] = 1'b0;
  assign \A[18][4] [2] = 1'b0;
  assign \A[18][4] [1] = 1'b0;
  assign \A[18][4] [0] = 1'b0;
  assign \A[18][5] [4] = 1'b0;
  assign \A[18][5] [3] = 1'b0;
  assign \A[18][5] [2] = 1'b0;
  assign \A[18][5] [1] = 1'b0;
  assign \A[18][5] [0] = 1'b0;
  assign \A[18][6] [4] = 1'b0;
  assign \A[18][6] [3] = 1'b0;
  assign \A[18][6] [2] = 1'b0;
  assign \A[18][6] [1] = 1'b0;
  assign \A[18][6] [0] = 1'b0;
  assign \A[18][8] [4] = 1'b0;
  assign \A[18][8] [3] = 1'b0;
  assign \A[18][8] [2] = 1'b0;
  assign \A[18][8] [1] = 1'b0;
  assign \A[18][8] [0] = 1'b0;
  assign \A[18][9] [4] = 1'b0;
  assign \A[18][9] [3] = 1'b0;
  assign \A[18][9] [2] = 1'b0;
  assign \A[18][9] [1] = 1'b0;
  assign \A[18][10] [4] = 1'b0;
  assign \A[18][10] [3] = 1'b0;
  assign \A[18][10] [2] = 1'b0;
  assign \A[18][10] [0] = 1'b0;
  assign \A[18][11] [4] = 1'b0;
  assign \A[18][11] [3] = 1'b0;
  assign \A[18][11] [2] = 1'b0;
  assign \A[18][11] [1] = 1'b0;
  assign \A[18][11] [0] = 1'b0;
  assign \A[18][12] [4] = 1'b0;
  assign \A[18][12] [3] = 1'b0;
  assign \A[18][12] [2] = 1'b0;
  assign \A[18][12] [0] = 1'b0;
  assign \A[18][14] [0] = 1'b0;
  assign \A[18][15] [4] = 1'b0;
  assign \A[18][15] [3] = 1'b0;
  assign \A[18][15] [2] = 1'b0;
  assign \A[18][15] [1] = 1'b0;
  assign \A[18][16] [1] = 1'b0;
  assign \A[18][17] [4] = 1'b0;
  assign \A[18][17] [3] = 1'b0;
  assign \A[18][17] [2] = 1'b0;
  assign \A[18][17] [0] = 1'b0;
  assign \A[18][19] [4] = 1'b0;
  assign \A[18][19] [3] = 1'b0;
  assign \A[18][19] [2] = 1'b0;
  assign \A[18][19] [0] = 1'b0;
  assign \A[18][20] [4] = 1'b0;
  assign \A[18][20] [3] = 1'b0;
  assign \A[18][20] [2] = 1'b0;
  assign \A[18][20] [1] = 1'b0;
  assign \A[18][20] [0] = 1'b0;
  assign \A[18][21] [4] = 1'b0;
  assign \A[18][21] [3] = 1'b0;
  assign \A[18][21] [2] = 1'b0;
  assign \A[18][21] [1] = 1'b0;
  assign \A[18][23] [4] = 1'b0;
  assign \A[18][23] [3] = 1'b0;
  assign \A[18][23] [2] = 1'b0;
  assign \A[18][23] [1] = 1'b0;
  assign \A[18][23] [0] = 1'b0;
  assign \A[18][24] [4] = 1'b0;
  assign \A[18][24] [3] = 1'b0;
  assign \A[18][24] [2] = 1'b0;
  assign \A[18][24] [0] = 1'b0;
  assign \A[18][25] [4] = 1'b0;
  assign \A[18][25] [3] = 1'b0;
  assign \A[18][25] [2] = 1'b0;
  assign \A[18][26] [4] = 1'b0;
  assign \A[18][26] [3] = 1'b0;
  assign \A[18][26] [2] = 1'b0;
  assign \A[18][26] [1] = 1'b0;
  assign \A[18][26] [0] = 1'b0;
  assign \A[18][27] [4] = 1'b0;
  assign \A[18][27] [3] = 1'b0;
  assign \A[18][27] [2] = 1'b0;
  assign \A[18][27] [1] = 1'b0;
  assign \A[18][27] [0] = 1'b0;
  assign \A[18][29] [4] = 1'b0;
  assign \A[18][29] [3] = 1'b0;
  assign \A[18][29] [2] = 1'b0;
  assign \A[18][29] [1] = 1'b0;
  assign \A[18][29] [0] = 1'b0;
  assign \A[18][30] [4] = 1'b0;
  assign \A[18][30] [3] = 1'b0;
  assign \A[18][30] [1] = 1'b0;
  assign \A[18][30] [0] = 1'b0;
  assign \A[18][31] [0] = 1'b0;
  assign \A[18][33] [1] = 1'b0;
  assign \A[18][36] [0] = 1'b0;
  assign \A[18][37] [1] = 1'b0;
  assign \A[18][38] [4] = 1'b0;
  assign \A[18][38] [3] = 1'b0;
  assign \A[18][38] [2] = 1'b0;
  assign \A[18][38] [1] = 1'b0;
  assign \A[18][38] [0] = 1'b0;
  assign \A[18][39] [4] = 1'b0;
  assign \A[18][39] [3] = 1'b0;
  assign \A[18][39] [2] = 1'b0;
  assign \A[18][39] [1] = 1'b0;
  assign \A[18][39] [0] = 1'b0;
  assign \A[18][41] [0] = 1'b0;
  assign \A[18][42] [4] = 1'b0;
  assign \A[18][42] [3] = 1'b0;
  assign \A[18][42] [2] = 1'b0;
  assign \A[18][42] [0] = 1'b0;
  assign \A[18][43] [4] = 1'b0;
  assign \A[18][43] [3] = 1'b0;
  assign \A[18][43] [2] = 1'b0;
  assign \A[18][43] [0] = 1'b0;
  assign \A[18][44] [4] = 1'b0;
  assign \A[18][44] [3] = 1'b0;
  assign \A[18][44] [2] = 1'b0;
  assign \A[18][44] [1] = 1'b0;
  assign \A[18][45] [4] = 1'b0;
  assign \A[18][45] [3] = 1'b0;
  assign \A[18][45] [2] = 1'b0;
  assign \A[18][45] [1] = 1'b0;
  assign \A[18][46] [4] = 1'b0;
  assign \A[18][46] [3] = 1'b0;
  assign \A[18][46] [2] = 1'b0;
  assign \A[18][46] [1] = 1'b0;
  assign \A[18][46] [0] = 1'b0;
  assign \A[18][47] [4] = 1'b0;
  assign \A[18][47] [3] = 1'b0;
  assign \A[18][47] [1] = 1'b0;
  assign \A[18][47] [0] = 1'b0;
  assign \A[18][48] [4] = 1'b0;
  assign \A[18][48] [3] = 1'b0;
  assign \A[18][48] [2] = 1'b0;
  assign \A[18][49] [4] = 1'b0;
  assign \A[18][49] [3] = 1'b0;
  assign \A[18][49] [2] = 1'b0;
  assign \A[18][49] [1] = 1'b0;
  assign \A[18][49] [0] = 1'b0;
  assign \A[18][50] [0] = 1'b0;
  assign \A[18][51] [4] = 1'b0;
  assign \A[18][51] [3] = 1'b0;
  assign \A[18][51] [2] = 1'b0;
  assign \A[18][51] [1] = 1'b0;
  assign \A[18][53] [4] = 1'b0;
  assign \A[18][53] [3] = 1'b0;
  assign \A[18][53] [2] = 1'b0;
  assign \A[18][53] [1] = 1'b0;
  assign \A[18][53] [0] = 1'b0;
  assign \A[18][54] [0] = 1'b0;
  assign \A[18][56] [4] = 1'b0;
  assign \A[18][56] [3] = 1'b0;
  assign \A[18][56] [2] = 1'b0;
  assign \A[18][56] [1] = 1'b0;
  assign \A[18][57] [4] = 1'b0;
  assign \A[18][57] [3] = 1'b0;
  assign \A[18][57] [2] = 1'b0;
  assign \A[18][57] [1] = 1'b0;
  assign \A[18][58] [4] = 1'b0;
  assign \A[18][58] [3] = 1'b0;
  assign \A[18][58] [1] = 1'b0;
  assign \A[18][58] [0] = 1'b0;
  assign \A[18][59] [4] = 1'b0;
  assign \A[18][59] [3] = 1'b0;
  assign \A[18][59] [2] = 1'b0;
  assign \A[18][59] [1] = 1'b0;
  assign \A[18][59] [0] = 1'b0;
  assign \A[18][60] [4] = 1'b0;
  assign \A[18][60] [3] = 1'b0;
  assign \A[18][60] [2] = 1'b0;
  assign \A[18][60] [1] = 1'b0;
  assign \A[18][61] [4] = 1'b0;
  assign \A[18][61] [3] = 1'b0;
  assign \A[18][61] [2] = 1'b0;
  assign \A[18][61] [1] = 1'b0;
  assign \A[18][62] [4] = 1'b0;
  assign \A[18][62] [3] = 1'b0;
  assign \A[18][62] [2] = 1'b0;
  assign \A[18][62] [1] = 1'b0;
  assign \A[18][63] [4] = 1'b0;
  assign \A[18][63] [3] = 1'b0;
  assign \A[18][63] [2] = 1'b0;
  assign \A[18][63] [1] = 1'b0;
  assign \A[18][64] [0] = 1'b0;
  assign \A[18][66] [1] = 1'b0;
  assign \A[18][66] [0] = 1'b0;
  assign \A[18][67] [4] = 1'b0;
  assign \A[18][67] [3] = 1'b0;
  assign \A[18][67] [2] = 1'b0;
  assign \A[18][67] [1] = 1'b0;
  assign \A[18][67] [0] = 1'b0;
  assign \A[18][68] [4] = 1'b0;
  assign \A[18][68] [3] = 1'b0;
  assign \A[18][68] [2] = 1'b0;
  assign \A[18][68] [1] = 1'b0;
  assign \A[18][69] [4] = 1'b0;
  assign \A[18][69] [3] = 1'b0;
  assign \A[18][69] [2] = 1'b0;
  assign \A[18][69] [1] = 1'b0;
  assign \A[18][70] [4] = 1'b0;
  assign \A[18][70] [3] = 1'b0;
  assign \A[18][70] [2] = 1'b0;
  assign \A[18][70] [1] = 1'b0;
  assign \A[18][70] [0] = 1'b0;
  assign \A[18][73] [0] = 1'b0;
  assign \A[18][74] [4] = 1'b0;
  assign \A[18][74] [3] = 1'b0;
  assign \A[18][74] [2] = 1'b0;
  assign \A[18][74] [1] = 1'b0;
  assign \A[18][74] [0] = 1'b0;
  assign \A[18][76] [4] = 1'b0;
  assign \A[18][76] [3] = 1'b0;
  assign \A[18][76] [2] = 1'b0;
  assign \A[18][76] [1] = 1'b0;
  assign \A[18][78] [4] = 1'b0;
  assign \A[18][78] [3] = 1'b0;
  assign \A[18][78] [2] = 1'b0;
  assign \A[18][78] [0] = 1'b0;
  assign \A[18][80] [4] = 1'b0;
  assign \A[18][80] [3] = 1'b0;
  assign \A[18][80] [2] = 1'b0;
  assign \A[18][80] [1] = 1'b0;
  assign \A[18][81] [4] = 1'b0;
  assign \A[18][81] [3] = 1'b0;
  assign \A[18][81] [2] = 1'b0;
  assign \A[18][81] [1] = 1'b0;
  assign \A[18][82] [4] = 1'b0;
  assign \A[18][82] [3] = 1'b0;
  assign \A[18][82] [2] = 1'b0;
  assign \A[18][82] [1] = 1'b0;
  assign \A[18][82] [0] = 1'b0;
  assign \A[18][85] [4] = 1'b0;
  assign \A[18][85] [3] = 1'b0;
  assign \A[18][85] [2] = 1'b0;
  assign \A[18][85] [1] = 1'b0;
  assign \A[18][85] [0] = 1'b0;
  assign \A[18][86] [4] = 1'b0;
  assign \A[18][86] [3] = 1'b0;
  assign \A[18][86] [2] = 1'b0;
  assign \A[18][86] [1] = 1'b0;
  assign \A[18][87] [4] = 1'b0;
  assign \A[18][87] [3] = 1'b0;
  assign \A[18][87] [2] = 1'b0;
  assign \A[18][87] [1] = 1'b0;
  assign \A[18][87] [0] = 1'b0;
  assign \A[18][88] [0] = 1'b0;
  assign \A[18][89] [1] = 1'b0;
  assign \A[18][89] [0] = 1'b0;
  assign \A[18][91] [1] = 1'b0;
  assign \A[18][92] [0] = 1'b0;
  assign \A[18][93] [0] = 1'b0;
  assign \A[18][94] [4] = 1'b0;
  assign \A[18][94] [3] = 1'b0;
  assign \A[18][94] [2] = 1'b0;
  assign \A[18][94] [1] = 1'b0;
  assign \A[18][94] [0] = 1'b0;
  assign \A[18][95] [4] = 1'b0;
  assign \A[18][95] [3] = 1'b0;
  assign \A[18][95] [2] = 1'b0;
  assign \A[18][97] [4] = 1'b0;
  assign \A[18][97] [3] = 1'b0;
  assign \A[18][97] [2] = 1'b0;
  assign \A[18][97] [1] = 1'b0;
  assign \A[18][99] [0] = 1'b0;
  assign \A[18][101] [4] = 1'b0;
  assign \A[18][101] [3] = 1'b0;
  assign \A[18][101] [2] = 1'b0;
  assign \A[18][101] [1] = 1'b0;
  assign \A[18][101] [0] = 1'b0;
  assign \A[18][102] [4] = 1'b0;
  assign \A[18][102] [3] = 1'b0;
  assign \A[18][102] [2] = 1'b0;
  assign \A[18][102] [1] = 1'b0;
  assign \A[18][102] [0] = 1'b0;
  assign \A[18][103] [1] = 1'b0;
  assign \A[18][104] [0] = 1'b0;
  assign \A[18][105] [0] = 1'b0;
  assign \A[18][106] [4] = 1'b0;
  assign \A[18][106] [3] = 1'b0;
  assign \A[18][106] [2] = 1'b0;
  assign \A[18][106] [1] = 1'b0;
  assign \A[18][107] [4] = 1'b0;
  assign \A[18][107] [3] = 1'b0;
  assign \A[18][107] [2] = 1'b0;
  assign \A[18][107] [1] = 1'b0;
  assign \A[18][107] [0] = 1'b0;
  assign \A[18][109] [4] = 1'b0;
  assign \A[18][109] [3] = 1'b0;
  assign \A[18][109] [2] = 1'b0;
  assign \A[18][109] [1] = 1'b0;
  assign \A[18][109] [0] = 1'b0;
  assign \A[18][110] [4] = 1'b0;
  assign \A[18][110] [3] = 1'b0;
  assign \A[18][110] [2] = 1'b0;
  assign \A[18][111] [4] = 1'b0;
  assign \A[18][111] [3] = 1'b0;
  assign \A[18][111] [2] = 1'b0;
  assign \A[18][111] [1] = 1'b0;
  assign \A[18][112] [4] = 1'b0;
  assign \A[18][112] [3] = 1'b0;
  assign \A[18][112] [2] = 1'b0;
  assign \A[18][113] [4] = 1'b0;
  assign \A[18][113] [3] = 1'b0;
  assign \A[18][113] [2] = 1'b0;
  assign \A[18][113] [1] = 1'b0;
  assign \A[18][114] [0] = 1'b0;
  assign \A[18][115] [4] = 1'b0;
  assign \A[18][115] [3] = 1'b0;
  assign \A[18][115] [2] = 1'b0;
  assign \A[18][115] [1] = 1'b0;
  assign \A[18][115] [0] = 1'b0;
  assign \A[18][116] [4] = 1'b0;
  assign \A[18][116] [3] = 1'b0;
  assign \A[18][116] [2] = 1'b0;
  assign \A[18][116] [1] = 1'b0;
  assign \A[18][117] [0] = 1'b0;
  assign \A[18][119] [4] = 1'b0;
  assign \A[18][119] [3] = 1'b0;
  assign \A[18][119] [2] = 1'b0;
  assign \A[18][119] [1] = 1'b0;
  assign \A[18][119] [0] = 1'b0;
  assign \A[18][120] [4] = 1'b0;
  assign \A[18][120] [3] = 1'b0;
  assign \A[18][120] [2] = 1'b0;
  assign \A[18][120] [1] = 1'b0;
  assign \A[18][120] [0] = 1'b0;
  assign \A[18][121] [4] = 1'b0;
  assign \A[18][121] [3] = 1'b0;
  assign \A[18][121] [2] = 1'b0;
  assign \A[18][121] [1] = 1'b0;
  assign \A[18][121] [0] = 1'b0;
  assign \A[18][122] [1] = 1'b0;
  assign \A[18][123] [0] = 1'b0;
  assign \A[18][124] [0] = 1'b0;
  assign \A[18][125] [4] = 1'b0;
  assign \A[18][125] [3] = 1'b0;
  assign \A[18][125] [2] = 1'b0;
  assign \A[18][125] [0] = 1'b0;
  assign \A[18][126] [4] = 1'b0;
  assign \A[18][126] [3] = 1'b0;
  assign \A[18][126] [1] = 1'b0;
  assign \A[18][129] [4] = 1'b0;
  assign \A[18][129] [3] = 1'b0;
  assign \A[18][129] [2] = 1'b0;
  assign \A[18][130] [4] = 1'b0;
  assign \A[18][130] [3] = 1'b0;
  assign \A[18][130] [2] = 1'b0;
  assign \A[18][130] [1] = 1'b0;
  assign \A[18][131] [1] = 1'b0;
  assign \A[18][132] [1] = 1'b0;
  assign \A[18][136] [4] = 1'b0;
  assign \A[18][136] [3] = 1'b0;
  assign \A[18][136] [2] = 1'b0;
  assign \A[18][136] [1] = 1'b0;
  assign \A[18][140] [4] = 1'b0;
  assign \A[18][140] [3] = 1'b0;
  assign \A[18][140] [2] = 1'b0;
  assign \A[18][140] [1] = 1'b0;
  assign \A[18][140] [0] = 1'b0;
  assign \A[18][142] [4] = 1'b0;
  assign \A[18][142] [3] = 1'b0;
  assign \A[18][142] [2] = 1'b0;
  assign \A[18][142] [1] = 1'b0;
  assign \A[18][143] [4] = 1'b0;
  assign \A[18][143] [3] = 1'b0;
  assign \A[18][143] [2] = 1'b0;
  assign \A[18][143] [1] = 1'b0;
  assign \A[18][144] [4] = 1'b0;
  assign \A[18][144] [3] = 1'b0;
  assign \A[18][144] [2] = 1'b0;
  assign \A[18][144] [1] = 1'b0;
  assign \A[18][145] [4] = 1'b0;
  assign \A[18][145] [3] = 1'b0;
  assign \A[18][145] [2] = 1'b0;
  assign \A[18][145] [1] = 1'b0;
  assign \A[18][147] [4] = 1'b0;
  assign \A[18][147] [3] = 1'b0;
  assign \A[18][147] [2] = 1'b0;
  assign \A[18][147] [1] = 1'b0;
  assign \A[18][147] [0] = 1'b0;
  assign \A[18][148] [4] = 1'b0;
  assign \A[18][148] [3] = 1'b0;
  assign \A[18][148] [2] = 1'b0;
  assign \A[18][148] [1] = 1'b0;
  assign \A[18][150] [4] = 1'b0;
  assign \A[18][150] [3] = 1'b0;
  assign \A[18][150] [2] = 1'b0;
  assign \A[18][150] [1] = 1'b0;
  assign \A[18][150] [0] = 1'b0;
  assign \A[18][151] [1] = 1'b0;
  assign \A[18][152] [0] = 1'b0;
  assign \A[18][153] [4] = 1'b0;
  assign \A[18][153] [3] = 1'b0;
  assign \A[18][153] [2] = 1'b0;
  assign \A[18][154] [4] = 1'b0;
  assign \A[18][154] [3] = 1'b0;
  assign \A[18][154] [2] = 1'b0;
  assign \A[18][154] [1] = 1'b0;
  assign \A[18][154] [0] = 1'b0;
  assign \A[18][155] [4] = 1'b0;
  assign \A[18][155] [3] = 1'b0;
  assign \A[18][155] [2] = 1'b0;
  assign \A[18][155] [0] = 1'b0;
  assign \A[18][157] [4] = 1'b0;
  assign \A[18][157] [3] = 1'b0;
  assign \A[18][157] [2] = 1'b0;
  assign \A[18][157] [1] = 1'b0;
  assign \A[18][158] [4] = 1'b0;
  assign \A[18][158] [3] = 1'b0;
  assign \A[18][158] [2] = 1'b0;
  assign \A[18][158] [1] = 1'b0;
  assign \A[18][159] [4] = 1'b0;
  assign \A[18][159] [3] = 1'b0;
  assign \A[18][159] [1] = 1'b0;
  assign \A[18][159] [0] = 1'b0;
  assign \A[18][160] [4] = 1'b0;
  assign \A[18][160] [3] = 1'b0;
  assign \A[18][160] [2] = 1'b0;
  assign \A[18][160] [0] = 1'b0;
  assign \A[18][161] [4] = 1'b0;
  assign \A[18][161] [3] = 1'b0;
  assign \A[18][161] [2] = 1'b0;
  assign \A[18][161] [1] = 1'b0;
  assign \A[18][161] [0] = 1'b0;
  assign \A[18][162] [4] = 1'b0;
  assign \A[18][162] [3] = 1'b0;
  assign \A[18][162] [2] = 1'b0;
  assign \A[18][162] [0] = 1'b0;
  assign \A[18][163] [0] = 1'b0;
  assign \A[18][164] [4] = 1'b0;
  assign \A[18][164] [3] = 1'b0;
  assign \A[18][164] [2] = 1'b0;
  assign \A[18][164] [1] = 1'b0;
  assign \A[18][164] [0] = 1'b0;
  assign \A[18][165] [1] = 1'b0;
  assign \A[18][167] [1] = 1'b0;
  assign \A[18][168] [4] = 1'b0;
  assign \A[18][168] [3] = 1'b0;
  assign \A[18][168] [2] = 1'b0;
  assign \A[18][168] [1] = 1'b0;
  assign \A[18][168] [0] = 1'b0;
  assign \A[18][169] [4] = 1'b0;
  assign \A[18][169] [3] = 1'b0;
  assign \A[18][169] [2] = 1'b0;
  assign \A[18][169] [1] = 1'b0;
  assign \A[18][169] [0] = 1'b0;
  assign \A[18][170] [4] = 1'b0;
  assign \A[18][170] [3] = 1'b0;
  assign \A[18][170] [2] = 1'b0;
  assign \A[18][170] [1] = 1'b0;
  assign \A[18][170] [0] = 1'b0;
  assign \A[18][171] [1] = 1'b0;
  assign \A[18][174] [4] = 1'b0;
  assign \A[18][174] [3] = 1'b0;
  assign \A[18][174] [2] = 1'b0;
  assign \A[18][174] [1] = 1'b0;
  assign \A[18][174] [0] = 1'b0;
  assign \A[18][175] [4] = 1'b0;
  assign \A[18][175] [3] = 1'b0;
  assign \A[18][175] [2] = 1'b0;
  assign \A[18][175] [1] = 1'b0;
  assign \A[18][177] [1] = 1'b0;
  assign \A[18][178] [4] = 1'b0;
  assign \A[18][178] [3] = 1'b0;
  assign \A[18][178] [2] = 1'b0;
  assign \A[18][178] [1] = 1'b0;
  assign \A[18][178] [0] = 1'b0;
  assign \A[18][179] [4] = 1'b0;
  assign \A[18][179] [3] = 1'b0;
  assign \A[18][179] [2] = 1'b0;
  assign \A[18][179] [1] = 1'b0;
  assign \A[18][180] [4] = 1'b0;
  assign \A[18][180] [3] = 1'b0;
  assign \A[18][180] [2] = 1'b0;
  assign \A[18][181] [4] = 1'b0;
  assign \A[18][181] [3] = 1'b0;
  assign \A[18][181] [2] = 1'b0;
  assign \A[18][181] [0] = 1'b0;
  assign \A[18][182] [4] = 1'b0;
  assign \A[18][182] [3] = 1'b0;
  assign \A[18][182] [2] = 1'b0;
  assign \A[18][182] [1] = 1'b0;
  assign \A[18][182] [0] = 1'b0;
  assign \A[18][183] [0] = 1'b0;
  assign \A[18][184] [4] = 1'b0;
  assign \A[18][184] [3] = 1'b0;
  assign \A[18][184] [2] = 1'b0;
  assign \A[18][184] [1] = 1'b0;
  assign \A[18][184] [0] = 1'b0;
  assign \A[18][185] [4] = 1'b0;
  assign \A[18][185] [3] = 1'b0;
  assign \A[18][185] [2] = 1'b0;
  assign \A[18][185] [0] = 1'b0;
  assign \A[18][186] [4] = 1'b0;
  assign \A[18][186] [3] = 1'b0;
  assign \A[18][186] [2] = 1'b0;
  assign \A[18][187] [4] = 1'b0;
  assign \A[18][187] [3] = 1'b0;
  assign \A[18][187] [2] = 1'b0;
  assign \A[18][187] [1] = 1'b0;
  assign \A[18][187] [0] = 1'b0;
  assign \A[18][190] [4] = 1'b0;
  assign \A[18][190] [3] = 1'b0;
  assign \A[18][190] [2] = 1'b0;
  assign \A[18][190] [1] = 1'b0;
  assign \A[18][192] [4] = 1'b0;
  assign \A[18][192] [3] = 1'b0;
  assign \A[18][192] [2] = 1'b0;
  assign \A[18][193] [4] = 1'b0;
  assign \A[18][193] [3] = 1'b0;
  assign \A[18][193] [2] = 1'b0;
  assign \A[18][193] [1] = 1'b0;
  assign \A[18][193] [0] = 1'b0;
  assign \A[18][195] [4] = 1'b0;
  assign \A[18][195] [3] = 1'b0;
  assign \A[18][195] [2] = 1'b0;
  assign \A[18][195] [1] = 1'b0;
  assign \A[18][195] [0] = 1'b0;
  assign \A[18][196] [4] = 1'b0;
  assign \A[18][196] [3] = 1'b0;
  assign \A[18][196] [2] = 1'b0;
  assign \A[18][196] [1] = 1'b0;
  assign \A[18][196] [0] = 1'b0;
  assign \A[18][197] [4] = 1'b0;
  assign \A[18][197] [3] = 1'b0;
  assign \A[18][197] [2] = 1'b0;
  assign \A[18][197] [1] = 1'b0;
  assign \A[18][198] [4] = 1'b0;
  assign \A[18][198] [3] = 1'b0;
  assign \A[18][198] [2] = 1'b0;
  assign \A[18][198] [1] = 1'b0;
  assign \A[18][199] [4] = 1'b0;
  assign \A[18][199] [3] = 1'b0;
  assign \A[18][199] [2] = 1'b0;
  assign \A[18][199] [1] = 1'b0;
  assign \A[18][200] [4] = 1'b0;
  assign \A[18][200] [3] = 1'b0;
  assign \A[18][200] [2] = 1'b0;
  assign \A[18][200] [1] = 1'b0;
  assign \A[18][200] [0] = 1'b0;
  assign \A[18][201] [4] = 1'b0;
  assign \A[18][201] [3] = 1'b0;
  assign \A[18][201] [2] = 1'b0;
  assign \A[18][201] [1] = 1'b0;
  assign \A[18][202] [4] = 1'b0;
  assign \A[18][202] [3] = 1'b0;
  assign \A[18][202] [2] = 1'b0;
  assign \A[18][202] [1] = 1'b0;
  assign \A[18][203] [4] = 1'b0;
  assign \A[18][203] [3] = 1'b0;
  assign \A[18][203] [2] = 1'b0;
  assign \A[18][203] [0] = 1'b0;
  assign \A[18][204] [4] = 1'b0;
  assign \A[18][204] [3] = 1'b0;
  assign \A[18][204] [2] = 1'b0;
  assign \A[18][204] [0] = 1'b0;
  assign \A[18][205] [4] = 1'b0;
  assign \A[18][205] [3] = 1'b0;
  assign \A[18][205] [2] = 1'b0;
  assign \A[18][205] [1] = 1'b0;
  assign \A[18][208] [4] = 1'b0;
  assign \A[18][208] [3] = 1'b0;
  assign \A[18][208] [2] = 1'b0;
  assign \A[18][208] [1] = 1'b0;
  assign \A[18][209] [4] = 1'b0;
  assign \A[18][209] [3] = 1'b0;
  assign \A[18][209] [2] = 1'b0;
  assign \A[18][210] [4] = 1'b0;
  assign \A[18][210] [3] = 1'b0;
  assign \A[18][210] [2] = 1'b0;
  assign \A[18][210] [1] = 1'b0;
  assign \A[18][211] [4] = 1'b0;
  assign \A[18][211] [3] = 1'b0;
  assign \A[18][211] [2] = 1'b0;
  assign \A[18][211] [0] = 1'b0;
  assign \A[18][212] [4] = 1'b0;
  assign \A[18][212] [3] = 1'b0;
  assign \A[18][212] [2] = 1'b0;
  assign \A[18][213] [4] = 1'b0;
  assign \A[18][213] [3] = 1'b0;
  assign \A[18][213] [2] = 1'b0;
  assign \A[18][213] [1] = 1'b0;
  assign \A[18][213] [0] = 1'b0;
  assign \A[18][215] [4] = 1'b0;
  assign \A[18][215] [3] = 1'b0;
  assign \A[18][215] [2] = 1'b0;
  assign \A[18][216] [4] = 1'b0;
  assign \A[18][216] [3] = 1'b0;
  assign \A[18][216] [2] = 1'b0;
  assign \A[18][216] [1] = 1'b0;
  assign \A[18][216] [0] = 1'b0;
  assign \A[18][218] [4] = 1'b0;
  assign \A[18][218] [3] = 1'b0;
  assign \A[18][218] [2] = 1'b0;
  assign \A[18][218] [1] = 1'b0;
  assign \A[18][218] [0] = 1'b0;
  assign \A[18][219] [0] = 1'b0;
  assign \A[18][220] [4] = 1'b0;
  assign \A[18][220] [3] = 1'b0;
  assign \A[18][220] [2] = 1'b0;
  assign \A[18][220] [1] = 1'b0;
  assign \A[18][220] [0] = 1'b0;
  assign \A[18][222] [4] = 1'b0;
  assign \A[18][222] [3] = 1'b0;
  assign \A[18][222] [2] = 1'b0;
  assign \A[18][222] [1] = 1'b0;
  assign \A[18][222] [0] = 1'b0;
  assign \A[18][223] [0] = 1'b0;
  assign \A[18][224] [4] = 1'b0;
  assign \A[18][224] [3] = 1'b0;
  assign \A[18][224] [2] = 1'b0;
  assign \A[18][224] [0] = 1'b0;
  assign \A[18][225] [4] = 1'b0;
  assign \A[18][225] [3] = 1'b0;
  assign \A[18][225] [2] = 1'b0;
  assign \A[18][225] [0] = 1'b0;
  assign \A[18][226] [4] = 1'b0;
  assign \A[18][226] [3] = 1'b0;
  assign \A[18][226] [2] = 1'b0;
  assign \A[18][226] [1] = 1'b0;
  assign \A[18][227] [4] = 1'b0;
  assign \A[18][227] [3] = 1'b0;
  assign \A[18][227] [2] = 1'b0;
  assign \A[18][227] [1] = 1'b0;
  assign \A[18][227] [0] = 1'b0;
  assign \A[18][229] [4] = 1'b0;
  assign \A[18][229] [3] = 1'b0;
  assign \A[18][229] [2] = 1'b0;
  assign \A[18][229] [0] = 1'b0;
  assign \A[18][231] [4] = 1'b0;
  assign \A[18][231] [3] = 1'b0;
  assign \A[18][231] [2] = 1'b0;
  assign \A[18][232] [4] = 1'b0;
  assign \A[18][232] [3] = 1'b0;
  assign \A[18][232] [2] = 1'b0;
  assign \A[18][232] [1] = 1'b0;
  assign \A[18][232] [0] = 1'b0;
  assign \A[18][233] [4] = 1'b0;
  assign \A[18][233] [3] = 1'b0;
  assign \A[18][233] [2] = 1'b0;
  assign \A[18][233] [0] = 1'b0;
  assign \A[18][234] [4] = 1'b0;
  assign \A[18][234] [3] = 1'b0;
  assign \A[18][234] [2] = 1'b0;
  assign \A[18][234] [1] = 1'b0;
  assign \A[18][234] [0] = 1'b0;
  assign \A[18][235] [0] = 1'b0;
  assign \A[18][236] [4] = 1'b0;
  assign \A[18][236] [3] = 1'b0;
  assign \A[18][236] [2] = 1'b0;
  assign \A[18][236] [1] = 1'b0;
  assign \A[18][236] [0] = 1'b0;
  assign \A[18][237] [0] = 1'b0;
  assign \A[18][240] [4] = 1'b0;
  assign \A[18][240] [3] = 1'b0;
  assign \A[18][240] [2] = 1'b0;
  assign \A[18][240] [1] = 1'b0;
  assign \A[18][241] [4] = 1'b0;
  assign \A[18][241] [3] = 1'b0;
  assign \A[18][241] [2] = 1'b0;
  assign \A[18][241] [0] = 1'b0;
  assign \A[18][242] [4] = 1'b0;
  assign \A[18][242] [3] = 1'b0;
  assign \A[18][242] [2] = 1'b0;
  assign \A[18][242] [1] = 1'b0;
  assign \A[18][243] [4] = 1'b0;
  assign \A[18][243] [3] = 1'b0;
  assign \A[18][243] [2] = 1'b0;
  assign \A[18][243] [1] = 1'b0;
  assign \A[18][243] [0] = 1'b0;
  assign \A[18][244] [0] = 1'b0;
  assign \A[18][246] [4] = 1'b0;
  assign \A[18][246] [3] = 1'b0;
  assign \A[18][246] [2] = 1'b0;
  assign \A[18][247] [4] = 1'b0;
  assign \A[18][247] [3] = 1'b0;
  assign \A[18][247] [2] = 1'b0;
  assign \A[18][247] [0] = 1'b0;
  assign \A[18][248] [4] = 1'b0;
  assign \A[18][248] [3] = 1'b0;
  assign \A[18][248] [2] = 1'b0;
  assign \A[18][248] [1] = 1'b0;
  assign \A[18][248] [0] = 1'b0;
  assign \A[18][249] [4] = 1'b0;
  assign \A[18][249] [3] = 1'b0;
  assign \A[18][249] [2] = 1'b0;
  assign \A[18][249] [1] = 1'b0;
  assign \A[18][249] [0] = 1'b0;
  assign \A[18][251] [4] = 1'b0;
  assign \A[18][251] [3] = 1'b0;
  assign \A[18][251] [2] = 1'b0;
  assign \A[18][251] [1] = 1'b0;
  assign \A[18][252] [4] = 1'b0;
  assign \A[18][252] [3] = 1'b0;
  assign \A[18][252] [2] = 1'b0;
  assign \A[18][252] [1] = 1'b0;
  assign \A[18][252] [0] = 1'b0;
  assign \A[18][255] [4] = 1'b0;
  assign \A[18][255] [3] = 1'b0;
  assign \A[18][255] [2] = 1'b0;
  assign \A[18][255] [1] = 1'b0;
  assign \A[19][0] [4] = 1'b0;
  assign \A[19][0] [3] = 1'b0;
  assign \A[19][0] [1] = 1'b0;
  assign \A[19][0] [0] = 1'b0;
  assign \A[19][2] [4] = 1'b0;
  assign \A[19][2] [3] = 1'b0;
  assign \A[19][2] [2] = 1'b0;
  assign \A[19][3] [4] = 1'b0;
  assign \A[19][3] [3] = 1'b0;
  assign \A[19][3] [2] = 1'b0;
  assign \A[19][3] [1] = 1'b0;
  assign \A[19][5] [4] = 1'b0;
  assign \A[19][5] [3] = 1'b0;
  assign \A[19][5] [2] = 1'b0;
  assign \A[19][5] [1] = 1'b0;
  assign \A[19][6] [4] = 1'b0;
  assign \A[19][6] [3] = 1'b0;
  assign \A[19][6] [1] = 1'b0;
  assign \A[19][6] [0] = 1'b0;
  assign \A[19][7] [4] = 1'b0;
  assign \A[19][7] [3] = 1'b0;
  assign \A[19][7] [2] = 1'b0;
  assign \A[19][7] [0] = 1'b0;
  assign \A[19][8] [4] = 1'b0;
  assign \A[19][8] [3] = 1'b0;
  assign \A[19][8] [2] = 1'b0;
  assign \A[19][8] [1] = 1'b0;
  assign \A[19][8] [0] = 1'b0;
  assign \A[19][9] [4] = 1'b0;
  assign \A[19][9] [3] = 1'b0;
  assign \A[19][9] [2] = 1'b0;
  assign \A[19][9] [1] = 1'b0;
  assign \A[19][9] [0] = 1'b0;
  assign \A[19][10] [4] = 1'b0;
  assign \A[19][10] [3] = 1'b0;
  assign \A[19][10] [2] = 1'b0;
  assign \A[19][10] [1] = 1'b0;
  assign \A[19][10] [0] = 1'b0;
  assign \A[19][11] [4] = 1'b0;
  assign \A[19][11] [3] = 1'b0;
  assign \A[19][11] [2] = 1'b0;
  assign \A[19][11] [0] = 1'b0;
  assign \A[19][12] [4] = 1'b0;
  assign \A[19][12] [3] = 1'b0;
  assign \A[19][12] [2] = 1'b0;
  assign \A[19][13] [4] = 1'b0;
  assign \A[19][13] [3] = 1'b0;
  assign \A[19][13] [2] = 1'b0;
  assign \A[19][13] [1] = 1'b0;
  assign \A[19][14] [4] = 1'b0;
  assign \A[19][14] [3] = 1'b0;
  assign \A[19][14] [2] = 1'b0;
  assign \A[19][14] [1] = 1'b0;
  assign \A[19][14] [0] = 1'b0;
  assign \A[19][15] [4] = 1'b0;
  assign \A[19][15] [3] = 1'b0;
  assign \A[19][15] [1] = 1'b0;
  assign \A[19][15] [0] = 1'b0;
  assign \A[19][16] [4] = 1'b0;
  assign \A[19][16] [3] = 1'b0;
  assign \A[19][16] [2] = 1'b0;
  assign \A[19][16] [1] = 1'b0;
  assign \A[19][17] [0] = 1'b0;
  assign \A[19][18] [4] = 1'b0;
  assign \A[19][18] [3] = 1'b0;
  assign \A[19][18] [2] = 1'b0;
  assign \A[19][18] [1] = 1'b0;
  assign \A[19][19] [4] = 1'b0;
  assign \A[19][19] [3] = 1'b0;
  assign \A[19][19] [2] = 1'b0;
  assign \A[19][19] [1] = 1'b0;
  assign \A[19][20] [4] = 1'b0;
  assign \A[19][20] [3] = 1'b0;
  assign \A[19][20] [2] = 1'b0;
  assign \A[19][20] [1] = 1'b0;
  assign \A[19][20] [0] = 1'b0;
  assign \A[19][21] [4] = 1'b0;
  assign \A[19][21] [3] = 1'b0;
  assign \A[19][21] [2] = 1'b0;
  assign \A[19][21] [0] = 1'b0;
  assign \A[19][22] [4] = 1'b0;
  assign \A[19][22] [3] = 1'b0;
  assign \A[19][22] [2] = 1'b0;
  assign \A[19][22] [0] = 1'b0;
  assign \A[19][24] [4] = 1'b0;
  assign \A[19][24] [3] = 1'b0;
  assign \A[19][24] [2] = 1'b0;
  assign \A[19][24] [1] = 1'b0;
  assign \A[19][25] [4] = 1'b0;
  assign \A[19][25] [3] = 1'b0;
  assign \A[19][25] [2] = 1'b0;
  assign \A[19][25] [0] = 1'b0;
  assign \A[19][26] [1] = 1'b0;
  assign \A[19][26] [0] = 1'b0;
  assign \A[19][27] [4] = 1'b0;
  assign \A[19][27] [3] = 1'b0;
  assign \A[19][27] [2] = 1'b0;
  assign \A[19][27] [0] = 1'b0;
  assign \A[19][30] [4] = 1'b0;
  assign \A[19][30] [3] = 1'b0;
  assign \A[19][30] [2] = 1'b0;
  assign \A[19][30] [1] = 1'b0;
  assign \A[19][31] [1] = 1'b0;
  assign \A[19][32] [4] = 1'b0;
  assign \A[19][32] [3] = 1'b0;
  assign \A[19][32] [2] = 1'b0;
  assign \A[19][32] [1] = 1'b0;
  assign \A[19][35] [4] = 1'b0;
  assign \A[19][35] [3] = 1'b0;
  assign \A[19][35] [2] = 1'b0;
  assign \A[19][35] [1] = 1'b0;
  assign \A[19][35] [0] = 1'b0;
  assign \A[19][36] [4] = 1'b0;
  assign \A[19][36] [3] = 1'b0;
  assign \A[19][36] [2] = 1'b0;
  assign \A[19][36] [1] = 1'b0;
  assign \A[19][37] [1] = 1'b0;
  assign \A[19][38] [4] = 1'b0;
  assign \A[19][38] [3] = 1'b0;
  assign \A[19][38] [2] = 1'b0;
  assign \A[19][38] [1] = 1'b0;
  assign \A[19][38] [0] = 1'b0;
  assign \A[19][39] [4] = 1'b0;
  assign \A[19][39] [3] = 1'b0;
  assign \A[19][39] [1] = 1'b0;
  assign \A[19][39] [0] = 1'b0;
  assign \A[19][40] [4] = 1'b0;
  assign \A[19][40] [3] = 1'b0;
  assign \A[19][40] [2] = 1'b0;
  assign \A[19][40] [1] = 1'b0;
  assign \A[19][40] [0] = 1'b0;
  assign \A[19][42] [4] = 1'b0;
  assign \A[19][42] [3] = 1'b0;
  assign \A[19][42] [2] = 1'b0;
  assign \A[19][42] [1] = 1'b0;
  assign \A[19][42] [0] = 1'b0;
  assign \A[19][43] [4] = 1'b0;
  assign \A[19][43] [3] = 1'b0;
  assign \A[19][43] [2] = 1'b0;
  assign \A[19][43] [1] = 1'b0;
  assign \A[19][43] [0] = 1'b0;
  assign \A[19][44] [1] = 1'b0;
  assign \A[19][45] [4] = 1'b0;
  assign \A[19][45] [3] = 1'b0;
  assign \A[19][45] [2] = 1'b0;
  assign \A[19][45] [0] = 1'b0;
  assign \A[19][46] [1] = 1'b0;
  assign \A[19][46] [0] = 1'b0;
  assign \A[19][47] [0] = 1'b0;
  assign \A[19][48] [0] = 1'b0;
  assign \A[19][49] [0] = 1'b0;
  assign \A[19][50] [4] = 1'b0;
  assign \A[19][50] [3] = 1'b0;
  assign \A[19][50] [2] = 1'b0;
  assign \A[19][50] [1] = 1'b0;
  assign \A[19][50] [0] = 1'b0;
  assign \A[19][51] [4] = 1'b0;
  assign \A[19][51] [3] = 1'b0;
  assign \A[19][51] [2] = 1'b0;
  assign \A[19][51] [1] = 1'b0;
  assign \A[19][51] [0] = 1'b0;
  assign \A[19][53] [4] = 1'b0;
  assign \A[19][53] [3] = 1'b0;
  assign \A[19][53] [2] = 1'b0;
  assign \A[19][53] [1] = 1'b0;
  assign \A[19][53] [0] = 1'b0;
  assign \A[19][54] [0] = 1'b0;
  assign \A[19][55] [4] = 1'b0;
  assign \A[19][55] [3] = 1'b0;
  assign \A[19][55] [2] = 1'b0;
  assign \A[19][55] [1] = 1'b0;
  assign \A[19][55] [0] = 1'b0;
  assign \A[19][56] [1] = 1'b0;
  assign \A[19][57] [1] = 1'b0;
  assign \A[19][57] [0] = 1'b0;
  assign \A[19][58] [0] = 1'b0;
  assign \A[19][59] [2] = 1'b0;
  assign \A[19][59] [0] = 1'b0;
  assign \A[19][60] [1] = 1'b0;
  assign \A[19][60] [0] = 1'b0;
  assign \A[19][61] [0] = 1'b0;
  assign \A[19][62] [0] = 1'b0;
  assign \A[19][63] [4] = 1'b0;
  assign \A[19][63] [3] = 1'b0;
  assign \A[19][63] [2] = 1'b0;
  assign \A[19][63] [1] = 1'b0;
  assign \A[19][63] [0] = 1'b0;
  assign \A[19][64] [4] = 1'b0;
  assign \A[19][64] [3] = 1'b0;
  assign \A[19][64] [2] = 1'b0;
  assign \A[19][64] [1] = 1'b0;
  assign \A[19][64] [0] = 1'b0;
  assign \A[19][67] [4] = 1'b0;
  assign \A[19][67] [3] = 1'b0;
  assign \A[19][67] [2] = 1'b0;
  assign \A[19][67] [1] = 1'b0;
  assign \A[19][67] [0] = 1'b0;
  assign \A[19][73] [1] = 1'b0;
  assign \A[19][74] [4] = 1'b0;
  assign \A[19][74] [3] = 1'b0;
  assign \A[19][74] [2] = 1'b0;
  assign \A[19][74] [0] = 1'b0;
  assign \A[19][76] [1] = 1'b0;
  assign \A[19][77] [2] = 1'b0;
  assign \A[19][78] [2] = 1'b0;
  assign \A[19][78] [1] = 1'b0;
  assign \A[19][79] [2] = 1'b0;
  assign \A[19][80] [0] = 1'b0;
  assign \A[19][82] [1] = 1'b0;
  assign \A[19][82] [0] = 1'b0;
  assign \A[19][83] [0] = 1'b0;
  assign \A[19][84] [4] = 1'b0;
  assign \A[19][84] [3] = 1'b0;
  assign \A[19][84] [2] = 1'b0;
  assign \A[19][84] [1] = 1'b0;
  assign \A[19][86] [4] = 1'b0;
  assign \A[19][86] [3] = 1'b0;
  assign \A[19][86] [2] = 1'b0;
  assign \A[19][86] [0] = 1'b0;
  assign \A[19][87] [2] = 1'b0;
  assign \A[19][89] [4] = 1'b0;
  assign \A[19][89] [3] = 1'b0;
  assign \A[19][89] [2] = 1'b0;
  assign \A[19][89] [1] = 1'b0;
  assign \A[19][89] [0] = 1'b0;
  assign \A[19][91] [0] = 1'b0;
  assign \A[19][93] [0] = 1'b0;
  assign \A[19][94] [2] = 1'b0;
  assign \A[19][94] [1] = 1'b0;
  assign \A[19][94] [0] = 1'b0;
  assign \A[19][95] [1] = 1'b0;
  assign \A[19][95] [0] = 1'b0;
  assign \A[19][97] [4] = 1'b0;
  assign \A[19][97] [3] = 1'b0;
  assign \A[19][97] [2] = 1'b0;
  assign \A[19][97] [1] = 1'b0;
  assign \A[19][98] [4] = 1'b0;
  assign \A[19][98] [3] = 1'b0;
  assign \A[19][98] [2] = 1'b0;
  assign \A[19][98] [1] = 1'b0;
  assign \A[19][98] [0] = 1'b0;
  assign \A[19][99] [4] = 1'b0;
  assign \A[19][99] [3] = 1'b0;
  assign \A[19][99] [2] = 1'b0;
  assign \A[19][99] [1] = 1'b0;
  assign \A[19][99] [0] = 1'b0;
  assign \A[19][100] [0] = 1'b0;
  assign \A[19][101] [4] = 1'b0;
  assign \A[19][101] [3] = 1'b0;
  assign \A[19][101] [2] = 1'b0;
  assign \A[19][101] [1] = 1'b0;
  assign \A[19][101] [0] = 1'b0;
  assign \A[19][103] [4] = 1'b0;
  assign \A[19][103] [3] = 1'b0;
  assign \A[19][103] [2] = 1'b0;
  assign \A[19][103] [1] = 1'b0;
  assign \A[19][103] [0] = 1'b0;
  assign \A[19][105] [4] = 1'b0;
  assign \A[19][105] [3] = 1'b0;
  assign \A[19][105] [2] = 1'b0;
  assign \A[19][105] [1] = 1'b0;
  assign \A[19][105] [0] = 1'b0;
  assign \A[19][107] [4] = 1'b0;
  assign \A[19][107] [3] = 1'b0;
  assign \A[19][107] [2] = 1'b0;
  assign \A[19][107] [1] = 1'b0;
  assign \A[19][107] [0] = 1'b0;
  assign \A[19][109] [4] = 1'b0;
  assign \A[19][109] [3] = 1'b0;
  assign \A[19][109] [2] = 1'b0;
  assign \A[19][109] [1] = 1'b0;
  assign \A[19][109] [0] = 1'b0;
  assign \A[19][110] [1] = 1'b0;
  assign \A[19][110] [0] = 1'b0;
  assign \A[19][111] [2] = 1'b0;
  assign \A[19][111] [1] = 1'b0;
  assign \A[19][112] [4] = 1'b0;
  assign \A[19][112] [3] = 1'b0;
  assign \A[19][112] [2] = 1'b0;
  assign \A[19][112] [1] = 1'b0;
  assign \A[19][112] [0] = 1'b0;
  assign \A[19][113] [4] = 1'b0;
  assign \A[19][113] [3] = 1'b0;
  assign \A[19][113] [2] = 1'b0;
  assign \A[19][113] [1] = 1'b0;
  assign \A[19][113] [0] = 1'b0;
  assign \A[19][114] [4] = 1'b0;
  assign \A[19][114] [3] = 1'b0;
  assign \A[19][114] [2] = 1'b0;
  assign \A[19][114] [1] = 1'b0;
  assign \A[19][116] [4] = 1'b0;
  assign \A[19][116] [3] = 1'b0;
  assign \A[19][116] [2] = 1'b0;
  assign \A[19][116] [1] = 1'b0;
  assign \A[19][116] [0] = 1'b0;
  assign \A[19][117] [4] = 1'b0;
  assign \A[19][117] [3] = 1'b0;
  assign \A[19][117] [2] = 1'b0;
  assign \A[19][117] [1] = 1'b0;
  assign \A[19][119] [0] = 1'b0;
  assign \A[19][120] [0] = 1'b0;
  assign \A[19][121] [4] = 1'b0;
  assign \A[19][121] [3] = 1'b0;
  assign \A[19][121] [2] = 1'b0;
  assign \A[19][121] [1] = 1'b0;
  assign \A[19][121] [0] = 1'b0;
  assign \A[19][122] [4] = 1'b0;
  assign \A[19][122] [3] = 1'b0;
  assign \A[19][122] [2] = 1'b0;
  assign \A[19][122] [1] = 1'b0;
  assign \A[19][122] [0] = 1'b0;
  assign \A[19][124] [4] = 1'b0;
  assign \A[19][124] [3] = 1'b0;
  assign \A[19][124] [2] = 1'b0;
  assign \A[19][124] [1] = 1'b0;
  assign \A[19][124] [0] = 1'b0;
  assign \A[19][125] [4] = 1'b0;
  assign \A[19][125] [3] = 1'b0;
  assign \A[19][125] [2] = 1'b0;
  assign \A[19][125] [1] = 1'b0;
  assign \A[19][126] [4] = 1'b0;
  assign \A[19][126] [3] = 1'b0;
  assign \A[19][126] [2] = 1'b0;
  assign \A[19][126] [1] = 1'b0;
  assign \A[19][126] [0] = 1'b0;
  assign \A[19][128] [1] = 1'b0;
  assign \A[19][129] [4] = 1'b0;
  assign \A[19][129] [3] = 1'b0;
  assign \A[19][129] [2] = 1'b0;
  assign \A[19][129] [1] = 1'b0;
  assign \A[19][129] [0] = 1'b0;
  assign \A[19][130] [4] = 1'b0;
  assign \A[19][130] [3] = 1'b0;
  assign \A[19][130] [2] = 1'b0;
  assign \A[19][130] [1] = 1'b0;
  assign \A[19][131] [4] = 1'b0;
  assign \A[19][131] [3] = 1'b0;
  assign \A[19][131] [2] = 1'b0;
  assign \A[19][131] [1] = 1'b0;
  assign \A[19][132] [0] = 1'b0;
  assign \A[19][134] [0] = 1'b0;
  assign \A[19][135] [4] = 1'b0;
  assign \A[19][135] [3] = 1'b0;
  assign \A[19][135] [2] = 1'b0;
  assign \A[19][135] [1] = 1'b0;
  assign \A[19][135] [0] = 1'b0;
  assign \A[19][136] [0] = 1'b0;
  assign \A[19][137] [4] = 1'b0;
  assign \A[19][137] [3] = 1'b0;
  assign \A[19][137] [2] = 1'b0;
  assign \A[19][137] [1] = 1'b0;
  assign \A[19][137] [0] = 1'b0;
  assign \A[19][138] [4] = 1'b0;
  assign \A[19][138] [3] = 1'b0;
  assign \A[19][138] [2] = 1'b0;
  assign \A[19][140] [4] = 1'b0;
  assign \A[19][140] [3] = 1'b0;
  assign \A[19][140] [2] = 1'b0;
  assign \A[19][140] [1] = 1'b0;
  assign \A[19][142] [4] = 1'b0;
  assign \A[19][142] [3] = 1'b0;
  assign \A[19][142] [2] = 1'b0;
  assign \A[19][142] [1] = 1'b0;
  assign \A[19][142] [0] = 1'b0;
  assign \A[19][144] [2] = 1'b0;
  assign \A[19][145] [1] = 1'b0;
  assign \A[19][146] [4] = 1'b0;
  assign \A[19][146] [3] = 1'b0;
  assign \A[19][146] [2] = 1'b0;
  assign \A[19][146] [1] = 1'b0;
  assign \A[19][147] [0] = 1'b0;
  assign \A[19][148] [4] = 1'b0;
  assign \A[19][148] [3] = 1'b0;
  assign \A[19][148] [2] = 1'b0;
  assign \A[19][148] [1] = 1'b0;
  assign \A[19][148] [0] = 1'b0;
  assign \A[19][149] [4] = 1'b0;
  assign \A[19][149] [3] = 1'b0;
  assign \A[19][149] [2] = 1'b0;
  assign \A[19][149] [1] = 1'b0;
  assign \A[19][149] [0] = 1'b0;
  assign \A[19][150] [4] = 1'b0;
  assign \A[19][150] [3] = 1'b0;
  assign \A[19][150] [2] = 1'b0;
  assign \A[19][150] [1] = 1'b0;
  assign \A[19][153] [4] = 1'b0;
  assign \A[19][153] [3] = 1'b0;
  assign \A[19][153] [2] = 1'b0;
  assign \A[19][153] [1] = 1'b0;
  assign \A[19][153] [0] = 1'b0;
  assign \A[19][156] [4] = 1'b0;
  assign \A[19][156] [3] = 1'b0;
  assign \A[19][156] [2] = 1'b0;
  assign \A[19][156] [1] = 1'b0;
  assign \A[19][156] [0] = 1'b0;
  assign \A[19][158] [4] = 1'b0;
  assign \A[19][158] [3] = 1'b0;
  assign \A[19][158] [2] = 1'b0;
  assign \A[19][158] [1] = 1'b0;
  assign \A[19][158] [0] = 1'b0;
  assign \A[19][159] [4] = 1'b0;
  assign \A[19][159] [3] = 1'b0;
  assign \A[19][159] [2] = 1'b0;
  assign \A[19][159] [1] = 1'b0;
  assign \A[19][159] [0] = 1'b0;
  assign \A[19][160] [0] = 1'b0;
  assign \A[19][161] [0] = 1'b0;
  assign \A[19][163] [4] = 1'b0;
  assign \A[19][163] [3] = 1'b0;
  assign \A[19][163] [2] = 1'b0;
  assign \A[19][163] [1] = 1'b0;
  assign \A[19][163] [0] = 1'b0;
  assign \A[19][164] [4] = 1'b0;
  assign \A[19][164] [3] = 1'b0;
  assign \A[19][164] [2] = 1'b0;
  assign \A[19][164] [1] = 1'b0;
  assign \A[19][164] [0] = 1'b0;
  assign \A[19][165] [4] = 1'b0;
  assign \A[19][165] [3] = 1'b0;
  assign \A[19][165] [2] = 1'b0;
  assign \A[19][165] [1] = 1'b0;
  assign \A[19][166] [4] = 1'b0;
  assign \A[19][166] [3] = 1'b0;
  assign \A[19][166] [2] = 1'b0;
  assign \A[19][166] [1] = 1'b0;
  assign \A[19][166] [0] = 1'b0;
  assign \A[19][167] [4] = 1'b0;
  assign \A[19][167] [3] = 1'b0;
  assign \A[19][167] [2] = 1'b0;
  assign \A[19][167] [1] = 1'b0;
  assign \A[19][167] [0] = 1'b0;
  assign \A[19][169] [4] = 1'b0;
  assign \A[19][169] [3] = 1'b0;
  assign \A[19][169] [2] = 1'b0;
  assign \A[19][169] [1] = 1'b0;
  assign \A[19][169] [0] = 1'b0;
  assign \A[19][170] [4] = 1'b0;
  assign \A[19][170] [3] = 1'b0;
  assign \A[19][170] [2] = 1'b0;
  assign \A[19][170] [1] = 1'b0;
  assign \A[19][171] [4] = 1'b0;
  assign \A[19][171] [3] = 1'b0;
  assign \A[19][171] [2] = 1'b0;
  assign \A[19][171] [1] = 1'b0;
  assign \A[19][171] [0] = 1'b0;
  assign \A[19][172] [4] = 1'b0;
  assign \A[19][172] [3] = 1'b0;
  assign \A[19][172] [2] = 1'b0;
  assign \A[19][172] [1] = 1'b0;
  assign \A[19][172] [0] = 1'b0;
  assign \A[19][173] [1] = 1'b0;
  assign \A[19][174] [0] = 1'b0;
  assign \A[19][175] [4] = 1'b0;
  assign \A[19][175] [3] = 1'b0;
  assign \A[19][175] [2] = 1'b0;
  assign \A[19][175] [1] = 1'b0;
  assign \A[19][175] [0] = 1'b0;
  assign \A[19][176] [0] = 1'b0;
  assign \A[19][177] [4] = 1'b0;
  assign \A[19][177] [3] = 1'b0;
  assign \A[19][177] [2] = 1'b0;
  assign \A[19][177] [1] = 1'b0;
  assign \A[19][177] [0] = 1'b0;
  assign \A[19][178] [0] = 1'b0;
  assign \A[19][179] [0] = 1'b0;
  assign \A[19][180] [4] = 1'b0;
  assign \A[19][180] [3] = 1'b0;
  assign \A[19][180] [2] = 1'b0;
  assign \A[19][180] [1] = 1'b0;
  assign \A[19][180] [0] = 1'b0;
  assign \A[19][184] [1] = 1'b0;
  assign \A[19][185] [4] = 1'b0;
  assign \A[19][185] [3] = 1'b0;
  assign \A[19][185] [2] = 1'b0;
  assign \A[19][185] [1] = 1'b0;
  assign \A[19][185] [0] = 1'b0;
  assign \A[19][186] [4] = 1'b0;
  assign \A[19][186] [3] = 1'b0;
  assign \A[19][186] [2] = 1'b0;
  assign \A[19][186] [1] = 1'b0;
  assign \A[19][186] [0] = 1'b0;
  assign \A[19][187] [4] = 1'b0;
  assign \A[19][187] [3] = 1'b0;
  assign \A[19][187] [2] = 1'b0;
  assign \A[19][187] [0] = 1'b0;
  assign \A[19][188] [0] = 1'b0;
  assign \A[19][189] [4] = 1'b0;
  assign \A[19][189] [3] = 1'b0;
  assign \A[19][189] [2] = 1'b0;
  assign \A[19][189] [1] = 1'b0;
  assign \A[19][190] [4] = 1'b0;
  assign \A[19][190] [3] = 1'b0;
  assign \A[19][190] [2] = 1'b0;
  assign \A[19][190] [0] = 1'b0;
  assign \A[19][191] [4] = 1'b0;
  assign \A[19][191] [3] = 1'b0;
  assign \A[19][191] [2] = 1'b0;
  assign \A[19][191] [0] = 1'b0;
  assign \A[19][192] [4] = 1'b0;
  assign \A[19][192] [3] = 1'b0;
  assign \A[19][192] [2] = 1'b0;
  assign \A[19][192] [0] = 1'b0;
  assign \A[19][193] [4] = 1'b0;
  assign \A[19][193] [3] = 1'b0;
  assign \A[19][193] [2] = 1'b0;
  assign \A[19][193] [1] = 1'b0;
  assign \A[19][194] [4] = 1'b0;
  assign \A[19][194] [3] = 1'b0;
  assign \A[19][194] [2] = 1'b0;
  assign \A[19][194] [1] = 1'b0;
  assign \A[19][194] [0] = 1'b0;
  assign \A[19][195] [1] = 1'b0;
  assign \A[19][196] [4] = 1'b0;
  assign \A[19][196] [3] = 1'b0;
  assign \A[19][196] [2] = 1'b0;
  assign \A[19][196] [1] = 1'b0;
  assign \A[19][196] [0] = 1'b0;
  assign \A[19][198] [4] = 1'b0;
  assign \A[19][198] [3] = 1'b0;
  assign \A[19][198] [2] = 1'b0;
  assign \A[19][198] [0] = 1'b0;
  assign \A[19][200] [4] = 1'b0;
  assign \A[19][200] [3] = 1'b0;
  assign \A[19][200] [2] = 1'b0;
  assign \A[19][200] [1] = 1'b0;
  assign \A[19][200] [0] = 1'b0;
  assign \A[19][201] [1] = 1'b0;
  assign \A[19][201] [0] = 1'b0;
  assign \A[19][202] [0] = 1'b0;
  assign \A[19][203] [4] = 1'b0;
  assign \A[19][203] [3] = 1'b0;
  assign \A[19][203] [2] = 1'b0;
  assign \A[19][203] [1] = 1'b0;
  assign \A[19][203] [0] = 1'b0;
  assign \A[19][204] [4] = 1'b0;
  assign \A[19][204] [3] = 1'b0;
  assign \A[19][204] [2] = 1'b0;
  assign \A[19][204] [1] = 1'b0;
  assign \A[19][205] [4] = 1'b0;
  assign \A[19][205] [3] = 1'b0;
  assign \A[19][205] [2] = 1'b0;
  assign \A[19][205] [0] = 1'b0;
  assign \A[19][207] [4] = 1'b0;
  assign \A[19][207] [3] = 1'b0;
  assign \A[19][207] [2] = 1'b0;
  assign \A[19][207] [0] = 1'b0;
  assign \A[19][209] [4] = 1'b0;
  assign \A[19][209] [3] = 1'b0;
  assign \A[19][209] [2] = 1'b0;
  assign \A[19][209] [1] = 1'b0;
  assign \A[19][209] [0] = 1'b0;
  assign \A[19][210] [0] = 1'b0;
  assign \A[19][211] [4] = 1'b0;
  assign \A[19][211] [3] = 1'b0;
  assign \A[19][211] [2] = 1'b0;
  assign \A[19][211] [0] = 1'b0;
  assign \A[19][212] [4] = 1'b0;
  assign \A[19][212] [3] = 1'b0;
  assign \A[19][212] [2] = 1'b0;
  assign \A[19][212] [1] = 1'b0;
  assign \A[19][213] [4] = 1'b0;
  assign \A[19][213] [3] = 1'b0;
  assign \A[19][213] [2] = 1'b0;
  assign \A[19][213] [1] = 1'b0;
  assign \A[19][214] [0] = 1'b0;
  assign \A[19][215] [4] = 1'b0;
  assign \A[19][215] [3] = 1'b0;
  assign \A[19][215] [2] = 1'b0;
  assign \A[19][216] [4] = 1'b0;
  assign \A[19][216] [3] = 1'b0;
  assign \A[19][216] [2] = 1'b0;
  assign \A[19][216] [1] = 1'b0;
  assign \A[19][216] [0] = 1'b0;
  assign \A[19][217] [4] = 1'b0;
  assign \A[19][217] [3] = 1'b0;
  assign \A[19][217] [2] = 1'b0;
  assign \A[19][217] [1] = 1'b0;
  assign \A[19][219] [0] = 1'b0;
  assign \A[19][220] [4] = 1'b0;
  assign \A[19][220] [3] = 1'b0;
  assign \A[19][220] [2] = 1'b0;
  assign \A[19][220] [1] = 1'b0;
  assign \A[19][220] [0] = 1'b0;
  assign \A[19][223] [4] = 1'b0;
  assign \A[19][223] [3] = 1'b0;
  assign \A[19][223] [2] = 1'b0;
  assign \A[19][223] [1] = 1'b0;
  assign \A[19][223] [0] = 1'b0;
  assign \A[19][224] [0] = 1'b0;
  assign \A[19][225] [4] = 1'b0;
  assign \A[19][225] [3] = 1'b0;
  assign \A[19][225] [2] = 1'b0;
  assign \A[19][225] [1] = 1'b0;
  assign \A[19][225] [0] = 1'b0;
  assign \A[19][226] [4] = 1'b0;
  assign \A[19][226] [3] = 1'b0;
  assign \A[19][226] [2] = 1'b0;
  assign \A[19][226] [1] = 1'b0;
  assign \A[19][226] [0] = 1'b0;
  assign \A[19][227] [4] = 1'b0;
  assign \A[19][227] [3] = 1'b0;
  assign \A[19][227] [2] = 1'b0;
  assign \A[19][228] [4] = 1'b0;
  assign \A[19][228] [3] = 1'b0;
  assign \A[19][228] [2] = 1'b0;
  assign \A[19][228] [1] = 1'b0;
  assign \A[19][228] [0] = 1'b0;
  assign \A[19][229] [0] = 1'b0;
  assign \A[19][230] [4] = 1'b0;
  assign \A[19][230] [3] = 1'b0;
  assign \A[19][230] [2] = 1'b0;
  assign \A[19][230] [1] = 1'b0;
  assign \A[19][230] [0] = 1'b0;
  assign \A[19][231] [4] = 1'b0;
  assign \A[19][231] [3] = 1'b0;
  assign \A[19][231] [2] = 1'b0;
  assign \A[19][231] [0] = 1'b0;
  assign \A[19][232] [1] = 1'b0;
  assign \A[19][233] [4] = 1'b0;
  assign \A[19][233] [3] = 1'b0;
  assign \A[19][233] [2] = 1'b0;
  assign \A[19][233] [1] = 1'b0;
  assign \A[19][234] [4] = 1'b0;
  assign \A[19][234] [3] = 1'b0;
  assign \A[19][234] [2] = 1'b0;
  assign \A[19][234] [0] = 1'b0;
  assign \A[19][236] [4] = 1'b0;
  assign \A[19][236] [3] = 1'b0;
  assign \A[19][236] [2] = 1'b0;
  assign \A[19][236] [1] = 1'b0;
  assign \A[19][237] [4] = 1'b0;
  assign \A[19][237] [3] = 1'b0;
  assign \A[19][237] [2] = 1'b0;
  assign \A[19][237] [1] = 1'b0;
  assign \A[19][238] [1] = 1'b0;
  assign \A[19][239] [4] = 1'b0;
  assign \A[19][239] [3] = 1'b0;
  assign \A[19][239] [2] = 1'b0;
  assign \A[19][239] [1] = 1'b0;
  assign \A[19][239] [0] = 1'b0;
  assign \A[19][240] [4] = 1'b0;
  assign \A[19][240] [3] = 1'b0;
  assign \A[19][240] [2] = 1'b0;
  assign \A[19][240] [1] = 1'b0;
  assign \A[19][240] [0] = 1'b0;
  assign \A[19][241] [4] = 1'b0;
  assign \A[19][241] [3] = 1'b0;
  assign \A[19][241] [2] = 1'b0;
  assign \A[19][241] [1] = 1'b0;
  assign \A[19][241] [0] = 1'b0;
  assign \A[19][242] [4] = 1'b0;
  assign \A[19][242] [3] = 1'b0;
  assign \A[19][242] [2] = 1'b0;
  assign \A[19][242] [0] = 1'b0;
  assign \A[19][243] [4] = 1'b0;
  assign \A[19][243] [3] = 1'b0;
  assign \A[19][243] [2] = 1'b0;
  assign \A[19][243] [1] = 1'b0;
  assign \A[19][243] [0] = 1'b0;
  assign \A[19][244] [0] = 1'b0;
  assign \A[19][245] [4] = 1'b0;
  assign \A[19][245] [3] = 1'b0;
  assign \A[19][245] [2] = 1'b0;
  assign \A[19][245] [1] = 1'b0;
  assign \A[19][245] [0] = 1'b0;
  assign \A[19][246] [4] = 1'b0;
  assign \A[19][246] [3] = 1'b0;
  assign \A[19][246] [2] = 1'b0;
  assign \A[19][246] [1] = 1'b0;
  assign \A[19][247] [4] = 1'b0;
  assign \A[19][247] [3] = 1'b0;
  assign \A[19][247] [2] = 1'b0;
  assign \A[19][247] [1] = 1'b0;
  assign \A[19][247] [0] = 1'b0;
  assign \A[19][248] [1] = 1'b0;
  assign \A[19][249] [4] = 1'b0;
  assign \A[19][249] [3] = 1'b0;
  assign \A[19][249] [2] = 1'b0;
  assign \A[19][249] [1] = 1'b0;
  assign \A[19][249] [0] = 1'b0;
  assign \A[19][250] [4] = 1'b0;
  assign \A[19][250] [3] = 1'b0;
  assign \A[19][250] [2] = 1'b0;
  assign \A[19][250] [1] = 1'b0;
  assign \A[19][251] [4] = 1'b0;
  assign \A[19][251] [3] = 1'b0;
  assign \A[19][251] [2] = 1'b0;
  assign \A[19][251] [1] = 1'b0;
  assign \A[19][251] [0] = 1'b0;
  assign \A[19][252] [4] = 1'b0;
  assign \A[19][252] [3] = 1'b0;
  assign \A[19][252] [2] = 1'b0;
  assign \A[19][252] [1] = 1'b0;
  assign \A[19][253] [0] = 1'b0;
  assign \A[19][255] [4] = 1'b0;
  assign \A[19][255] [3] = 1'b0;
  assign \A[19][255] [2] = 1'b0;
  assign \A[19][255] [1] = 1'b0;
  assign \A[19][255] [0] = 1'b0;
  assign \biases_l1[0] [6] = 1'b1;
  assign \biases_l1[0] [5] = 1'b1;
  assign \biases_l1[0] [4] = 1'b1;
  assign \biases_l1[0] [1] = 1'b1;
  assign \biases_l1[0] [0] = 1'b1;
  assign \biases_l1[1] [6] = 1'b1;
  assign \biases_l1[1] [5] = 1'b1;
  assign \biases_l1[1] [4] = 1'b1;
  assign \biases_l1[1] [3] = 1'b1;
  assign \biases_l1[1] [0] = 1'b1;
  assign \biases_l1[2] [4] = 1'b1;
  assign \biases_l1[2] [1] = 1'b1;
  assign \biases_l1[2] [0] = 1'b1;
  assign \biases_l1[3] [6] = 1'b1;
  assign \biases_l1[3] [5] = 1'b1;
  assign \biases_l1[3] [4] = 1'b1;
  assign \biases_l1[3] [3] = 1'b1;
  assign \biases_l1[4] [3] = 1'b1;
  assign \biases_l1[4] [1] = 1'b1;
  assign \biases_l1[4] [0] = 1'b1;
  assign \biases_l1[5] [2] = 1'b1;
  assign \biases_l1[5] [0] = 1'b1;
  assign \biases_l1[6] [1] = 1'b1;
  assign \biases_l1[6] [0] = 1'b1;
  assign \biases_l1[7] [3] = 1'b1;
  assign \biases_l1[7] [0] = 1'b1;
  assign \biases_l1[8] [4] = 1'b1;
  assign \biases_l1[8] [3] = 1'b1;
  assign \biases_l1[8] [2] = 1'b1;
  assign \biases_l1[8] [0] = 1'b1;
  assign \biases_l1[9] [4] = 1'b1;
  assign \biases_l1[9] [2] = 1'b1;
  assign \biases_l1[9] [1] = 1'b1;
  assign \biases_l1[10] [6] = 1'b1;
  assign \biases_l1[10] [5] = 1'b1;
  assign \biases_l1[10] [2] = 1'b1;
  assign \biases_l1[10] [1] = 1'b1;
  assign \biases_l1[10] [0] = 1'b1;
  assign \biases_l1[11] [2] = 1'b1;
  assign \biases_l1[11] [0] = 1'b1;
  assign \biases_l1[12] [6] = 1'b1;
  assign \biases_l1[12] [5] = 1'b1;
  assign \biases_l1[12] [3] = 1'b1;
  assign \biases_l1[12] [2] = 1'b1;
  assign \biases_l1[13] [6] = 1'b1;
  assign \biases_l1[13] [5] = 1'b1;
  assign \biases_l1[14] [6] = 1'b1;
  assign \biases_l1[14] [5] = 1'b1;
  assign \biases_l1[14] [3] = 1'b1;
  assign \biases_l1[14] [2] = 1'b1;
  assign \biases_l1[14] [0] = 1'b1;
  assign \biases_l1[15] [6] = 1'b1;
  assign \biases_l1[15] [4] = 1'b1;
  assign \biases_l1[15] [3] = 1'b1;
  assign \biases_l1[15] [2] = 1'b1;
  assign \biases_l1[15] [0] = 1'b1;
  assign \biases_l1[16] [6] = 1'b1;
  assign \biases_l1[16] [5] = 1'b1;
  assign \biases_l1[16] [3] = 1'b1;
  assign \biases_l1[16] [2] = 1'b1;
  assign \biases_l1[16] [1] = 1'b1;
  assign \biases_l1[17] [4] = 1'b1;
  assign \biases_l1[17] [1] = 1'b1;
  assign \biases_l1[18] [6] = 1'b1;
  assign \biases_l1[18] [5] = 1'b1;
  assign \biases_l1[18] [4] = 1'b1;
  assign \biases_l1[18] [3] = 1'b1;
  assign \biases_l1[18] [1] = 1'b1;
  assign \biases_l1[19] [5] = 1'b1;
  assign \biases_l1[19] [3] = 1'b1;
  assign \biases_l1[19] [0] = 1'b1;
  assign \A[0][0] [0] = 1'b1;
  assign \A[0][1] [0] = 1'b1;
  assign \A[0][3] [4] = 1'b1;
  assign \A[0][3] [3] = 1'b1;
  assign \A[0][3] [2] = 1'b1;
  assign \A[0][3] [1] = 1'b1;
  assign \A[0][4] [0] = 1'b1;
  assign \A[0][5] [0] = 1'b1;
  assign \A[0][6] [2] = 1'b1;
  assign \A[0][7] [4] = 1'b1;
  assign \A[0][7] [3] = 1'b1;
  assign \A[0][7] [2] = 1'b1;
  assign \A[0][7] [1] = 1'b1;
  assign \A[0][7] [0] = 1'b1;
  assign \A[0][8] [4] = 1'b1;
  assign \A[0][8] [3] = 1'b1;
  assign \A[0][8] [2] = 1'b1;
  assign \A[0][8] [1] = 1'b1;
  assign \A[0][8] [0] = 1'b1;
  assign \A[0][9] [4] = 1'b1;
  assign \A[0][9] [3] = 1'b1;
  assign \A[0][9] [2] = 1'b1;
  assign \A[0][9] [0] = 1'b1;
  assign \A[0][11] [4] = 1'b1;
  assign \A[0][11] [3] = 1'b1;
  assign \A[0][11] [2] = 1'b1;
  assign \A[0][11] [1] = 1'b1;
  assign \A[0][12] [4] = 1'b1;
  assign \A[0][12] [3] = 1'b1;
  assign \A[0][12] [2] = 1'b1;
  assign \A[0][12] [1] = 1'b1;
  assign \A[0][13] [0] = 1'b1;
  assign \A[0][14] [0] = 1'b1;
  assign \A[0][16] [4] = 1'b1;
  assign \A[0][16] [3] = 1'b1;
  assign \A[0][16] [2] = 1'b1;
  assign \A[0][16] [1] = 1'b1;
  assign \A[0][16] [0] = 1'b1;
  assign \A[0][17] [4] = 1'b1;
  assign \A[0][17] [3] = 1'b1;
  assign \A[0][17] [2] = 1'b1;
  assign \A[0][17] [1] = 1'b1;
  assign \A[0][18] [4] = 1'b1;
  assign \A[0][18] [3] = 1'b1;
  assign \A[0][18] [2] = 1'b1;
  assign \A[0][18] [1] = 1'b1;
  assign \A[0][18] [0] = 1'b1;
  assign \A[0][19] [1] = 1'b1;
  assign \A[0][19] [0] = 1'b1;
  assign \A[0][21] [4] = 1'b1;
  assign \A[0][21] [3] = 1'b1;
  assign \A[0][21] [2] = 1'b1;
  assign \A[0][21] [1] = 1'b1;
  assign \A[0][21] [0] = 1'b1;
  assign \A[0][22] [0] = 1'b1;
  assign \A[0][23] [4] = 1'b1;
  assign \A[0][23] [3] = 1'b1;
  assign \A[0][23] [2] = 1'b1;
  assign \A[0][23] [1] = 1'b1;
  assign \A[0][23] [0] = 1'b1;
  assign \A[0][26] [4] = 1'b1;
  assign \A[0][26] [3] = 1'b1;
  assign \A[0][26] [2] = 1'b1;
  assign \A[0][26] [1] = 1'b1;
  assign \A[0][27] [0] = 1'b1;
  assign \A[0][28] [4] = 1'b1;
  assign \A[0][28] [3] = 1'b1;
  assign \A[0][28] [2] = 1'b1;
  assign \A[0][28] [1] = 1'b1;
  assign \A[0][28] [0] = 1'b1;
  assign \A[0][29] [0] = 1'b1;
  assign \A[0][31] [0] = 1'b1;
  assign \A[0][32] [4] = 1'b1;
  assign \A[0][32] [3] = 1'b1;
  assign \A[0][32] [2] = 1'b1;
  assign \A[0][32] [1] = 1'b1;
  assign \A[0][32] [0] = 1'b1;
  assign \A[0][33] [1] = 1'b1;
  assign \A[0][33] [0] = 1'b1;
  assign \A[0][34] [4] = 1'b1;
  assign \A[0][34] [3] = 1'b1;
  assign \A[0][34] [2] = 1'b1;
  assign \A[0][34] [1] = 1'b1;
  assign \A[0][35] [1] = 1'b1;
  assign \A[0][37] [4] = 1'b1;
  assign \A[0][37] [3] = 1'b1;
  assign \A[0][37] [2] = 1'b1;
  assign \A[0][37] [1] = 1'b1;
  assign \A[0][37] [0] = 1'b1;
  assign \A[0][39] [0] = 1'b1;
  assign \A[0][41] [4] = 1'b1;
  assign \A[0][41] [3] = 1'b1;
  assign \A[0][41] [2] = 1'b1;
  assign \A[0][41] [1] = 1'b1;
  assign \A[0][41] [0] = 1'b1;
  assign \A[0][42] [1] = 1'b1;
  assign \A[0][43] [4] = 1'b1;
  assign \A[0][43] [3] = 1'b1;
  assign \A[0][43] [2] = 1'b1;
  assign \A[0][43] [1] = 1'b1;
  assign \A[0][46] [1] = 1'b1;
  assign \A[0][47] [1] = 1'b1;
  assign \A[0][48] [4] = 1'b1;
  assign \A[0][48] [3] = 1'b1;
  assign \A[0][48] [2] = 1'b1;
  assign \A[0][48] [1] = 1'b1;
  assign \A[0][48] [0] = 1'b1;
  assign \A[0][49] [4] = 1'b1;
  assign \A[0][49] [3] = 1'b1;
  assign \A[0][49] [2] = 1'b1;
  assign \A[0][49] [0] = 1'b1;
  assign \A[0][56] [0] = 1'b1;
  assign \A[0][57] [4] = 1'b1;
  assign \A[0][57] [3] = 1'b1;
  assign \A[0][57] [2] = 1'b1;
  assign \A[0][57] [1] = 1'b1;
  assign \A[0][57] [0] = 1'b1;
  assign \A[0][58] [4] = 1'b1;
  assign \A[0][58] [3] = 1'b1;
  assign \A[0][58] [2] = 1'b1;
  assign \A[0][58] [1] = 1'b1;
  assign \A[0][58] [0] = 1'b1;
  assign \A[0][59] [0] = 1'b1;
  assign \A[0][60] [1] = 1'b1;
  assign \A[0][61] [1] = 1'b1;
  assign \A[0][63] [1] = 1'b1;
  assign \A[0][65] [4] = 1'b1;
  assign \A[0][65] [3] = 1'b1;
  assign \A[0][65] [2] = 1'b1;
  assign \A[0][65] [1] = 1'b1;
  assign \A[0][65] [0] = 1'b1;
  assign \A[0][66] [4] = 1'b1;
  assign \A[0][66] [3] = 1'b1;
  assign \A[0][66] [2] = 1'b1;
  assign \A[0][66] [1] = 1'b1;
  assign \A[0][66] [0] = 1'b1;
  assign \A[0][67] [4] = 1'b1;
  assign \A[0][67] [3] = 1'b1;
  assign \A[0][67] [2] = 1'b1;
  assign \A[0][67] [1] = 1'b1;
  assign \A[0][67] [0] = 1'b1;
  assign \A[0][68] [0] = 1'b1;
  assign \A[0][70] [4] = 1'b1;
  assign \A[0][70] [3] = 1'b1;
  assign \A[0][70] [2] = 1'b1;
  assign \A[0][70] [1] = 1'b1;
  assign \A[0][71] [1] = 1'b1;
  assign \A[0][72] [0] = 1'b1;
  assign \A[0][74] [4] = 1'b1;
  assign \A[0][74] [3] = 1'b1;
  assign \A[0][74] [2] = 1'b1;
  assign \A[0][74] [1] = 1'b1;
  assign \A[0][74] [0] = 1'b1;
  assign \A[0][75] [4] = 1'b1;
  assign \A[0][75] [3] = 1'b1;
  assign \A[0][75] [2] = 1'b1;
  assign \A[0][75] [0] = 1'b1;
  assign \A[0][76] [0] = 1'b1;
  assign \A[0][77] [4] = 1'b1;
  assign \A[0][77] [3] = 1'b1;
  assign \A[0][77] [2] = 1'b1;
  assign \A[0][77] [1] = 1'b1;
  assign \A[0][80] [4] = 1'b1;
  assign \A[0][80] [3] = 1'b1;
  assign \A[0][80] [2] = 1'b1;
  assign \A[0][80] [0] = 1'b1;
  assign \A[0][81] [4] = 1'b1;
  assign \A[0][81] [3] = 1'b1;
  assign \A[0][81] [2] = 1'b1;
  assign \A[0][81] [1] = 1'b1;
  assign \A[0][81] [0] = 1'b1;
  assign \A[0][82] [0] = 1'b1;
  assign \A[0][83] [1] = 1'b1;
  assign \A[0][84] [4] = 1'b1;
  assign \A[0][84] [3] = 1'b1;
  assign \A[0][84] [2] = 1'b1;
  assign \A[0][84] [1] = 1'b1;
  assign \A[0][85] [4] = 1'b1;
  assign \A[0][85] [3] = 1'b1;
  assign \A[0][85] [2] = 1'b1;
  assign \A[0][85] [1] = 1'b1;
  assign \A[0][85] [0] = 1'b1;
  assign \A[0][86] [4] = 1'b1;
  assign \A[0][86] [3] = 1'b1;
  assign \A[0][86] [2] = 1'b1;
  assign \A[0][86] [1] = 1'b1;
  assign \A[0][86] [0] = 1'b1;
  assign \A[0][88] [1] = 1'b1;
  assign \A[0][89] [4] = 1'b1;
  assign \A[0][89] [3] = 1'b1;
  assign \A[0][89] [2] = 1'b1;
  assign \A[0][89] [1] = 1'b1;
  assign \A[0][90] [4] = 1'b1;
  assign \A[0][90] [3] = 1'b1;
  assign \A[0][90] [2] = 1'b1;
  assign \A[0][90] [1] = 1'b1;
  assign \A[0][90] [0] = 1'b1;
  assign \A[0][92] [0] = 1'b1;
  assign \A[0][93] [0] = 1'b1;
  assign \A[0][94] [4] = 1'b1;
  assign \A[0][94] [3] = 1'b1;
  assign \A[0][94] [2] = 1'b1;
  assign \A[0][94] [1] = 1'b1;
  assign \A[0][95] [1] = 1'b1;
  assign \A[0][96] [4] = 1'b1;
  assign \A[0][96] [3] = 1'b1;
  assign \A[0][96] [2] = 1'b1;
  assign \A[0][96] [1] = 1'b1;
  assign \A[0][96] [0] = 1'b1;
  assign \A[0][97] [4] = 1'b1;
  assign \A[0][97] [3] = 1'b1;
  assign \A[0][97] [2] = 1'b1;
  assign \A[0][97] [1] = 1'b1;
  assign \A[0][97] [0] = 1'b1;
  assign \A[0][98] [4] = 1'b1;
  assign \A[0][98] [3] = 1'b1;
  assign \A[0][98] [2] = 1'b1;
  assign \A[0][98] [1] = 1'b1;
  assign \A[0][98] [0] = 1'b1;
  assign \A[0][100] [0] = 1'b1;
  assign \A[0][101] [4] = 1'b1;
  assign \A[0][101] [3] = 1'b1;
  assign \A[0][101] [2] = 1'b1;
  assign \A[0][101] [1] = 1'b1;
  assign \A[0][101] [0] = 1'b1;
  assign \A[0][102] [0] = 1'b1;
  assign \A[0][103] [1] = 1'b1;
  assign \A[0][104] [4] = 1'b1;
  assign \A[0][104] [3] = 1'b1;
  assign \A[0][104] [2] = 1'b1;
  assign \A[0][104] [0] = 1'b1;
  assign \A[0][105] [4] = 1'b1;
  assign \A[0][105] [3] = 1'b1;
  assign \A[0][105] [2] = 1'b1;
  assign \A[0][105] [1] = 1'b1;
  assign \A[0][105] [0] = 1'b1;
  assign \A[0][106] [4] = 1'b1;
  assign \A[0][106] [3] = 1'b1;
  assign \A[0][106] [2] = 1'b1;
  assign \A[0][106] [0] = 1'b1;
  assign \A[0][108] [4] = 1'b1;
  assign \A[0][108] [3] = 1'b1;
  assign \A[0][108] [2] = 1'b1;
  assign \A[0][108] [1] = 1'b1;
  assign \A[0][111] [0] = 1'b1;
  assign \A[0][112] [4] = 1'b1;
  assign \A[0][112] [3] = 1'b1;
  assign \A[0][112] [2] = 1'b1;
  assign \A[0][112] [1] = 1'b1;
  assign \A[0][112] [0] = 1'b1;
  assign \A[0][114] [1] = 1'b1;
  assign \A[0][115] [4] = 1'b1;
  assign \A[0][115] [3] = 1'b1;
  assign \A[0][115] [2] = 1'b1;
  assign \A[0][115] [1] = 1'b1;
  assign \A[0][117] [4] = 1'b1;
  assign \A[0][117] [3] = 1'b1;
  assign \A[0][117] [2] = 1'b1;
  assign \A[0][117] [1] = 1'b1;
  assign \A[0][118] [4] = 1'b1;
  assign \A[0][118] [3] = 1'b1;
  assign \A[0][118] [2] = 1'b1;
  assign \A[0][118] [1] = 1'b1;
  assign \A[0][119] [4] = 1'b1;
  assign \A[0][119] [3] = 1'b1;
  assign \A[0][119] [2] = 1'b1;
  assign \A[0][119] [0] = 1'b1;
  assign \A[0][120] [0] = 1'b1;
  assign \A[0][121] [4] = 1'b1;
  assign \A[0][121] [3] = 1'b1;
  assign \A[0][121] [2] = 1'b1;
  assign \A[0][121] [1] = 1'b1;
  assign \A[0][121] [0] = 1'b1;
  assign \A[0][122] [4] = 1'b1;
  assign \A[0][122] [3] = 1'b1;
  assign \A[0][122] [2] = 1'b1;
  assign \A[0][122] [1] = 1'b1;
  assign \A[0][122] [0] = 1'b1;
  assign \A[0][123] [4] = 1'b1;
  assign \A[0][123] [3] = 1'b1;
  assign \A[0][123] [2] = 1'b1;
  assign \A[0][123] [1] = 1'b1;
  assign \A[0][123] [0] = 1'b1;
  assign \A[0][125] [4] = 1'b1;
  assign \A[0][125] [3] = 1'b1;
  assign \A[0][125] [2] = 1'b1;
  assign \A[0][125] [1] = 1'b1;
  assign \A[0][125] [0] = 1'b1;
  assign \A[0][126] [4] = 1'b1;
  assign \A[0][126] [3] = 1'b1;
  assign \A[0][126] [2] = 1'b1;
  assign \A[0][126] [1] = 1'b1;
  assign \A[0][126] [0] = 1'b1;
  assign \A[0][128] [0] = 1'b1;
  assign \A[0][130] [0] = 1'b1;
  assign \A[0][132] [0] = 1'b1;
  assign \A[0][134] [4] = 1'b1;
  assign \A[0][134] [3] = 1'b1;
  assign \A[0][134] [2] = 1'b1;
  assign \A[0][134] [1] = 1'b1;
  assign \A[0][134] [0] = 1'b1;
  assign \A[0][136] [0] = 1'b1;
  assign \A[0][137] [4] = 1'b1;
  assign \A[0][137] [3] = 1'b1;
  assign \A[0][137] [2] = 1'b1;
  assign \A[0][138] [1] = 1'b1;
  assign \A[0][139] [0] = 1'b1;
  assign \A[0][141] [4] = 1'b1;
  assign \A[0][141] [3] = 1'b1;
  assign \A[0][141] [2] = 1'b1;
  assign \A[0][141] [1] = 1'b1;
  assign \A[0][141] [0] = 1'b1;
  assign \A[0][142] [4] = 1'b1;
  assign \A[0][142] [3] = 1'b1;
  assign \A[0][142] [2] = 1'b1;
  assign \A[0][142] [1] = 1'b1;
  assign \A[0][142] [0] = 1'b1;
  assign \A[0][144] [0] = 1'b1;
  assign \A[0][145] [4] = 1'b1;
  assign \A[0][145] [3] = 1'b1;
  assign \A[0][145] [2] = 1'b1;
  assign \A[0][145] [1] = 1'b1;
  assign \A[0][146] [1] = 1'b1;
  assign \A[0][146] [0] = 1'b1;
  assign \A[0][149] [4] = 1'b1;
  assign \A[0][149] [3] = 1'b1;
  assign \A[0][149] [2] = 1'b1;
  assign \A[0][149] [1] = 1'b1;
  assign \A[0][150] [0] = 1'b1;
  assign \A[0][151] [4] = 1'b1;
  assign \A[0][151] [3] = 1'b1;
  assign \A[0][151] [2] = 1'b1;
  assign \A[0][151] [1] = 1'b1;
  assign \A[0][153] [0] = 1'b1;
  assign \A[0][154] [4] = 1'b1;
  assign \A[0][154] [3] = 1'b1;
  assign \A[0][154] [2] = 1'b1;
  assign \A[0][154] [0] = 1'b1;
  assign \A[0][155] [4] = 1'b1;
  assign \A[0][155] [3] = 1'b1;
  assign \A[0][155] [2] = 1'b1;
  assign \A[0][155] [1] = 1'b1;
  assign \A[0][155] [0] = 1'b1;
  assign \A[0][156] [4] = 1'b1;
  assign \A[0][156] [3] = 1'b1;
  assign \A[0][156] [2] = 1'b1;
  assign \A[0][156] [1] = 1'b1;
  assign \A[0][156] [0] = 1'b1;
  assign \A[0][157] [4] = 1'b1;
  assign \A[0][157] [3] = 1'b1;
  assign \A[0][157] [2] = 1'b1;
  assign \A[0][157] [1] = 1'b1;
  assign \A[0][157] [0] = 1'b1;
  assign \A[0][158] [4] = 1'b1;
  assign \A[0][158] [3] = 1'b1;
  assign \A[0][158] [2] = 1'b1;
  assign \A[0][158] [1] = 1'b1;
  assign \A[0][158] [0] = 1'b1;
  assign \A[0][159] [1] = 1'b1;
  assign \A[0][162] [4] = 1'b1;
  assign \A[0][162] [3] = 1'b1;
  assign \A[0][162] [2] = 1'b1;
  assign \A[0][162] [1] = 1'b1;
  assign \A[0][164] [4] = 1'b1;
  assign \A[0][164] [3] = 1'b1;
  assign \A[0][164] [2] = 1'b1;
  assign \A[0][164] [1] = 1'b1;
  assign \A[0][165] [4] = 1'b1;
  assign \A[0][165] [3] = 1'b1;
  assign \A[0][165] [2] = 1'b1;
  assign \A[0][165] [1] = 1'b1;
  assign \A[0][165] [0] = 1'b1;
  assign \A[0][166] [0] = 1'b1;
  assign \A[0][167] [4] = 1'b1;
  assign \A[0][167] [3] = 1'b1;
  assign \A[0][167] [2] = 1'b1;
  assign \A[0][167] [0] = 1'b1;
  assign \A[0][169] [4] = 1'b1;
  assign \A[0][169] [3] = 1'b1;
  assign \A[0][169] [2] = 1'b1;
  assign \A[0][169] [1] = 1'b1;
  assign \A[0][169] [0] = 1'b1;
  assign \A[0][170] [4] = 1'b1;
  assign \A[0][170] [3] = 1'b1;
  assign \A[0][170] [2] = 1'b1;
  assign \A[0][170] [1] = 1'b1;
  assign \A[0][170] [0] = 1'b1;
  assign \A[0][171] [0] = 1'b1;
  assign \A[0][172] [4] = 1'b1;
  assign \A[0][172] [3] = 1'b1;
  assign \A[0][172] [2] = 1'b1;
  assign \A[0][172] [1] = 1'b1;
  assign \A[0][172] [0] = 1'b1;
  assign \A[0][174] [0] = 1'b1;
  assign \A[0][175] [4] = 1'b1;
  assign \A[0][175] [3] = 1'b1;
  assign \A[0][175] [2] = 1'b1;
  assign \A[0][175] [1] = 1'b1;
  assign \A[0][175] [0] = 1'b1;
  assign \A[0][176] [4] = 1'b1;
  assign \A[0][176] [3] = 1'b1;
  assign \A[0][176] [2] = 1'b1;
  assign \A[0][176] [1] = 1'b1;
  assign \A[0][176] [0] = 1'b1;
  assign \A[0][177] [4] = 1'b1;
  assign \A[0][177] [3] = 1'b1;
  assign \A[0][177] [2] = 1'b1;
  assign \A[0][177] [0] = 1'b1;
  assign \A[0][179] [0] = 1'b1;
  assign \A[0][183] [0] = 1'b1;
  assign \A[0][184] [4] = 1'b1;
  assign \A[0][184] [3] = 1'b1;
  assign \A[0][184] [2] = 1'b1;
  assign \A[0][184] [1] = 1'b1;
  assign \A[0][184] [0] = 1'b1;
  assign \A[0][185] [4] = 1'b1;
  assign \A[0][185] [3] = 1'b1;
  assign \A[0][185] [2] = 1'b1;
  assign \A[0][185] [1] = 1'b1;
  assign \A[0][186] [4] = 1'b1;
  assign \A[0][186] [3] = 1'b1;
  assign \A[0][186] [2] = 1'b1;
  assign \A[0][186] [1] = 1'b1;
  assign \A[0][187] [0] = 1'b1;
  assign \A[0][189] [0] = 1'b1;
  assign \A[0][190] [4] = 1'b1;
  assign \A[0][190] [3] = 1'b1;
  assign \A[0][190] [2] = 1'b1;
  assign \A[0][190] [1] = 1'b1;
  assign \A[0][190] [0] = 1'b1;
  assign \A[0][191] [1] = 1'b1;
  assign \A[0][193] [4] = 1'b1;
  assign \A[0][193] [3] = 1'b1;
  assign \A[0][193] [2] = 1'b1;
  assign \A[0][193] [1] = 1'b1;
  assign \A[0][194] [4] = 1'b1;
  assign \A[0][194] [3] = 1'b1;
  assign \A[0][194] [2] = 1'b1;
  assign \A[0][194] [1] = 1'b1;
  assign \A[0][195] [4] = 1'b1;
  assign \A[0][195] [3] = 1'b1;
  assign \A[0][195] [2] = 1'b1;
  assign \A[0][195] [1] = 1'b1;
  assign \A[0][195] [0] = 1'b1;
  assign \A[0][196] [0] = 1'b1;
  assign \A[0][197] [4] = 1'b1;
  assign \A[0][197] [3] = 1'b1;
  assign \A[0][197] [2] = 1'b1;
  assign \A[0][199] [4] = 1'b1;
  assign \A[0][199] [3] = 1'b1;
  assign \A[0][199] [2] = 1'b1;
  assign \A[0][199] [1] = 1'b1;
  assign \A[0][199] [0] = 1'b1;
  assign \A[0][200] [1] = 1'b1;
  assign \A[0][201] [0] = 1'b1;
  assign \A[0][202] [0] = 1'b1;
  assign \A[0][203] [0] = 1'b1;
  assign \A[0][204] [0] = 1'b1;
  assign \A[0][205] [4] = 1'b1;
  assign \A[0][205] [3] = 1'b1;
  assign \A[0][205] [2] = 1'b1;
  assign \A[0][205] [1] = 1'b1;
  assign \A[0][208] [4] = 1'b1;
  assign \A[0][208] [3] = 1'b1;
  assign \A[0][208] [2] = 1'b1;
  assign \A[0][208] [1] = 1'b1;
  assign \A[0][208] [0] = 1'b1;
  assign \A[0][209] [4] = 1'b1;
  assign \A[0][209] [3] = 1'b1;
  assign \A[0][209] [2] = 1'b1;
  assign \A[0][209] [1] = 1'b1;
  assign \A[0][210] [4] = 1'b1;
  assign \A[0][210] [3] = 1'b1;
  assign \A[0][210] [2] = 1'b1;
  assign \A[0][210] [1] = 1'b1;
  assign \A[0][210] [0] = 1'b1;
  assign \A[0][211] [4] = 1'b1;
  assign \A[0][211] [3] = 1'b1;
  assign \A[0][211] [2] = 1'b1;
  assign \A[0][211] [1] = 1'b1;
  assign \A[0][211] [0] = 1'b1;
  assign \A[0][212] [0] = 1'b1;
  assign \A[0][213] [4] = 1'b1;
  assign \A[0][213] [3] = 1'b1;
  assign \A[0][213] [2] = 1'b1;
  assign \A[0][213] [1] = 1'b1;
  assign \A[0][216] [1] = 1'b1;
  assign \A[0][216] [0] = 1'b1;
  assign \A[0][219] [0] = 1'b1;
  assign \A[0][220] [4] = 1'b1;
  assign \A[0][220] [3] = 1'b1;
  assign \A[0][220] [2] = 1'b1;
  assign \A[0][220] [1] = 1'b1;
  assign \A[0][220] [0] = 1'b1;
  assign \A[0][222] [0] = 1'b1;
  assign \A[0][224] [1] = 1'b1;
  assign \A[0][224] [0] = 1'b1;
  assign \A[0][226] [4] = 1'b1;
  assign \A[0][226] [3] = 1'b1;
  assign \A[0][226] [2] = 1'b1;
  assign \A[0][226] [1] = 1'b1;
  assign \A[0][226] [0] = 1'b1;
  assign \A[0][227] [0] = 1'b1;
  assign \A[0][228] [0] = 1'b1;
  assign \A[0][230] [4] = 1'b1;
  assign \A[0][230] [3] = 1'b1;
  assign \A[0][230] [2] = 1'b1;
  assign \A[0][230] [0] = 1'b1;
  assign \A[0][232] [4] = 1'b1;
  assign \A[0][232] [3] = 1'b1;
  assign \A[0][232] [2] = 1'b1;
  assign \A[0][232] [1] = 1'b1;
  assign \A[0][233] [0] = 1'b1;
  assign \A[0][234] [4] = 1'b1;
  assign \A[0][234] [3] = 1'b1;
  assign \A[0][234] [2] = 1'b1;
  assign \A[0][234] [1] = 1'b1;
  assign \A[0][235] [0] = 1'b1;
  assign \A[0][237] [1] = 1'b1;
  assign \A[0][238] [0] = 1'b1;
  assign \A[0][239] [1] = 1'b1;
  assign \A[0][241] [4] = 1'b1;
  assign \A[0][241] [3] = 1'b1;
  assign \A[0][241] [2] = 1'b1;
  assign \A[0][241] [1] = 1'b1;
  assign \A[0][241] [0] = 1'b1;
  assign \A[0][242] [4] = 1'b1;
  assign \A[0][242] [3] = 1'b1;
  assign \A[0][242] [2] = 1'b1;
  assign \A[0][242] [1] = 1'b1;
  assign \A[0][242] [0] = 1'b1;
  assign \A[0][243] [4] = 1'b1;
  assign \A[0][243] [3] = 1'b1;
  assign \A[0][243] [2] = 1'b1;
  assign \A[0][243] [1] = 1'b1;
  assign \A[0][243] [0] = 1'b1;
  assign \A[0][244] [1] = 1'b1;
  assign \A[0][245] [0] = 1'b1;
  assign \A[0][246] [1] = 1'b1;
  assign \A[0][247] [0] = 1'b1;
  assign \A[0][248] [1] = 1'b1;
  assign \A[0][248] [0] = 1'b1;
  assign \A[0][250] [4] = 1'b1;
  assign \A[0][250] [3] = 1'b1;
  assign \A[0][250] [2] = 1'b1;
  assign \A[0][250] [1] = 1'b1;
  assign \A[0][250] [0] = 1'b1;
  assign \A[0][252] [4] = 1'b1;
  assign \A[0][252] [3] = 1'b1;
  assign \A[0][252] [2] = 1'b1;
  assign \A[0][252] [1] = 1'b1;
  assign \A[0][253] [0] = 1'b1;
  assign \A[0][254] [4] = 1'b1;
  assign \A[0][254] [3] = 1'b1;
  assign \A[0][254] [2] = 1'b1;
  assign \A[0][254] [1] = 1'b1;
  assign \A[0][255] [4] = 1'b1;
  assign \A[0][255] [3] = 1'b1;
  assign \A[0][255] [2] = 1'b1;
  assign \A[0][255] [1] = 1'b1;
  assign \A[0][255] [0] = 1'b1;
  assign \A[1][0] [1] = 1'b1;
  assign \A[1][1] [4] = 1'b1;
  assign \A[1][1] [3] = 1'b1;
  assign \A[1][1] [2] = 1'b1;
  assign \A[1][1] [1] = 1'b1;
  assign \A[1][2] [4] = 1'b1;
  assign \A[1][2] [3] = 1'b1;
  assign \A[1][2] [2] = 1'b1;
  assign \A[1][2] [1] = 1'b1;
  assign \A[1][2] [0] = 1'b1;
  assign \A[1][5] [4] = 1'b1;
  assign \A[1][5] [3] = 1'b1;
  assign \A[1][5] [2] = 1'b1;
  assign \A[1][5] [1] = 1'b1;
  assign \A[1][6] [0] = 1'b1;
  assign \A[1][7] [4] = 1'b1;
  assign \A[1][7] [3] = 1'b1;
  assign \A[1][7] [2] = 1'b1;
  assign \A[1][7] [1] = 1'b1;
  assign \A[1][7] [0] = 1'b1;
  assign \A[1][8] [4] = 1'b1;
  assign \A[1][8] [3] = 1'b1;
  assign \A[1][8] [2] = 1'b1;
  assign \A[1][8] [1] = 1'b1;
  assign \A[1][8] [0] = 1'b1;
  assign \A[1][10] [4] = 1'b1;
  assign \A[1][10] [3] = 1'b1;
  assign \A[1][10] [2] = 1'b1;
  assign \A[1][10] [1] = 1'b1;
  assign \A[1][11] [1] = 1'b1;
  assign \A[1][12] [0] = 1'b1;
  assign \A[1][13] [4] = 1'b1;
  assign \A[1][13] [3] = 1'b1;
  assign \A[1][13] [2] = 1'b1;
  assign \A[1][13] [0] = 1'b1;
  assign \A[1][14] [0] = 1'b1;
  assign \A[1][16] [4] = 1'b1;
  assign \A[1][16] [3] = 1'b1;
  assign \A[1][16] [2] = 1'b1;
  assign \A[1][16] [1] = 1'b1;
  assign \A[1][16] [0] = 1'b1;
  assign \A[1][17] [4] = 1'b1;
  assign \A[1][17] [3] = 1'b1;
  assign \A[1][17] [2] = 1'b1;
  assign \A[1][17] [1] = 1'b1;
  assign \A[1][17] [0] = 1'b1;
  assign \A[1][19] [1] = 1'b1;
  assign \A[1][21] [4] = 1'b1;
  assign \A[1][21] [3] = 1'b1;
  assign \A[1][21] [2] = 1'b1;
  assign \A[1][21] [1] = 1'b1;
  assign \A[1][21] [0] = 1'b1;
  assign \A[1][23] [1] = 1'b1;
  assign \A[1][24] [4] = 1'b1;
  assign \A[1][24] [3] = 1'b1;
  assign \A[1][24] [2] = 1'b1;
  assign \A[1][24] [1] = 1'b1;
  assign \A[1][24] [0] = 1'b1;
  assign \A[1][26] [4] = 1'b1;
  assign \A[1][26] [3] = 1'b1;
  assign \A[1][26] [2] = 1'b1;
  assign \A[1][26] [0] = 1'b1;
  assign \A[1][28] [4] = 1'b1;
  assign \A[1][28] [3] = 1'b1;
  assign \A[1][28] [2] = 1'b1;
  assign \A[1][28] [1] = 1'b1;
  assign \A[1][28] [0] = 1'b1;
  assign \A[1][29] [4] = 1'b1;
  assign \A[1][29] [3] = 1'b1;
  assign \A[1][29] [2] = 1'b1;
  assign \A[1][29] [1] = 1'b1;
  assign \A[1][29] [0] = 1'b1;
  assign \A[1][30] [1] = 1'b1;
  assign \A[1][32] [4] = 1'b1;
  assign \A[1][32] [3] = 1'b1;
  assign \A[1][32] [2] = 1'b1;
  assign \A[1][32] [1] = 1'b1;
  assign \A[1][33] [4] = 1'b1;
  assign \A[1][33] [3] = 1'b1;
  assign \A[1][33] [2] = 1'b1;
  assign \A[1][33] [0] = 1'b1;
  assign \A[1][39] [4] = 1'b1;
  assign \A[1][39] [3] = 1'b1;
  assign \A[1][39] [2] = 1'b1;
  assign \A[1][39] [1] = 1'b1;
  assign \A[1][39] [0] = 1'b1;
  assign \A[1][40] [4] = 1'b1;
  assign \A[1][40] [3] = 1'b1;
  assign \A[1][40] [2] = 1'b1;
  assign \A[1][40] [1] = 1'b1;
  assign \A[1][41] [4] = 1'b1;
  assign \A[1][41] [3] = 1'b1;
  assign \A[1][41] [2] = 1'b1;
  assign \A[1][41] [1] = 1'b1;
  assign \A[1][41] [0] = 1'b1;
  assign \A[1][44] [4] = 1'b1;
  assign \A[1][44] [3] = 1'b1;
  assign \A[1][44] [2] = 1'b1;
  assign \A[1][44] [1] = 1'b1;
  assign \A[1][44] [0] = 1'b1;
  assign \A[1][45] [4] = 1'b1;
  assign \A[1][45] [3] = 1'b1;
  assign \A[1][45] [2] = 1'b1;
  assign \A[1][45] [1] = 1'b1;
  assign \A[1][45] [0] = 1'b1;
  assign \A[1][48] [4] = 1'b1;
  assign \A[1][48] [3] = 1'b1;
  assign \A[1][48] [2] = 1'b1;
  assign \A[1][48] [1] = 1'b1;
  assign \A[1][48] [0] = 1'b1;
  assign \A[1][49] [1] = 1'b1;
  assign \A[1][49] [0] = 1'b1;
  assign \A[1][50] [4] = 1'b1;
  assign \A[1][50] [3] = 1'b1;
  assign \A[1][50] [2] = 1'b1;
  assign \A[1][50] [1] = 1'b1;
  assign \A[1][50] [0] = 1'b1;
  assign \A[1][51] [4] = 1'b1;
  assign \A[1][51] [3] = 1'b1;
  assign \A[1][51] [2] = 1'b1;
  assign \A[1][51] [1] = 1'b1;
  assign \A[1][51] [0] = 1'b1;
  assign \A[1][52] [4] = 1'b1;
  assign \A[1][52] [3] = 1'b1;
  assign \A[1][52] [2] = 1'b1;
  assign \A[1][52] [0] = 1'b1;
  assign \A[1][54] [0] = 1'b1;
  assign \A[1][55] [4] = 1'b1;
  assign \A[1][55] [3] = 1'b1;
  assign \A[1][55] [2] = 1'b1;
  assign \A[1][55] [1] = 1'b1;
  assign \A[1][55] [0] = 1'b1;
  assign \A[1][56] [4] = 1'b1;
  assign \A[1][56] [3] = 1'b1;
  assign \A[1][56] [2] = 1'b1;
  assign \A[1][56] [1] = 1'b1;
  assign \A[1][58] [4] = 1'b1;
  assign \A[1][58] [3] = 1'b1;
  assign \A[1][58] [2] = 1'b1;
  assign \A[1][58] [1] = 1'b1;
  assign \A[1][58] [0] = 1'b1;
  assign \A[1][59] [4] = 1'b1;
  assign \A[1][59] [3] = 1'b1;
  assign \A[1][59] [2] = 1'b1;
  assign \A[1][59] [1] = 1'b1;
  assign \A[1][60] [4] = 1'b1;
  assign \A[1][60] [3] = 1'b1;
  assign \A[1][60] [2] = 1'b1;
  assign \A[1][60] [1] = 1'b1;
  assign \A[1][60] [0] = 1'b1;
  assign \A[1][61] [0] = 1'b1;
  assign \A[1][62] [4] = 1'b1;
  assign \A[1][62] [3] = 1'b1;
  assign \A[1][62] [2] = 1'b1;
  assign \A[1][62] [0] = 1'b1;
  assign \A[1][65] [0] = 1'b1;
  assign \A[1][66] [4] = 1'b1;
  assign \A[1][66] [3] = 1'b1;
  assign \A[1][66] [2] = 1'b1;
  assign \A[1][66] [1] = 1'b1;
  assign \A[1][67] [4] = 1'b1;
  assign \A[1][67] [3] = 1'b1;
  assign \A[1][67] [2] = 1'b1;
  assign \A[1][67] [1] = 1'b1;
  assign \A[1][68] [4] = 1'b1;
  assign \A[1][68] [3] = 1'b1;
  assign \A[1][68] [2] = 1'b1;
  assign \A[1][68] [0] = 1'b1;
  assign \A[1][69] [1] = 1'b1;
  assign \A[1][70] [0] = 1'b1;
  assign \A[1][71] [4] = 1'b1;
  assign \A[1][71] [3] = 1'b1;
  assign \A[1][71] [2] = 1'b1;
  assign \A[1][71] [1] = 1'b1;
  assign \A[1][73] [4] = 1'b1;
  assign \A[1][73] [3] = 1'b1;
  assign \A[1][73] [2] = 1'b1;
  assign \A[1][73] [1] = 1'b1;
  assign \A[1][73] [0] = 1'b1;
  assign \A[1][74] [4] = 1'b1;
  assign \A[1][74] [3] = 1'b1;
  assign \A[1][74] [2] = 1'b1;
  assign \A[1][74] [1] = 1'b1;
  assign \A[1][75] [0] = 1'b1;
  assign \A[1][76] [4] = 1'b1;
  assign \A[1][76] [3] = 1'b1;
  assign \A[1][76] [2] = 1'b1;
  assign \A[1][76] [1] = 1'b1;
  assign \A[1][77] [4] = 1'b1;
  assign \A[1][77] [3] = 1'b1;
  assign \A[1][77] [2] = 1'b1;
  assign \A[1][77] [1] = 1'b1;
  assign \A[1][77] [0] = 1'b1;
  assign \A[1][78] [4] = 1'b1;
  assign \A[1][78] [3] = 1'b1;
  assign \A[1][78] [2] = 1'b1;
  assign \A[1][78] [1] = 1'b1;
  assign \A[1][78] [0] = 1'b1;
  assign \A[1][79] [4] = 1'b1;
  assign \A[1][79] [3] = 1'b1;
  assign \A[1][79] [2] = 1'b1;
  assign \A[1][79] [0] = 1'b1;
  assign \A[1][81] [4] = 1'b1;
  assign \A[1][81] [3] = 1'b1;
  assign \A[1][81] [2] = 1'b1;
  assign \A[1][81] [0] = 1'b1;
  assign \A[1][82] [0] = 1'b1;
  assign \A[1][83] [4] = 1'b1;
  assign \A[1][83] [3] = 1'b1;
  assign \A[1][83] [2] = 1'b1;
  assign \A[1][83] [1] = 1'b1;
  assign \A[1][84] [4] = 1'b1;
  assign \A[1][84] [3] = 1'b1;
  assign \A[1][84] [2] = 1'b1;
  assign \A[1][84] [1] = 1'b1;
  assign \A[1][85] [0] = 1'b1;
  assign \A[1][88] [4] = 1'b1;
  assign \A[1][88] [3] = 1'b1;
  assign \A[1][88] [2] = 1'b1;
  assign \A[1][88] [1] = 1'b1;
  assign \A[1][88] [0] = 1'b1;
  assign \A[1][89] [4] = 1'b1;
  assign \A[1][89] [3] = 1'b1;
  assign \A[1][89] [2] = 1'b1;
  assign \A[1][89] [1] = 1'b1;
  assign \A[1][90] [0] = 1'b1;
  assign \A[1][91] [0] = 1'b1;
  assign \A[1][93] [0] = 1'b1;
  assign \A[1][94] [4] = 1'b1;
  assign \A[1][94] [3] = 1'b1;
  assign \A[1][94] [2] = 1'b1;
  assign \A[1][94] [1] = 1'b1;
  assign \A[1][94] [0] = 1'b1;
  assign \A[1][95] [1] = 1'b1;
  assign \A[1][96] [4] = 1'b1;
  assign \A[1][96] [3] = 1'b1;
  assign \A[1][96] [2] = 1'b1;
  assign \A[1][96] [1] = 1'b1;
  assign \A[1][96] [0] = 1'b1;
  assign \A[1][99] [0] = 1'b1;
  assign \A[1][100] [1] = 1'b1;
  assign \A[1][102] [1] = 1'b1;
  assign \A[1][103] [1] = 1'b1;
  assign \A[1][104] [1] = 1'b1;
  assign \A[1][104] [0] = 1'b1;
  assign \A[1][105] [4] = 1'b1;
  assign \A[1][105] [3] = 1'b1;
  assign \A[1][105] [2] = 1'b1;
  assign \A[1][105] [1] = 1'b1;
  assign \A[1][106] [0] = 1'b1;
  assign \A[1][107] [4] = 1'b1;
  assign \A[1][107] [3] = 1'b1;
  assign \A[1][107] [2] = 1'b1;
  assign \A[1][107] [1] = 1'b1;
  assign \A[1][108] [0] = 1'b1;
  assign \A[1][109] [4] = 1'b1;
  assign \A[1][109] [3] = 1'b1;
  assign \A[1][109] [2] = 1'b1;
  assign \A[1][109] [1] = 1'b1;
  assign \A[1][109] [0] = 1'b1;
  assign \A[1][110] [4] = 1'b1;
  assign \A[1][110] [3] = 1'b1;
  assign \A[1][110] [2] = 1'b1;
  assign \A[1][110] [1] = 1'b1;
  assign \A[1][110] [0] = 1'b1;
  assign \A[1][111] [4] = 1'b1;
  assign \A[1][111] [3] = 1'b1;
  assign \A[1][111] [2] = 1'b1;
  assign \A[1][111] [1] = 1'b1;
  assign \A[1][111] [0] = 1'b1;
  assign \A[1][112] [4] = 1'b1;
  assign \A[1][112] [3] = 1'b1;
  assign \A[1][112] [2] = 1'b1;
  assign \A[1][112] [1] = 1'b1;
  assign \A[1][112] [0] = 1'b1;
  assign \A[1][113] [4] = 1'b1;
  assign \A[1][113] [3] = 1'b1;
  assign \A[1][113] [2] = 1'b1;
  assign \A[1][113] [1] = 1'b1;
  assign \A[1][113] [0] = 1'b1;
  assign \A[1][114] [4] = 1'b1;
  assign \A[1][114] [3] = 1'b1;
  assign \A[1][114] [2] = 1'b1;
  assign \A[1][114] [1] = 1'b1;
  assign \A[1][115] [4] = 1'b1;
  assign \A[1][115] [3] = 1'b1;
  assign \A[1][115] [2] = 1'b1;
  assign \A[1][115] [1] = 1'b1;
  assign \A[1][115] [0] = 1'b1;
  assign \A[1][118] [0] = 1'b1;
  assign \A[1][119] [0] = 1'b1;
  assign \A[1][122] [0] = 1'b1;
  assign \A[1][123] [4] = 1'b1;
  assign \A[1][123] [3] = 1'b1;
  assign \A[1][123] [2] = 1'b1;
  assign \A[1][123] [1] = 1'b1;
  assign \A[1][130] [0] = 1'b1;
  assign \A[1][131] [0] = 1'b1;
  assign \A[1][132] [4] = 1'b1;
  assign \A[1][132] [3] = 1'b1;
  assign \A[1][132] [2] = 1'b1;
  assign \A[1][132] [1] = 1'b1;
  assign \A[1][133] [0] = 1'b1;
  assign \A[1][134] [4] = 1'b1;
  assign \A[1][134] [3] = 1'b1;
  assign \A[1][134] [2] = 1'b1;
  assign \A[1][134] [1] = 1'b1;
  assign \A[1][134] [0] = 1'b1;
  assign \A[1][135] [4] = 1'b1;
  assign \A[1][135] [3] = 1'b1;
  assign \A[1][135] [2] = 1'b1;
  assign \A[1][135] [1] = 1'b1;
  assign \A[1][135] [0] = 1'b1;
  assign \A[1][137] [4] = 1'b1;
  assign \A[1][137] [3] = 1'b1;
  assign \A[1][137] [2] = 1'b1;
  assign \A[1][137] [1] = 1'b1;
  assign \A[1][137] [0] = 1'b1;
  assign \A[1][138] [0] = 1'b1;
  assign \A[1][141] [1] = 1'b1;
  assign \A[1][143] [1] = 1'b1;
  assign \A[1][143] [0] = 1'b1;
  assign \A[1][145] [1] = 1'b1;
  assign \A[1][146] [1] = 1'b1;
  assign \A[1][146] [0] = 1'b1;
  assign \A[1][147] [4] = 1'b1;
  assign \A[1][147] [3] = 1'b1;
  assign \A[1][147] [2] = 1'b1;
  assign \A[1][147] [0] = 1'b1;
  assign \A[1][148] [4] = 1'b1;
  assign \A[1][148] [3] = 1'b1;
  assign \A[1][148] [2] = 1'b1;
  assign \A[1][148] [0] = 1'b1;
  assign \A[1][149] [4] = 1'b1;
  assign \A[1][149] [3] = 1'b1;
  assign \A[1][149] [2] = 1'b1;
  assign \A[1][149] [1] = 1'b1;
  assign \A[1][149] [0] = 1'b1;
  assign \A[1][151] [1] = 1'b1;
  assign \A[1][151] [0] = 1'b1;
  assign \A[1][152] [0] = 1'b1;
  assign \A[1][154] [1] = 1'b1;
  assign \A[1][155] [4] = 1'b1;
  assign \A[1][155] [3] = 1'b1;
  assign \A[1][155] [2] = 1'b1;
  assign \A[1][155] [1] = 1'b1;
  assign \A[1][156] [4] = 1'b1;
  assign \A[1][156] [3] = 1'b1;
  assign \A[1][156] [2] = 1'b1;
  assign \A[1][156] [1] = 1'b1;
  assign \A[1][156] [0] = 1'b1;
  assign \A[1][157] [0] = 1'b1;
  assign \A[1][158] [0] = 1'b1;
  assign \A[1][160] [1] = 1'b1;
  assign \A[1][161] [4] = 1'b1;
  assign \A[1][161] [3] = 1'b1;
  assign \A[1][161] [2] = 1'b1;
  assign \A[1][161] [1] = 1'b1;
  assign \A[1][161] [0] = 1'b1;
  assign \A[1][162] [4] = 1'b1;
  assign \A[1][162] [3] = 1'b1;
  assign \A[1][162] [2] = 1'b1;
  assign \A[1][162] [1] = 1'b1;
  assign \A[1][162] [0] = 1'b1;
  assign \A[1][164] [4] = 1'b1;
  assign \A[1][164] [3] = 1'b1;
  assign \A[1][164] [2] = 1'b1;
  assign \A[1][164] [1] = 1'b1;
  assign \A[1][164] [0] = 1'b1;
  assign \A[1][166] [1] = 1'b1;
  assign \A[1][167] [4] = 1'b1;
  assign \A[1][167] [3] = 1'b1;
  assign \A[1][167] [2] = 1'b1;
  assign \A[1][167] [1] = 1'b1;
  assign \A[1][169] [4] = 1'b1;
  assign \A[1][169] [3] = 1'b1;
  assign \A[1][169] [2] = 1'b1;
  assign \A[1][169] [1] = 1'b1;
  assign \A[1][170] [0] = 1'b1;
  assign \A[1][171] [4] = 1'b1;
  assign \A[1][171] [3] = 1'b1;
  assign \A[1][171] [2] = 1'b1;
  assign \A[1][171] [1] = 1'b1;
  assign \A[1][173] [0] = 1'b1;
  assign \A[1][174] [1] = 1'b1;
  assign \A[1][174] [0] = 1'b1;
  assign \A[1][176] [0] = 1'b1;
  assign \A[1][177] [4] = 1'b1;
  assign \A[1][177] [3] = 1'b1;
  assign \A[1][177] [2] = 1'b1;
  assign \A[1][177] [1] = 1'b1;
  assign \A[1][177] [0] = 1'b1;
  assign \A[1][178] [4] = 1'b1;
  assign \A[1][178] [3] = 1'b1;
  assign \A[1][178] [2] = 1'b1;
  assign \A[1][178] [1] = 1'b1;
  assign \A[1][178] [0] = 1'b1;
  assign \A[1][179] [4] = 1'b1;
  assign \A[1][179] [3] = 1'b1;
  assign \A[1][179] [2] = 1'b1;
  assign \A[1][179] [1] = 1'b1;
  assign \A[1][179] [0] = 1'b1;
  assign \A[1][182] [4] = 1'b1;
  assign \A[1][182] [3] = 1'b1;
  assign \A[1][182] [2] = 1'b1;
  assign \A[1][182] [1] = 1'b1;
  assign \A[1][183] [1] = 1'b1;
  assign \A[1][184] [4] = 1'b1;
  assign \A[1][184] [3] = 1'b1;
  assign \A[1][184] [2] = 1'b1;
  assign \A[1][184] [1] = 1'b1;
  assign \A[1][184] [0] = 1'b1;
  assign \A[1][185] [4] = 1'b1;
  assign \A[1][185] [3] = 1'b1;
  assign \A[1][185] [2] = 1'b1;
  assign \A[1][185] [1] = 1'b1;
  assign \A[1][185] [0] = 1'b1;
  assign \A[1][186] [4] = 1'b1;
  assign \A[1][186] [3] = 1'b1;
  assign \A[1][186] [2] = 1'b1;
  assign \A[1][186] [0] = 1'b1;
  assign \A[1][187] [1] = 1'b1;
  assign \A[1][187] [0] = 1'b1;
  assign \A[1][188] [1] = 1'b1;
  assign \A[1][189] [4] = 1'b1;
  assign \A[1][189] [3] = 1'b1;
  assign \A[1][189] [2] = 1'b1;
  assign \A[1][189] [0] = 1'b1;
  assign \A[1][190] [1] = 1'b1;
  assign \A[1][190] [0] = 1'b1;
  assign \A[1][191] [1] = 1'b1;
  assign \A[1][192] [1] = 1'b1;
  assign \A[1][192] [0] = 1'b1;
  assign \A[1][193] [4] = 1'b1;
  assign \A[1][193] [3] = 1'b1;
  assign \A[1][193] [2] = 1'b1;
  assign \A[1][193] [1] = 1'b1;
  assign \A[1][193] [0] = 1'b1;
  assign \A[1][194] [4] = 1'b1;
  assign \A[1][194] [3] = 1'b1;
  assign \A[1][194] [2] = 1'b1;
  assign \A[1][194] [1] = 1'b1;
  assign \A[1][194] [0] = 1'b1;
  assign \A[1][195] [1] = 1'b1;
  assign \A[1][195] [0] = 1'b1;
  assign \A[1][196] [1] = 1'b1;
  assign \A[1][196] [0] = 1'b1;
  assign \A[1][197] [4] = 1'b1;
  assign \A[1][197] [3] = 1'b1;
  assign \A[1][197] [2] = 1'b1;
  assign \A[1][197] [0] = 1'b1;
  assign \A[1][198] [0] = 1'b1;
  assign \A[1][199] [4] = 1'b1;
  assign \A[1][199] [3] = 1'b1;
  assign \A[1][199] [2] = 1'b1;
  assign \A[1][199] [1] = 1'b1;
  assign \A[1][199] [0] = 1'b1;
  assign \A[1][200] [0] = 1'b1;
  assign \A[1][202] [0] = 1'b1;
  assign \A[1][204] [4] = 1'b1;
  assign \A[1][204] [3] = 1'b1;
  assign \A[1][204] [2] = 1'b1;
  assign \A[1][204] [1] = 1'b1;
  assign \A[1][204] [0] = 1'b1;
  assign \A[1][207] [4] = 1'b1;
  assign \A[1][207] [3] = 1'b1;
  assign \A[1][207] [2] = 1'b1;
  assign \A[1][207] [1] = 1'b1;
  assign \A[1][207] [0] = 1'b1;
  assign \A[1][208] [4] = 1'b1;
  assign \A[1][208] [3] = 1'b1;
  assign \A[1][208] [2] = 1'b1;
  assign \A[1][208] [1] = 1'b1;
  assign \A[1][208] [0] = 1'b1;
  assign \A[1][209] [4] = 1'b1;
  assign \A[1][209] [3] = 1'b1;
  assign \A[1][209] [2] = 1'b1;
  assign \A[1][209] [1] = 1'b1;
  assign \A[1][209] [0] = 1'b1;
  assign \A[1][210] [4] = 1'b1;
  assign \A[1][210] [3] = 1'b1;
  assign \A[1][210] [2] = 1'b1;
  assign \A[1][210] [1] = 1'b1;
  assign \A[1][210] [0] = 1'b1;
  assign \A[1][211] [4] = 1'b1;
  assign \A[1][211] [3] = 1'b1;
  assign \A[1][211] [2] = 1'b1;
  assign \A[1][211] [1] = 1'b1;
  assign \A[1][211] [0] = 1'b1;
  assign \A[1][212] [0] = 1'b1;
  assign \A[1][214] [4] = 1'b1;
  assign \A[1][214] [3] = 1'b1;
  assign \A[1][214] [2] = 1'b1;
  assign \A[1][214] [1] = 1'b1;
  assign \A[1][216] [4] = 1'b1;
  assign \A[1][216] [3] = 1'b1;
  assign \A[1][216] [2] = 1'b1;
  assign \A[1][216] [1] = 1'b1;
  assign \A[1][216] [0] = 1'b1;
  assign \A[1][217] [4] = 1'b1;
  assign \A[1][217] [3] = 1'b1;
  assign \A[1][217] [2] = 1'b1;
  assign \A[1][217] [1] = 1'b1;
  assign \A[1][218] [0] = 1'b1;
  assign \A[1][219] [4] = 1'b1;
  assign \A[1][219] [3] = 1'b1;
  assign \A[1][219] [2] = 1'b1;
  assign \A[1][219] [1] = 1'b1;
  assign \A[1][219] [0] = 1'b1;
  assign \A[1][220] [4] = 1'b1;
  assign \A[1][220] [3] = 1'b1;
  assign \A[1][220] [2] = 1'b1;
  assign \A[1][220] [1] = 1'b1;
  assign \A[1][220] [0] = 1'b1;
  assign \A[1][221] [0] = 1'b1;
  assign \A[1][223] [0] = 1'b1;
  assign \A[1][224] [4] = 1'b1;
  assign \A[1][224] [3] = 1'b1;
  assign \A[1][224] [2] = 1'b1;
  assign \A[1][224] [0] = 1'b1;
  assign \A[1][225] [4] = 1'b1;
  assign \A[1][225] [3] = 1'b1;
  assign \A[1][225] [2] = 1'b1;
  assign \A[1][225] [1] = 1'b1;
  assign \A[1][227] [4] = 1'b1;
  assign \A[1][227] [3] = 1'b1;
  assign \A[1][227] [2] = 1'b1;
  assign \A[1][227] [1] = 1'b1;
  assign \A[1][227] [0] = 1'b1;
  assign \A[1][228] [2] = 1'b1;
  assign \A[1][230] [0] = 1'b1;
  assign \A[1][231] [4] = 1'b1;
  assign \A[1][231] [3] = 1'b1;
  assign \A[1][231] [2] = 1'b1;
  assign \A[1][231] [1] = 1'b1;
  assign \A[1][232] [1] = 1'b1;
  assign \A[1][233] [1] = 1'b1;
  assign \A[1][234] [0] = 1'b1;
  assign \A[1][236] [0] = 1'b1;
  assign \A[1][237] [4] = 1'b1;
  assign \A[1][237] [3] = 1'b1;
  assign \A[1][237] [2] = 1'b1;
  assign \A[1][237] [1] = 1'b1;
  assign \A[1][237] [0] = 1'b1;
  assign \A[1][238] [1] = 1'b1;
  assign \A[1][238] [0] = 1'b1;
  assign \A[1][239] [4] = 1'b1;
  assign \A[1][239] [3] = 1'b1;
  assign \A[1][239] [2] = 1'b1;
  assign \A[1][239] [1] = 1'b1;
  assign \A[1][240] [4] = 1'b1;
  assign \A[1][240] [3] = 1'b1;
  assign \A[1][240] [2] = 1'b1;
  assign \A[1][240] [1] = 1'b1;
  assign \A[1][240] [0] = 1'b1;
  assign \A[1][241] [4] = 1'b1;
  assign \A[1][241] [3] = 1'b1;
  assign \A[1][241] [2] = 1'b1;
  assign \A[1][241] [0] = 1'b1;
  assign \A[1][242] [4] = 1'b1;
  assign \A[1][242] [3] = 1'b1;
  assign \A[1][242] [2] = 1'b1;
  assign \A[1][242] [1] = 1'b1;
  assign \A[1][243] [4] = 1'b1;
  assign \A[1][243] [3] = 1'b1;
  assign \A[1][243] [2] = 1'b1;
  assign \A[1][243] [0] = 1'b1;
  assign \A[1][244] [4] = 1'b1;
  assign \A[1][244] [3] = 1'b1;
  assign \A[1][244] [2] = 1'b1;
  assign \A[1][244] [1] = 1'b1;
  assign \A[1][244] [0] = 1'b1;
  assign \A[1][245] [0] = 1'b1;
  assign \A[1][247] [4] = 1'b1;
  assign \A[1][247] [3] = 1'b1;
  assign \A[1][247] [2] = 1'b1;
  assign \A[1][247] [1] = 1'b1;
  assign \A[1][247] [0] = 1'b1;
  assign \A[1][248] [4] = 1'b1;
  assign \A[1][248] [3] = 1'b1;
  assign \A[1][248] [2] = 1'b1;
  assign \A[1][248] [1] = 1'b1;
  assign \A[1][248] [0] = 1'b1;
  assign \A[1][250] [4] = 1'b1;
  assign \A[1][250] [3] = 1'b1;
  assign \A[1][250] [2] = 1'b1;
  assign \A[1][250] [1] = 1'b1;
  assign \A[1][250] [0] = 1'b1;
  assign \A[1][251] [4] = 1'b1;
  assign \A[1][251] [3] = 1'b1;
  assign \A[1][251] [2] = 1'b1;
  assign \A[1][251] [1] = 1'b1;
  assign \A[1][251] [0] = 1'b1;
  assign \A[1][252] [4] = 1'b1;
  assign \A[1][252] [3] = 1'b1;
  assign \A[1][252] [2] = 1'b1;
  assign \A[1][252] [1] = 1'b1;
  assign \A[1][252] [0] = 1'b1;
  assign \A[1][253] [0] = 1'b1;
  assign \A[1][254] [4] = 1'b1;
  assign \A[1][254] [3] = 1'b1;
  assign \A[1][254] [2] = 1'b1;
  assign \A[1][254] [1] = 1'b1;
  assign \A[1][254] [0] = 1'b1;
  assign \A[1][255] [4] = 1'b1;
  assign \A[1][255] [3] = 1'b1;
  assign \A[1][255] [2] = 1'b1;
  assign \A[1][255] [1] = 1'b1;
  assign \A[2][0] [4] = 1'b1;
  assign \A[2][0] [3] = 1'b1;
  assign \A[2][0] [1] = 1'b1;
  assign \A[2][2] [4] = 1'b1;
  assign \A[2][2] [3] = 1'b1;
  assign \A[2][2] [2] = 1'b1;
  assign \A[2][2] [1] = 1'b1;
  assign \A[2][2] [0] = 1'b1;
  assign \A[2][4] [4] = 1'b1;
  assign \A[2][4] [3] = 1'b1;
  assign \A[2][4] [2] = 1'b1;
  assign \A[2][4] [1] = 1'b1;
  assign \A[2][4] [0] = 1'b1;
  assign \A[2][5] [4] = 1'b1;
  assign \A[2][5] [3] = 1'b1;
  assign \A[2][5] [2] = 1'b1;
  assign \A[2][5] [0] = 1'b1;
  assign \A[2][6] [4] = 1'b1;
  assign \A[2][6] [3] = 1'b1;
  assign \A[2][6] [2] = 1'b1;
  assign \A[2][6] [1] = 1'b1;
  assign \A[2][6] [0] = 1'b1;
  assign \A[2][7] [4] = 1'b1;
  assign \A[2][7] [3] = 1'b1;
  assign \A[2][7] [2] = 1'b1;
  assign \A[2][7] [0] = 1'b1;
  assign \A[2][8] [0] = 1'b1;
  assign \A[2][9] [4] = 1'b1;
  assign \A[2][9] [3] = 1'b1;
  assign \A[2][9] [2] = 1'b1;
  assign \A[2][9] [1] = 1'b1;
  assign \A[2][10] [4] = 1'b1;
  assign \A[2][10] [3] = 1'b1;
  assign \A[2][10] [2] = 1'b1;
  assign \A[2][10] [1] = 1'b1;
  assign \A[2][11] [4] = 1'b1;
  assign \A[2][11] [3] = 1'b1;
  assign \A[2][11] [2] = 1'b1;
  assign \A[2][11] [1] = 1'b1;
  assign \A[2][12] [4] = 1'b1;
  assign \A[2][12] [3] = 1'b1;
  assign \A[2][12] [2] = 1'b1;
  assign \A[2][12] [1] = 1'b1;
  assign \A[2][12] [0] = 1'b1;
  assign \A[2][13] [4] = 1'b1;
  assign \A[2][13] [3] = 1'b1;
  assign \A[2][13] [1] = 1'b1;
  assign \A[2][13] [0] = 1'b1;
  assign \A[2][14] [4] = 1'b1;
  assign \A[2][14] [3] = 1'b1;
  assign \A[2][14] [2] = 1'b1;
  assign \A[2][14] [1] = 1'b1;
  assign \A[2][14] [0] = 1'b1;
  assign \A[2][15] [4] = 1'b1;
  assign \A[2][15] [3] = 1'b1;
  assign \A[2][15] [2] = 1'b1;
  assign \A[2][15] [1] = 1'b1;
  assign \A[2][15] [0] = 1'b1;
  assign \A[2][16] [4] = 1'b1;
  assign \A[2][16] [3] = 1'b1;
  assign \A[2][16] [2] = 1'b1;
  assign \A[2][16] [1] = 1'b1;
  assign \A[2][16] [0] = 1'b1;
  assign \A[2][17] [4] = 1'b1;
  assign \A[2][17] [3] = 1'b1;
  assign \A[2][17] [2] = 1'b1;
  assign \A[2][17] [1] = 1'b1;
  assign \A[2][17] [0] = 1'b1;
  assign \A[2][18] [4] = 1'b1;
  assign \A[2][18] [3] = 1'b1;
  assign \A[2][18] [2] = 1'b1;
  assign \A[2][18] [1] = 1'b1;
  assign \A[2][19] [4] = 1'b1;
  assign \A[2][19] [3] = 1'b1;
  assign \A[2][19] [2] = 1'b1;
  assign \A[2][19] [1] = 1'b1;
  assign \A[2][19] [0] = 1'b1;
  assign \A[2][20] [4] = 1'b1;
  assign \A[2][20] [3] = 1'b1;
  assign \A[2][20] [2] = 1'b1;
  assign \A[2][20] [0] = 1'b1;
  assign \A[2][21] [1] = 1'b1;
  assign \A[2][22] [4] = 1'b1;
  assign \A[2][22] [3] = 1'b1;
  assign \A[2][22] [2] = 1'b1;
  assign \A[2][22] [1] = 1'b1;
  assign \A[2][25] [4] = 1'b1;
  assign \A[2][25] [3] = 1'b1;
  assign \A[2][25] [2] = 1'b1;
  assign \A[2][25] [1] = 1'b1;
  assign \A[2][27] [4] = 1'b1;
  assign \A[2][27] [3] = 1'b1;
  assign \A[2][27] [2] = 1'b1;
  assign \A[2][27] [1] = 1'b1;
  assign \A[2][29] [1] = 1'b1;
  assign \A[2][30] [4] = 1'b1;
  assign \A[2][30] [3] = 1'b1;
  assign \A[2][30] [2] = 1'b1;
  assign \A[2][30] [1] = 1'b1;
  assign \A[2][30] [0] = 1'b1;
  assign \A[2][31] [4] = 1'b1;
  assign \A[2][31] [3] = 1'b1;
  assign \A[2][31] [2] = 1'b1;
  assign \A[2][31] [1] = 1'b1;
  assign \A[2][32] [4] = 1'b1;
  assign \A[2][32] [3] = 1'b1;
  assign \A[2][32] [2] = 1'b1;
  assign \A[2][33] [4] = 1'b1;
  assign \A[2][33] [3] = 1'b1;
  assign \A[2][33] [2] = 1'b1;
  assign \A[2][33] [1] = 1'b1;
  assign \A[2][33] [0] = 1'b1;
  assign \A[2][34] [4] = 1'b1;
  assign \A[2][34] [3] = 1'b1;
  assign \A[2][34] [2] = 1'b1;
  assign \A[2][34] [1] = 1'b1;
  assign \A[2][34] [0] = 1'b1;
  assign \A[2][35] [4] = 1'b1;
  assign \A[2][35] [3] = 1'b1;
  assign \A[2][35] [2] = 1'b1;
  assign \A[2][35] [1] = 1'b1;
  assign \A[2][35] [0] = 1'b1;
  assign \A[2][37] [4] = 1'b1;
  assign \A[2][37] [3] = 1'b1;
  assign \A[2][37] [2] = 1'b1;
  assign \A[2][37] [1] = 1'b1;
  assign \A[2][39] [4] = 1'b1;
  assign \A[2][39] [3] = 1'b1;
  assign \A[2][39] [2] = 1'b1;
  assign \A[2][39] [1] = 1'b1;
  assign \A[2][39] [0] = 1'b1;
  assign \A[2][40] [4] = 1'b1;
  assign \A[2][40] [3] = 1'b1;
  assign \A[2][40] [2] = 1'b1;
  assign \A[2][40] [1] = 1'b1;
  assign \A[2][40] [0] = 1'b1;
  assign \A[2][42] [0] = 1'b1;
  assign \A[2][43] [4] = 1'b1;
  assign \A[2][43] [3] = 1'b1;
  assign \A[2][43] [2] = 1'b1;
  assign \A[2][43] [1] = 1'b1;
  assign \A[2][43] [0] = 1'b1;
  assign \A[2][44] [4] = 1'b1;
  assign \A[2][44] [3] = 1'b1;
  assign \A[2][44] [2] = 1'b1;
  assign \A[2][44] [1] = 1'b1;
  assign \A[2][45] [4] = 1'b1;
  assign \A[2][45] [3] = 1'b1;
  assign \A[2][45] [2] = 1'b1;
  assign \A[2][45] [0] = 1'b1;
  assign \A[2][46] [4] = 1'b1;
  assign \A[2][46] [3] = 1'b1;
  assign \A[2][46] [2] = 1'b1;
  assign \A[2][46] [1] = 1'b1;
  assign \A[2][46] [0] = 1'b1;
  assign \A[2][48] [0] = 1'b1;
  assign \A[2][50] [0] = 1'b1;
  assign \A[2][51] [4] = 1'b1;
  assign \A[2][51] [3] = 1'b1;
  assign \A[2][51] [2] = 1'b1;
  assign \A[2][51] [1] = 1'b1;
  assign \A[2][51] [0] = 1'b1;
  assign \A[2][52] [4] = 1'b1;
  assign \A[2][52] [3] = 1'b1;
  assign \A[2][52] [2] = 1'b1;
  assign \A[2][52] [1] = 1'b1;
  assign \A[2][52] [0] = 1'b1;
  assign \A[2][54] [0] = 1'b1;
  assign \A[2][55] [0] = 1'b1;
  assign \A[2][57] [0] = 1'b1;
  assign \A[2][58] [4] = 1'b1;
  assign \A[2][58] [3] = 1'b1;
  assign \A[2][58] [2] = 1'b1;
  assign \A[2][58] [1] = 1'b1;
  assign \A[2][58] [0] = 1'b1;
  assign \A[2][59] [1] = 1'b1;
  assign \A[2][60] [0] = 1'b1;
  assign \A[2][61] [4] = 1'b1;
  assign \A[2][61] [3] = 1'b1;
  assign \A[2][61] [2] = 1'b1;
  assign \A[2][61] [1] = 1'b1;
  assign \A[2][61] [0] = 1'b1;
  assign \A[2][62] [4] = 1'b1;
  assign \A[2][62] [3] = 1'b1;
  assign \A[2][62] [2] = 1'b1;
  assign \A[2][62] [1] = 1'b1;
  assign \A[2][62] [0] = 1'b1;
  assign \A[2][63] [0] = 1'b1;
  assign \A[2][64] [4] = 1'b1;
  assign \A[2][64] [3] = 1'b1;
  assign \A[2][64] [2] = 1'b1;
  assign \A[2][64] [1] = 1'b1;
  assign \A[2][64] [0] = 1'b1;
  assign \A[2][66] [1] = 1'b1;
  assign \A[2][67] [0] = 1'b1;
  assign \A[2][69] [4] = 1'b1;
  assign \A[2][69] [3] = 1'b1;
  assign \A[2][69] [2] = 1'b1;
  assign \A[2][69] [1] = 1'b1;
  assign \A[2][69] [0] = 1'b1;
  assign \A[2][70] [4] = 1'b1;
  assign \A[2][70] [3] = 1'b1;
  assign \A[2][70] [2] = 1'b1;
  assign \A[2][70] [1] = 1'b1;
  assign \A[2][70] [0] = 1'b1;
  assign \A[2][71] [1] = 1'b1;
  assign \A[2][72] [0] = 1'b1;
  assign \A[2][73] [0] = 1'b1;
  assign \A[2][74] [4] = 1'b1;
  assign \A[2][74] [3] = 1'b1;
  assign \A[2][74] [2] = 1'b1;
  assign \A[2][74] [1] = 1'b1;
  assign \A[2][74] [0] = 1'b1;
  assign \A[2][78] [4] = 1'b1;
  assign \A[2][78] [3] = 1'b1;
  assign \A[2][78] [2] = 1'b1;
  assign \A[2][78] [1] = 1'b1;
  assign \A[2][78] [0] = 1'b1;
  assign \A[2][79] [4] = 1'b1;
  assign \A[2][79] [3] = 1'b1;
  assign \A[2][79] [2] = 1'b1;
  assign \A[2][79] [0] = 1'b1;
  assign \A[2][80] [4] = 1'b1;
  assign \A[2][80] [3] = 1'b1;
  assign \A[2][80] [2] = 1'b1;
  assign \A[2][80] [1] = 1'b1;
  assign \A[2][80] [0] = 1'b1;
  assign \A[2][81] [4] = 1'b1;
  assign \A[2][81] [3] = 1'b1;
  assign \A[2][81] [2] = 1'b1;
  assign \A[2][81] [1] = 1'b1;
  assign \A[2][82] [0] = 1'b1;
  assign \A[2][83] [4] = 1'b1;
  assign \A[2][83] [3] = 1'b1;
  assign \A[2][83] [2] = 1'b1;
  assign \A[2][84] [1] = 1'b1;
  assign \A[2][85] [4] = 1'b1;
  assign \A[2][85] [3] = 1'b1;
  assign \A[2][85] [2] = 1'b1;
  assign \A[2][85] [1] = 1'b1;
  assign \A[2][85] [0] = 1'b1;
  assign \A[2][88] [1] = 1'b1;
  assign \A[2][88] [0] = 1'b1;
  assign \A[2][90] [1] = 1'b1;
  assign \A[2][90] [0] = 1'b1;
  assign \A[2][91] [4] = 1'b1;
  assign \A[2][91] [3] = 1'b1;
  assign \A[2][91] [2] = 1'b1;
  assign \A[2][91] [1] = 1'b1;
  assign \A[2][93] [0] = 1'b1;
  assign \A[2][94] [4] = 1'b1;
  assign \A[2][94] [3] = 1'b1;
  assign \A[2][94] [2] = 1'b1;
  assign \A[2][94] [1] = 1'b1;
  assign \A[2][95] [4] = 1'b1;
  assign \A[2][95] [3] = 1'b1;
  assign \A[2][95] [2] = 1'b1;
  assign \A[2][95] [1] = 1'b1;
  assign \A[2][95] [0] = 1'b1;
  assign \A[2][96] [4] = 1'b1;
  assign \A[2][96] [3] = 1'b1;
  assign \A[2][96] [2] = 1'b1;
  assign \A[2][96] [1] = 1'b1;
  assign \A[2][97] [1] = 1'b1;
  assign \A[2][97] [0] = 1'b1;
  assign \A[2][98] [4] = 1'b1;
  assign \A[2][98] [3] = 1'b1;
  assign \A[2][98] [2] = 1'b1;
  assign \A[2][98] [1] = 1'b1;
  assign \A[2][99] [0] = 1'b1;
  assign \A[2][100] [0] = 1'b1;
  assign \A[2][101] [4] = 1'b1;
  assign \A[2][101] [3] = 1'b1;
  assign \A[2][101] [2] = 1'b1;
  assign \A[2][101] [1] = 1'b1;
  assign \A[2][102] [4] = 1'b1;
  assign \A[2][102] [3] = 1'b1;
  assign \A[2][102] [2] = 1'b1;
  assign \A[2][102] [1] = 1'b1;
  assign \A[2][102] [0] = 1'b1;
  assign \A[2][104] [1] = 1'b1;
  assign \A[2][105] [4] = 1'b1;
  assign \A[2][105] [3] = 1'b1;
  assign \A[2][105] [2] = 1'b1;
  assign \A[2][105] [1] = 1'b1;
  assign \A[2][105] [0] = 1'b1;
  assign \A[2][106] [0] = 1'b1;
  assign \A[2][108] [0] = 1'b1;
  assign \A[2][109] [4] = 1'b1;
  assign \A[2][109] [3] = 1'b1;
  assign \A[2][109] [2] = 1'b1;
  assign \A[2][109] [1] = 1'b1;
  assign \A[2][109] [0] = 1'b1;
  assign \A[2][110] [1] = 1'b1;
  assign \A[2][110] [0] = 1'b1;
  assign \A[2][112] [1] = 1'b1;
  assign \A[2][112] [0] = 1'b1;
  assign \A[2][113] [4] = 1'b1;
  assign \A[2][113] [3] = 1'b1;
  assign \A[2][113] [2] = 1'b1;
  assign \A[2][113] [1] = 1'b1;
  assign \A[2][114] [1] = 1'b1;
  assign \A[2][115] [4] = 1'b1;
  assign \A[2][115] [3] = 1'b1;
  assign \A[2][115] [2] = 1'b1;
  assign \A[2][115] [1] = 1'b1;
  assign \A[2][115] [0] = 1'b1;
  assign \A[2][116] [0] = 1'b1;
  assign \A[2][117] [0] = 1'b1;
  assign \A[2][118] [4] = 1'b1;
  assign \A[2][118] [3] = 1'b1;
  assign \A[2][118] [2] = 1'b1;
  assign \A[2][118] [1] = 1'b1;
  assign \A[2][119] [1] = 1'b1;
  assign \A[2][121] [1] = 1'b1;
  assign \A[2][122] [0] = 1'b1;
  assign \A[2][124] [0] = 1'b1;
  assign \A[2][125] [0] = 1'b1;
  assign \A[2][127] [4] = 1'b1;
  assign \A[2][127] [3] = 1'b1;
  assign \A[2][127] [2] = 1'b1;
  assign \A[2][127] [1] = 1'b1;
  assign \A[2][127] [0] = 1'b1;
  assign \A[2][128] [4] = 1'b1;
  assign \A[2][128] [3] = 1'b1;
  assign \A[2][128] [2] = 1'b1;
  assign \A[2][128] [1] = 1'b1;
  assign \A[2][128] [0] = 1'b1;
  assign \A[2][129] [1] = 1'b1;
  assign \A[2][129] [0] = 1'b1;
  assign \A[2][130] [0] = 1'b1;
  assign \A[2][131] [1] = 1'b1;
  assign \A[2][132] [0] = 1'b1;
  assign \A[2][134] [4] = 1'b1;
  assign \A[2][134] [3] = 1'b1;
  assign \A[2][134] [2] = 1'b1;
  assign \A[2][134] [1] = 1'b1;
  assign \A[2][136] [4] = 1'b1;
  assign \A[2][136] [3] = 1'b1;
  assign \A[2][136] [2] = 1'b1;
  assign \A[2][136] [1] = 1'b1;
  assign \A[2][136] [0] = 1'b1;
  assign \A[2][137] [2] = 1'b1;
  assign \A[2][138] [0] = 1'b1;
  assign \A[2][140] [4] = 1'b1;
  assign \A[2][140] [3] = 1'b1;
  assign \A[2][140] [2] = 1'b1;
  assign \A[2][140] [1] = 1'b1;
  assign \A[2][141] [0] = 1'b1;
  assign \A[2][143] [4] = 1'b1;
  assign \A[2][143] [3] = 1'b1;
  assign \A[2][143] [2] = 1'b1;
  assign \A[2][143] [1] = 1'b1;
  assign \A[2][143] [0] = 1'b1;
  assign \A[2][144] [4] = 1'b1;
  assign \A[2][144] [3] = 1'b1;
  assign \A[2][144] [2] = 1'b1;
  assign \A[2][144] [0] = 1'b1;
  assign \A[2][145] [1] = 1'b1;
  assign \A[2][145] [0] = 1'b1;
  assign \A[2][146] [4] = 1'b1;
  assign \A[2][146] [3] = 1'b1;
  assign \A[2][146] [2] = 1'b1;
  assign \A[2][146] [0] = 1'b1;
  assign \A[2][147] [4] = 1'b1;
  assign \A[2][147] [3] = 1'b1;
  assign \A[2][147] [2] = 1'b1;
  assign \A[2][147] [1] = 1'b1;
  assign \A[2][147] [0] = 1'b1;
  assign \A[2][148] [1] = 1'b1;
  assign \A[2][149] [0] = 1'b1;
  assign \A[2][153] [4] = 1'b1;
  assign \A[2][153] [3] = 1'b1;
  assign \A[2][153] [2] = 1'b1;
  assign \A[2][153] [1] = 1'b1;
  assign \A[2][153] [0] = 1'b1;
  assign \A[2][154] [0] = 1'b1;
  assign \A[2][155] [1] = 1'b1;
  assign \A[2][156] [0] = 1'b1;
  assign \A[2][158] [1] = 1'b1;
  assign \A[2][159] [4] = 1'b1;
  assign \A[2][159] [3] = 1'b1;
  assign \A[2][159] [2] = 1'b1;
  assign \A[2][159] [0] = 1'b1;
  assign \A[2][161] [2] = 1'b1;
  assign \A[2][163] [0] = 1'b1;
  assign \A[2][164] [4] = 1'b1;
  assign \A[2][164] [3] = 1'b1;
  assign \A[2][164] [2] = 1'b1;
  assign \A[2][164] [1] = 1'b1;
  assign \A[2][164] [0] = 1'b1;
  assign \A[2][165] [0] = 1'b1;
  assign \A[2][166] [0] = 1'b1;
  assign \A[2][167] [1] = 1'b1;
  assign \A[2][167] [0] = 1'b1;
  assign \A[2][168] [1] = 1'b1;
  assign \A[2][169] [1] = 1'b1;
  assign \A[2][169] [0] = 1'b1;
  assign \A[2][171] [0] = 1'b1;
  assign \A[2][172] [1] = 1'b1;
  assign \A[2][173] [4] = 1'b1;
  assign \A[2][173] [3] = 1'b1;
  assign \A[2][173] [2] = 1'b1;
  assign \A[2][173] [1] = 1'b1;
  assign \A[2][173] [0] = 1'b1;
  assign \A[2][174] [4] = 1'b1;
  assign \A[2][174] [3] = 1'b1;
  assign \A[2][174] [2] = 1'b1;
  assign \A[2][174] [1] = 1'b1;
  assign \A[2][175] [0] = 1'b1;
  assign \A[2][176] [4] = 1'b1;
  assign \A[2][176] [3] = 1'b1;
  assign \A[2][176] [2] = 1'b1;
  assign \A[2][176] [1] = 1'b1;
  assign \A[2][176] [0] = 1'b1;
  assign \A[2][177] [4] = 1'b1;
  assign \A[2][177] [3] = 1'b1;
  assign \A[2][177] [2] = 1'b1;
  assign \A[2][177] [1] = 1'b1;
  assign \A[2][178] [4] = 1'b1;
  assign \A[2][178] [3] = 1'b1;
  assign \A[2][178] [2] = 1'b1;
  assign \A[2][178] [1] = 1'b1;
  assign \A[2][178] [0] = 1'b1;
  assign \A[2][179] [4] = 1'b1;
  assign \A[2][179] [3] = 1'b1;
  assign \A[2][179] [2] = 1'b1;
  assign \A[2][179] [1] = 1'b1;
  assign \A[2][179] [0] = 1'b1;
  assign \A[2][180] [4] = 1'b1;
  assign \A[2][180] [3] = 1'b1;
  assign \A[2][180] [2] = 1'b1;
  assign \A[2][180] [1] = 1'b1;
  assign \A[2][181] [1] = 1'b1;
  assign \A[2][181] [0] = 1'b1;
  assign \A[2][182] [0] = 1'b1;
  assign \A[2][183] [0] = 1'b1;
  assign \A[2][186] [0] = 1'b1;
  assign \A[2][187] [0] = 1'b1;
  assign \A[2][188] [0] = 1'b1;
  assign \A[2][189] [4] = 1'b1;
  assign \A[2][189] [3] = 1'b1;
  assign \A[2][189] [2] = 1'b1;
  assign \A[2][189] [1] = 1'b1;
  assign \A[2][189] [0] = 1'b1;
  assign \A[2][190] [4] = 1'b1;
  assign \A[2][190] [3] = 1'b1;
  assign \A[2][190] [2] = 1'b1;
  assign \A[2][190] [1] = 1'b1;
  assign \A[2][190] [0] = 1'b1;
  assign \A[2][191] [0] = 1'b1;
  assign \A[2][192] [1] = 1'b1;
  assign \A[2][193] [4] = 1'b1;
  assign \A[2][193] [3] = 1'b1;
  assign \A[2][193] [2] = 1'b1;
  assign \A[2][193] [1] = 1'b1;
  assign \A[2][193] [0] = 1'b1;
  assign \A[2][194] [1] = 1'b1;
  assign \A[2][195] [1] = 1'b1;
  assign \A[2][196] [0] = 1'b1;
  assign \A[2][197] [0] = 1'b1;
  assign \A[2][200] [4] = 1'b1;
  assign \A[2][200] [3] = 1'b1;
  assign \A[2][200] [2] = 1'b1;
  assign \A[2][200] [1] = 1'b1;
  assign \A[2][201] [1] = 1'b1;
  assign \A[2][201] [0] = 1'b1;
  assign \A[2][203] [1] = 1'b1;
  assign \A[2][203] [0] = 1'b1;
  assign \A[2][204] [0] = 1'b1;
  assign \A[2][205] [0] = 1'b1;
  assign \A[2][206] [0] = 1'b1;
  assign \A[2][207] [4] = 1'b1;
  assign \A[2][207] [3] = 1'b1;
  assign \A[2][207] [2] = 1'b1;
  assign \A[2][207] [1] = 1'b1;
  assign \A[2][207] [0] = 1'b1;
  assign \A[2][209] [0] = 1'b1;
  assign \A[2][210] [4] = 1'b1;
  assign \A[2][210] [3] = 1'b1;
  assign \A[2][210] [2] = 1'b1;
  assign \A[2][210] [1] = 1'b1;
  assign \A[2][211] [1] = 1'b1;
  assign \A[2][213] [4] = 1'b1;
  assign \A[2][213] [3] = 1'b1;
  assign \A[2][213] [2] = 1'b1;
  assign \A[2][213] [1] = 1'b1;
  assign \A[2][213] [0] = 1'b1;
  assign \A[2][214] [4] = 1'b1;
  assign \A[2][214] [3] = 1'b1;
  assign \A[2][214] [2] = 1'b1;
  assign \A[2][214] [0] = 1'b1;
  assign \A[2][215] [4] = 1'b1;
  assign \A[2][215] [3] = 1'b1;
  assign \A[2][215] [2] = 1'b1;
  assign \A[2][215] [1] = 1'b1;
  assign \A[2][216] [4] = 1'b1;
  assign \A[2][216] [3] = 1'b1;
  assign \A[2][216] [2] = 1'b1;
  assign \A[2][216] [1] = 1'b1;
  assign \A[2][216] [0] = 1'b1;
  assign \A[2][217] [4] = 1'b1;
  assign \A[2][217] [3] = 1'b1;
  assign \A[2][217] [2] = 1'b1;
  assign \A[2][217] [1] = 1'b1;
  assign \A[2][218] [4] = 1'b1;
  assign \A[2][218] [3] = 1'b1;
  assign \A[2][218] [2] = 1'b1;
  assign \A[2][218] [1] = 1'b1;
  assign \A[2][218] [0] = 1'b1;
  assign \A[2][219] [4] = 1'b1;
  assign \A[2][219] [3] = 1'b1;
  assign \A[2][219] [2] = 1'b1;
  assign \A[2][219] [1] = 1'b1;
  assign \A[2][220] [1] = 1'b1;
  assign \A[2][220] [0] = 1'b1;
  assign \A[2][221] [0] = 1'b1;
  assign \A[2][222] [4] = 1'b1;
  assign \A[2][222] [3] = 1'b1;
  assign \A[2][222] [2] = 1'b1;
  assign \A[2][222] [1] = 1'b1;
  assign \A[2][222] [0] = 1'b1;
  assign \A[2][224] [4] = 1'b1;
  assign \A[2][224] [3] = 1'b1;
  assign \A[2][224] [2] = 1'b1;
  assign \A[2][224] [1] = 1'b1;
  assign \A[2][224] [0] = 1'b1;
  assign \A[2][225] [4] = 1'b1;
  assign \A[2][225] [3] = 1'b1;
  assign \A[2][225] [2] = 1'b1;
  assign \A[2][225] [1] = 1'b1;
  assign \A[2][225] [0] = 1'b1;
  assign \A[2][226] [0] = 1'b1;
  assign \A[2][227] [4] = 1'b1;
  assign \A[2][227] [3] = 1'b1;
  assign \A[2][227] [2] = 1'b1;
  assign \A[2][227] [1] = 1'b1;
  assign \A[2][227] [0] = 1'b1;
  assign \A[2][228] [4] = 1'b1;
  assign \A[2][228] [3] = 1'b1;
  assign \A[2][228] [2] = 1'b1;
  assign \A[2][230] [4] = 1'b1;
  assign \A[2][230] [3] = 1'b1;
  assign \A[2][230] [2] = 1'b1;
  assign \A[2][230] [1] = 1'b1;
  assign \A[2][230] [0] = 1'b1;
  assign \A[2][231] [4] = 1'b1;
  assign \A[2][231] [3] = 1'b1;
  assign \A[2][231] [2] = 1'b1;
  assign \A[2][231] [1] = 1'b1;
  assign \A[2][232] [4] = 1'b1;
  assign \A[2][232] [3] = 1'b1;
  assign \A[2][232] [2] = 1'b1;
  assign \A[2][232] [1] = 1'b1;
  assign \A[2][232] [0] = 1'b1;
  assign \A[2][233] [4] = 1'b1;
  assign \A[2][233] [3] = 1'b1;
  assign \A[2][233] [2] = 1'b1;
  assign \A[2][233] [1] = 1'b1;
  assign \A[2][234] [4] = 1'b1;
  assign \A[2][234] [3] = 1'b1;
  assign \A[2][234] [2] = 1'b1;
  assign \A[2][235] [4] = 1'b1;
  assign \A[2][235] [3] = 1'b1;
  assign \A[2][235] [2] = 1'b1;
  assign \A[2][235] [1] = 1'b1;
  assign \A[2][235] [0] = 1'b1;
  assign \A[2][236] [4] = 1'b1;
  assign \A[2][236] [3] = 1'b1;
  assign \A[2][236] [2] = 1'b1;
  assign \A[2][238] [4] = 1'b1;
  assign \A[2][238] [3] = 1'b1;
  assign \A[2][238] [2] = 1'b1;
  assign \A[2][238] [1] = 1'b1;
  assign \A[2][238] [0] = 1'b1;
  assign \A[2][239] [0] = 1'b1;
  assign \A[2][240] [4] = 1'b1;
  assign \A[2][240] [3] = 1'b1;
  assign \A[2][240] [2] = 1'b1;
  assign \A[2][240] [1] = 1'b1;
  assign \A[2][240] [0] = 1'b1;
  assign \A[2][242] [4] = 1'b1;
  assign \A[2][242] [3] = 1'b1;
  assign \A[2][242] [2] = 1'b1;
  assign \A[2][242] [1] = 1'b1;
  assign \A[2][243] [4] = 1'b1;
  assign \A[2][243] [3] = 1'b1;
  assign \A[2][243] [2] = 1'b1;
  assign \A[2][243] [0] = 1'b1;
  assign \A[2][244] [4] = 1'b1;
  assign \A[2][244] [3] = 1'b1;
  assign \A[2][244] [2] = 1'b1;
  assign \A[2][245] [4] = 1'b1;
  assign \A[2][245] [3] = 1'b1;
  assign \A[2][245] [2] = 1'b1;
  assign \A[2][245] [1] = 1'b1;
  assign \A[2][245] [0] = 1'b1;
  assign \A[2][247] [4] = 1'b1;
  assign \A[2][247] [3] = 1'b1;
  assign \A[2][247] [2] = 1'b1;
  assign \A[2][247] [0] = 1'b1;
  assign \A[2][250] [0] = 1'b1;
  assign \A[2][251] [1] = 1'b1;
  assign \A[2][252] [4] = 1'b1;
  assign \A[2][252] [3] = 1'b1;
  assign \A[2][252] [2] = 1'b1;
  assign \A[2][252] [1] = 1'b1;
  assign \A[2][252] [0] = 1'b1;
  assign \A[2][253] [4] = 1'b1;
  assign \A[2][253] [3] = 1'b1;
  assign \A[2][253] [2] = 1'b1;
  assign \A[2][253] [1] = 1'b1;
  assign \A[2][253] [0] = 1'b1;
  assign \A[2][254] [4] = 1'b1;
  assign \A[2][254] [3] = 1'b1;
  assign \A[2][254] [2] = 1'b1;
  assign \A[2][254] [1] = 1'b1;
  assign \A[3][1] [0] = 1'b1;
  assign \A[3][2] [4] = 1'b1;
  assign \A[3][2] [3] = 1'b1;
  assign \A[3][2] [2] = 1'b1;
  assign \A[3][2] [1] = 1'b1;
  assign \A[3][2] [0] = 1'b1;
  assign \A[3][4] [0] = 1'b1;
  assign \A[3][5] [4] = 1'b1;
  assign \A[3][5] [3] = 1'b1;
  assign \A[3][5] [2] = 1'b1;
  assign \A[3][5] [1] = 1'b1;
  assign \A[3][6] [4] = 1'b1;
  assign \A[3][6] [3] = 1'b1;
  assign \A[3][6] [2] = 1'b1;
  assign \A[3][6] [0] = 1'b1;
  assign \A[3][7] [4] = 1'b1;
  assign \A[3][7] [3] = 1'b1;
  assign \A[3][7] [2] = 1'b1;
  assign \A[3][7] [1] = 1'b1;
  assign \A[3][7] [0] = 1'b1;
  assign \A[3][8] [1] = 1'b1;
  assign \A[3][9] [4] = 1'b1;
  assign \A[3][9] [3] = 1'b1;
  assign \A[3][9] [2] = 1'b1;
  assign \A[3][9] [1] = 1'b1;
  assign \A[3][10] [4] = 1'b1;
  assign \A[3][10] [3] = 1'b1;
  assign \A[3][10] [2] = 1'b1;
  assign \A[3][10] [1] = 1'b1;
  assign \A[3][10] [0] = 1'b1;
  assign \A[3][11] [4] = 1'b1;
  assign \A[3][11] [3] = 1'b1;
  assign \A[3][11] [2] = 1'b1;
  assign \A[3][11] [1] = 1'b1;
  assign \A[3][11] [0] = 1'b1;
  assign \A[3][13] [4] = 1'b1;
  assign \A[3][13] [3] = 1'b1;
  assign \A[3][13] [2] = 1'b1;
  assign \A[3][13] [1] = 1'b1;
  assign \A[3][13] [0] = 1'b1;
  assign \A[3][14] [1] = 1'b1;
  assign \A[3][15] [1] = 1'b1;
  assign \A[3][15] [0] = 1'b1;
  assign \A[3][16] [4] = 1'b1;
  assign \A[3][16] [3] = 1'b1;
  assign \A[3][16] [2] = 1'b1;
  assign \A[3][16] [1] = 1'b1;
  assign \A[3][16] [0] = 1'b1;
  assign \A[3][18] [4] = 1'b1;
  assign \A[3][18] [3] = 1'b1;
  assign \A[3][18] [2] = 1'b1;
  assign \A[3][18] [1] = 1'b1;
  assign \A[3][20] [4] = 1'b1;
  assign \A[3][20] [3] = 1'b1;
  assign \A[3][20] [2] = 1'b1;
  assign \A[3][20] [1] = 1'b1;
  assign \A[3][25] [0] = 1'b1;
  assign \A[3][26] [4] = 1'b1;
  assign \A[3][26] [3] = 1'b1;
  assign \A[3][26] [2] = 1'b1;
  assign \A[3][26] [1] = 1'b1;
  assign \A[3][28] [1] = 1'b1;
  assign \A[3][29] [4] = 1'b1;
  assign \A[3][29] [3] = 1'b1;
  assign \A[3][29] [2] = 1'b1;
  assign \A[3][29] [1] = 1'b1;
  assign \A[3][31] [0] = 1'b1;
  assign \A[3][33] [4] = 1'b1;
  assign \A[3][33] [3] = 1'b1;
  assign \A[3][33] [2] = 1'b1;
  assign \A[3][33] [1] = 1'b1;
  assign \A[3][34] [4] = 1'b1;
  assign \A[3][34] [3] = 1'b1;
  assign \A[3][34] [2] = 1'b1;
  assign \A[3][34] [1] = 1'b1;
  assign \A[3][34] [0] = 1'b1;
  assign \A[3][35] [4] = 1'b1;
  assign \A[3][35] [3] = 1'b1;
  assign \A[3][35] [2] = 1'b1;
  assign \A[3][35] [1] = 1'b1;
  assign \A[3][35] [0] = 1'b1;
  assign \A[3][36] [4] = 1'b1;
  assign \A[3][36] [3] = 1'b1;
  assign \A[3][36] [2] = 1'b1;
  assign \A[3][36] [1] = 1'b1;
  assign \A[3][36] [0] = 1'b1;
  assign \A[3][37] [4] = 1'b1;
  assign \A[3][37] [3] = 1'b1;
  assign \A[3][37] [2] = 1'b1;
  assign \A[3][37] [1] = 1'b1;
  assign \A[3][37] [0] = 1'b1;
  assign \A[3][38] [0] = 1'b1;
  assign \A[3][39] [4] = 1'b1;
  assign \A[3][39] [3] = 1'b1;
  assign \A[3][39] [2] = 1'b1;
  assign \A[3][39] [1] = 1'b1;
  assign \A[3][41] [4] = 1'b1;
  assign \A[3][41] [3] = 1'b1;
  assign \A[3][41] [2] = 1'b1;
  assign \A[3][41] [1] = 1'b1;
  assign \A[3][41] [0] = 1'b1;
  assign \A[3][43] [4] = 1'b1;
  assign \A[3][43] [3] = 1'b1;
  assign \A[3][43] [2] = 1'b1;
  assign \A[3][43] [1] = 1'b1;
  assign \A[3][43] [0] = 1'b1;
  assign \A[3][44] [0] = 1'b1;
  assign \A[3][45] [1] = 1'b1;
  assign \A[3][46] [0] = 1'b1;
  assign \A[3][47] [4] = 1'b1;
  assign \A[3][47] [3] = 1'b1;
  assign \A[3][47] [2] = 1'b1;
  assign \A[3][47] [1] = 1'b1;
  assign \A[3][48] [4] = 1'b1;
  assign \A[3][48] [3] = 1'b1;
  assign \A[3][48] [2] = 1'b1;
  assign \A[3][48] [1] = 1'b1;
  assign \A[3][48] [0] = 1'b1;
  assign \A[3][49] [4] = 1'b1;
  assign \A[3][49] [3] = 1'b1;
  assign \A[3][49] [2] = 1'b1;
  assign \A[3][49] [1] = 1'b1;
  assign \A[3][49] [0] = 1'b1;
  assign \A[3][50] [4] = 1'b1;
  assign \A[3][50] [3] = 1'b1;
  assign \A[3][50] [2] = 1'b1;
  assign \A[3][50] [1] = 1'b1;
  assign \A[3][50] [0] = 1'b1;
  assign \A[3][52] [4] = 1'b1;
  assign \A[3][52] [3] = 1'b1;
  assign \A[3][52] [2] = 1'b1;
  assign \A[3][52] [1] = 1'b1;
  assign \A[3][52] [0] = 1'b1;
  assign \A[3][53] [1] = 1'b1;
  assign \A[3][54] [4] = 1'b1;
  assign \A[3][54] [3] = 1'b1;
  assign \A[3][54] [2] = 1'b1;
  assign \A[3][54] [0] = 1'b1;
  assign \A[3][55] [4] = 1'b1;
  assign \A[3][55] [3] = 1'b1;
  assign \A[3][55] [2] = 1'b1;
  assign \A[3][55] [1] = 1'b1;
  assign \A[3][55] [0] = 1'b1;
  assign \A[3][56] [1] = 1'b1;
  assign \A[3][56] [0] = 1'b1;
  assign \A[3][57] [0] = 1'b1;
  assign \A[3][58] [0] = 1'b1;
  assign \A[3][61] [0] = 1'b1;
  assign \A[3][64] [0] = 1'b1;
  assign \A[3][65] [1] = 1'b1;
  assign \A[3][66] [4] = 1'b1;
  assign \A[3][66] [3] = 1'b1;
  assign \A[3][66] [2] = 1'b1;
  assign \A[3][66] [1] = 1'b1;
  assign \A[3][66] [0] = 1'b1;
  assign \A[3][67] [4] = 1'b1;
  assign \A[3][67] [3] = 1'b1;
  assign \A[3][67] [2] = 1'b1;
  assign \A[3][67] [1] = 1'b1;
  assign \A[3][67] [0] = 1'b1;
  assign \A[3][68] [0] = 1'b1;
  assign \A[3][69] [1] = 1'b1;
  assign \A[3][70] [1] = 1'b1;
  assign \A[3][70] [0] = 1'b1;
  assign \A[3][72] [1] = 1'b1;
  assign \A[3][72] [0] = 1'b1;
  assign \A[3][73] [4] = 1'b1;
  assign \A[3][73] [3] = 1'b1;
  assign \A[3][73] [2] = 1'b1;
  assign \A[3][73] [1] = 1'b1;
  assign \A[3][74] [4] = 1'b1;
  assign \A[3][74] [3] = 1'b1;
  assign \A[3][74] [2] = 1'b1;
  assign \A[3][76] [1] = 1'b1;
  assign \A[3][77] [0] = 1'b1;
  assign \A[3][78] [4] = 1'b1;
  assign \A[3][78] [3] = 1'b1;
  assign \A[3][78] [2] = 1'b1;
  assign \A[3][78] [1] = 1'b1;
  assign \A[3][79] [1] = 1'b1;
  assign \A[3][80] [4] = 1'b1;
  assign \A[3][80] [3] = 1'b1;
  assign \A[3][80] [2] = 1'b1;
  assign \A[3][80] [1] = 1'b1;
  assign \A[3][80] [0] = 1'b1;
  assign \A[3][81] [0] = 1'b1;
  assign \A[3][83] [4] = 1'b1;
  assign \A[3][83] [3] = 1'b1;
  assign \A[3][83] [2] = 1'b1;
  assign \A[3][83] [1] = 1'b1;
  assign \A[3][83] [0] = 1'b1;
  assign \A[3][84] [4] = 1'b1;
  assign \A[3][84] [3] = 1'b1;
  assign \A[3][84] [2] = 1'b1;
  assign \A[3][84] [1] = 1'b1;
  assign \A[3][84] [0] = 1'b1;
  assign \A[3][85] [1] = 1'b1;
  assign \A[3][86] [0] = 1'b1;
  assign \A[3][87] [0] = 1'b1;
  assign \A[3][89] [4] = 1'b1;
  assign \A[3][89] [3] = 1'b1;
  assign \A[3][89] [2] = 1'b1;
  assign \A[3][89] [1] = 1'b1;
  assign \A[3][90] [0] = 1'b1;
  assign \A[3][91] [1] = 1'b1;
  assign \A[3][92] [4] = 1'b1;
  assign \A[3][92] [3] = 1'b1;
  assign \A[3][92] [2] = 1'b1;
  assign \A[3][92] [1] = 1'b1;
  assign \A[3][92] [0] = 1'b1;
  assign \A[3][93] [4] = 1'b1;
  assign \A[3][93] [3] = 1'b1;
  assign \A[3][93] [2] = 1'b1;
  assign \A[3][93] [1] = 1'b1;
  assign \A[3][93] [0] = 1'b1;
  assign \A[3][95] [4] = 1'b1;
  assign \A[3][95] [3] = 1'b1;
  assign \A[3][95] [2] = 1'b1;
  assign \A[3][95] [1] = 1'b1;
  assign \A[3][95] [0] = 1'b1;
  assign \A[3][96] [4] = 1'b1;
  assign \A[3][96] [3] = 1'b1;
  assign \A[3][96] [2] = 1'b1;
  assign \A[3][96] [1] = 1'b1;
  assign \A[3][96] [0] = 1'b1;
  assign \A[3][98] [4] = 1'b1;
  assign \A[3][98] [3] = 1'b1;
  assign \A[3][98] [2] = 1'b1;
  assign \A[3][98] [1] = 1'b1;
  assign \A[3][98] [0] = 1'b1;
  assign \A[3][99] [4] = 1'b1;
  assign \A[3][99] [3] = 1'b1;
  assign \A[3][99] [2] = 1'b1;
  assign \A[3][99] [1] = 1'b1;
  assign \A[3][99] [0] = 1'b1;
  assign \A[3][100] [4] = 1'b1;
  assign \A[3][100] [3] = 1'b1;
  assign \A[3][100] [2] = 1'b1;
  assign \A[3][100] [1] = 1'b1;
  assign \A[3][101] [4] = 1'b1;
  assign \A[3][101] [3] = 1'b1;
  assign \A[3][101] [2] = 1'b1;
  assign \A[3][101] [1] = 1'b1;
  assign \A[3][101] [0] = 1'b1;
  assign \A[3][102] [1] = 1'b1;
  assign \A[3][104] [0] = 1'b1;
  assign \A[3][105] [4] = 1'b1;
  assign \A[3][105] [3] = 1'b1;
  assign \A[3][105] [2] = 1'b1;
  assign \A[3][105] [1] = 1'b1;
  assign \A[3][105] [0] = 1'b1;
  assign \A[3][106] [1] = 1'b1;
  assign \A[3][108] [2] = 1'b1;
  assign \A[3][109] [1] = 1'b1;
  assign \A[3][109] [0] = 1'b1;
  assign \A[3][110] [4] = 1'b1;
  assign \A[3][110] [3] = 1'b1;
  assign \A[3][110] [2] = 1'b1;
  assign \A[3][110] [0] = 1'b1;
  assign \A[3][111] [4] = 1'b1;
  assign \A[3][111] [3] = 1'b1;
  assign \A[3][111] [2] = 1'b1;
  assign \A[3][111] [1] = 1'b1;
  assign \A[3][111] [0] = 1'b1;
  assign \A[3][113] [0] = 1'b1;
  assign \A[3][114] [4] = 1'b1;
  assign \A[3][114] [3] = 1'b1;
  assign \A[3][114] [2] = 1'b1;
  assign \A[3][114] [0] = 1'b1;
  assign \A[3][115] [4] = 1'b1;
  assign \A[3][115] [3] = 1'b1;
  assign \A[3][115] [2] = 1'b1;
  assign \A[3][115] [1] = 1'b1;
  assign \A[3][115] [0] = 1'b1;
  assign \A[3][117] [4] = 1'b1;
  assign \A[3][117] [3] = 1'b1;
  assign \A[3][117] [2] = 1'b1;
  assign \A[3][117] [1] = 1'b1;
  assign \A[3][117] [0] = 1'b1;
  assign \A[3][119] [4] = 1'b1;
  assign \A[3][119] [3] = 1'b1;
  assign \A[3][119] [2] = 1'b1;
  assign \A[3][119] [1] = 1'b1;
  assign \A[3][119] [0] = 1'b1;
  assign \A[3][120] [4] = 1'b1;
  assign \A[3][120] [3] = 1'b1;
  assign \A[3][120] [2] = 1'b1;
  assign \A[3][120] [1] = 1'b1;
  assign \A[3][121] [0] = 1'b1;
  assign \A[3][123] [1] = 1'b1;
  assign \A[3][127] [0] = 1'b1;
  assign \A[3][128] [4] = 1'b1;
  assign \A[3][128] [3] = 1'b1;
  assign \A[3][128] [2] = 1'b1;
  assign \A[3][128] [1] = 1'b1;
  assign \A[3][128] [0] = 1'b1;
  assign \A[3][129] [4] = 1'b1;
  assign \A[3][129] [3] = 1'b1;
  assign \A[3][129] [2] = 1'b1;
  assign \A[3][129] [1] = 1'b1;
  assign \A[3][130] [4] = 1'b1;
  assign \A[3][130] [3] = 1'b1;
  assign \A[3][130] [2] = 1'b1;
  assign \A[3][130] [1] = 1'b1;
  assign \A[3][132] [4] = 1'b1;
  assign \A[3][132] [3] = 1'b1;
  assign \A[3][132] [2] = 1'b1;
  assign \A[3][132] [1] = 1'b1;
  assign \A[3][132] [0] = 1'b1;
  assign \A[3][135] [4] = 1'b1;
  assign \A[3][135] [3] = 1'b1;
  assign \A[3][135] [2] = 1'b1;
  assign \A[3][135] [1] = 1'b1;
  assign \A[3][136] [1] = 1'b1;
  assign \A[3][137] [0] = 1'b1;
  assign \A[3][139] [0] = 1'b1;
  assign \A[3][140] [4] = 1'b1;
  assign \A[3][140] [3] = 1'b1;
  assign \A[3][140] [2] = 1'b1;
  assign \A[3][140] [1] = 1'b1;
  assign \A[3][141] [4] = 1'b1;
  assign \A[3][141] [3] = 1'b1;
  assign \A[3][141] [2] = 1'b1;
  assign \A[3][141] [1] = 1'b1;
  assign \A[3][142] [4] = 1'b1;
  assign \A[3][142] [3] = 1'b1;
  assign \A[3][142] [2] = 1'b1;
  assign \A[3][142] [1] = 1'b1;
  assign \A[3][142] [0] = 1'b1;
  assign \A[3][144] [4] = 1'b1;
  assign \A[3][144] [3] = 1'b1;
  assign \A[3][144] [2] = 1'b1;
  assign \A[3][144] [1] = 1'b1;
  assign \A[3][145] [1] = 1'b1;
  assign \A[3][146] [4] = 1'b1;
  assign \A[3][146] [3] = 1'b1;
  assign \A[3][146] [2] = 1'b1;
  assign \A[3][146] [1] = 1'b1;
  assign \A[3][146] [0] = 1'b1;
  assign \A[3][147] [4] = 1'b1;
  assign \A[3][147] [3] = 1'b1;
  assign \A[3][147] [2] = 1'b1;
  assign \A[3][147] [1] = 1'b1;
  assign \A[3][147] [0] = 1'b1;
  assign \A[3][148] [0] = 1'b1;
  assign \A[3][149] [1] = 1'b1;
  assign \A[3][149] [0] = 1'b1;
  assign \A[3][150] [1] = 1'b1;
  assign \A[3][151] [4] = 1'b1;
  assign \A[3][151] [3] = 1'b1;
  assign \A[3][151] [2] = 1'b1;
  assign \A[3][151] [1] = 1'b1;
  assign \A[3][151] [0] = 1'b1;
  assign \A[3][152] [0] = 1'b1;
  assign \A[3][154] [1] = 1'b1;
  assign \A[3][155] [4] = 1'b1;
  assign \A[3][155] [3] = 1'b1;
  assign \A[3][155] [2] = 1'b1;
  assign \A[3][155] [1] = 1'b1;
  assign \A[3][155] [0] = 1'b1;
  assign \A[3][156] [4] = 1'b1;
  assign \A[3][156] [3] = 1'b1;
  assign \A[3][156] [2] = 1'b1;
  assign \A[3][156] [1] = 1'b1;
  assign \A[3][156] [0] = 1'b1;
  assign \A[3][157] [4] = 1'b1;
  assign \A[3][157] [3] = 1'b1;
  assign \A[3][157] [2] = 1'b1;
  assign \A[3][157] [1] = 1'b1;
  assign \A[3][157] [0] = 1'b1;
  assign \A[3][158] [4] = 1'b1;
  assign \A[3][158] [3] = 1'b1;
  assign \A[3][158] [2] = 1'b1;
  assign \A[3][158] [1] = 1'b1;
  assign \A[3][159] [4] = 1'b1;
  assign \A[3][159] [3] = 1'b1;
  assign \A[3][159] [2] = 1'b1;
  assign \A[3][159] [1] = 1'b1;
  assign \A[3][160] [4] = 1'b1;
  assign \A[3][160] [3] = 1'b1;
  assign \A[3][160] [2] = 1'b1;
  assign \A[3][160] [1] = 1'b1;
  assign \A[3][160] [0] = 1'b1;
  assign \A[3][161] [4] = 1'b1;
  assign \A[3][161] [3] = 1'b1;
  assign \A[3][161] [2] = 1'b1;
  assign \A[3][161] [0] = 1'b1;
  assign \A[3][162] [0] = 1'b1;
  assign \A[3][164] [0] = 1'b1;
  assign \A[3][165] [4] = 1'b1;
  assign \A[3][165] [3] = 1'b1;
  assign \A[3][165] [2] = 1'b1;
  assign \A[3][165] [1] = 1'b1;
  assign \A[3][165] [0] = 1'b1;
  assign \A[3][168] [4] = 1'b1;
  assign \A[3][168] [3] = 1'b1;
  assign \A[3][168] [2] = 1'b1;
  assign \A[3][168] [1] = 1'b1;
  assign \A[3][168] [0] = 1'b1;
  assign \A[3][170] [4] = 1'b1;
  assign \A[3][170] [3] = 1'b1;
  assign \A[3][170] [2] = 1'b1;
  assign \A[3][170] [0] = 1'b1;
  assign \A[3][172] [0] = 1'b1;
  assign \A[3][174] [4] = 1'b1;
  assign \A[3][174] [3] = 1'b1;
  assign \A[3][174] [2] = 1'b1;
  assign \A[3][174] [1] = 1'b1;
  assign \A[3][175] [4] = 1'b1;
  assign \A[3][175] [3] = 1'b1;
  assign \A[3][175] [2] = 1'b1;
  assign \A[3][175] [0] = 1'b1;
  assign \A[3][178] [0] = 1'b1;
  assign \A[3][179] [1] = 1'b1;
  assign \A[3][180] [1] = 1'b1;
  assign \A[3][181] [0] = 1'b1;
  assign \A[3][183] [4] = 1'b1;
  assign \A[3][183] [3] = 1'b1;
  assign \A[3][183] [2] = 1'b1;
  assign \A[3][183] [1] = 1'b1;
  assign \A[3][183] [0] = 1'b1;
  assign \A[3][184] [4] = 1'b1;
  assign \A[3][184] [3] = 1'b1;
  assign \A[3][184] [2] = 1'b1;
  assign \A[3][184] [1] = 1'b1;
  assign \A[3][185] [4] = 1'b1;
  assign \A[3][185] [3] = 1'b1;
  assign \A[3][185] [2] = 1'b1;
  assign \A[3][185] [1] = 1'b1;
  assign \A[3][185] [0] = 1'b1;
  assign \A[3][186] [1] = 1'b1;
  assign \A[3][187] [1] = 1'b1;
  assign \A[3][188] [4] = 1'b1;
  assign \A[3][188] [3] = 1'b1;
  assign \A[3][188] [2] = 1'b1;
  assign \A[3][188] [1] = 1'b1;
  assign \A[3][188] [0] = 1'b1;
  assign \A[3][191] [4] = 1'b1;
  assign \A[3][191] [3] = 1'b1;
  assign \A[3][191] [2] = 1'b1;
  assign \A[3][191] [1] = 1'b1;
  assign \A[3][192] [0] = 1'b1;
  assign \A[3][194] [4] = 1'b1;
  assign \A[3][194] [3] = 1'b1;
  assign \A[3][194] [2] = 1'b1;
  assign \A[3][194] [1] = 1'b1;
  assign \A[3][195] [1] = 1'b1;
  assign \A[3][197] [1] = 1'b1;
  assign \A[3][198] [4] = 1'b1;
  assign \A[3][198] [3] = 1'b1;
  assign \A[3][198] [2] = 1'b1;
  assign \A[3][198] [0] = 1'b1;
  assign \A[3][200] [4] = 1'b1;
  assign \A[3][200] [3] = 1'b1;
  assign \A[3][200] [2] = 1'b1;
  assign \A[3][200] [1] = 1'b1;
  assign \A[3][200] [0] = 1'b1;
  assign \A[3][201] [0] = 1'b1;
  assign \A[3][203] [4] = 1'b1;
  assign \A[3][203] [3] = 1'b1;
  assign \A[3][203] [2] = 1'b1;
  assign \A[3][203] [1] = 1'b1;
  assign \A[3][204] [0] = 1'b1;
  assign \A[3][205] [4] = 1'b1;
  assign \A[3][205] [3] = 1'b1;
  assign \A[3][205] [2] = 1'b1;
  assign \A[3][205] [1] = 1'b1;
  assign \A[3][205] [0] = 1'b1;
  assign \A[3][206] [4] = 1'b1;
  assign \A[3][206] [3] = 1'b1;
  assign \A[3][206] [2] = 1'b1;
  assign \A[3][206] [1] = 1'b1;
  assign \A[3][209] [4] = 1'b1;
  assign \A[3][209] [3] = 1'b1;
  assign \A[3][209] [2] = 1'b1;
  assign \A[3][209] [1] = 1'b1;
  assign \A[3][209] [0] = 1'b1;
  assign \A[3][210] [4] = 1'b1;
  assign \A[3][210] [3] = 1'b1;
  assign \A[3][210] [2] = 1'b1;
  assign \A[3][210] [1] = 1'b1;
  assign \A[3][210] [0] = 1'b1;
  assign \A[3][211] [1] = 1'b1;
  assign \A[3][212] [4] = 1'b1;
  assign \A[3][212] [3] = 1'b1;
  assign \A[3][212] [2] = 1'b1;
  assign \A[3][212] [1] = 1'b1;
  assign \A[3][212] [0] = 1'b1;
  assign \A[3][214] [4] = 1'b1;
  assign \A[3][214] [3] = 1'b1;
  assign \A[3][214] [2] = 1'b1;
  assign \A[3][214] [1] = 1'b1;
  assign \A[3][215] [4] = 1'b1;
  assign \A[3][215] [3] = 1'b1;
  assign \A[3][215] [2] = 1'b1;
  assign \A[3][215] [1] = 1'b1;
  assign \A[3][215] [0] = 1'b1;
  assign \A[3][216] [1] = 1'b1;
  assign \A[3][218] [4] = 1'b1;
  assign \A[3][218] [3] = 1'b1;
  assign \A[3][218] [2] = 1'b1;
  assign \A[3][218] [1] = 1'b1;
  assign \A[3][218] [0] = 1'b1;
  assign \A[3][219] [4] = 1'b1;
  assign \A[3][219] [3] = 1'b1;
  assign \A[3][219] [2] = 1'b1;
  assign \A[3][219] [1] = 1'b1;
  assign \A[3][219] [0] = 1'b1;
  assign \A[3][220] [4] = 1'b1;
  assign \A[3][220] [3] = 1'b1;
  assign \A[3][220] [2] = 1'b1;
  assign \A[3][220] [1] = 1'b1;
  assign \A[3][220] [0] = 1'b1;
  assign \A[3][221] [4] = 1'b1;
  assign \A[3][221] [3] = 1'b1;
  assign \A[3][221] [2] = 1'b1;
  assign \A[3][221] [1] = 1'b1;
  assign \A[3][221] [0] = 1'b1;
  assign \A[3][222] [4] = 1'b1;
  assign \A[3][222] [3] = 1'b1;
  assign \A[3][222] [2] = 1'b1;
  assign \A[3][222] [1] = 1'b1;
  assign \A[3][222] [0] = 1'b1;
  assign \A[3][223] [0] = 1'b1;
  assign \A[3][224] [0] = 1'b1;
  assign \A[3][225] [0] = 1'b1;
  assign \A[3][226] [4] = 1'b1;
  assign \A[3][226] [3] = 1'b1;
  assign \A[3][226] [2] = 1'b1;
  assign \A[3][226] [1] = 1'b1;
  assign \A[3][226] [0] = 1'b1;
  assign \A[3][229] [4] = 1'b1;
  assign \A[3][229] [3] = 1'b1;
  assign \A[3][229] [2] = 1'b1;
  assign \A[3][229] [1] = 1'b1;
  assign \A[3][229] [0] = 1'b1;
  assign \A[3][230] [4] = 1'b1;
  assign \A[3][230] [3] = 1'b1;
  assign \A[3][230] [2] = 1'b1;
  assign \A[3][230] [1] = 1'b1;
  assign \A[3][233] [0] = 1'b1;
  assign \A[3][235] [0] = 1'b1;
  assign \A[3][238] [4] = 1'b1;
  assign \A[3][238] [3] = 1'b1;
  assign \A[3][238] [2] = 1'b1;
  assign \A[3][238] [1] = 1'b1;
  assign \A[3][238] [0] = 1'b1;
  assign \A[3][239] [4] = 1'b1;
  assign \A[3][239] [3] = 1'b1;
  assign \A[3][239] [2] = 1'b1;
  assign \A[3][239] [1] = 1'b1;
  assign \A[3][239] [0] = 1'b1;
  assign \A[3][240] [1] = 1'b1;
  assign \A[3][242] [4] = 1'b1;
  assign \A[3][242] [3] = 1'b1;
  assign \A[3][242] [2] = 1'b1;
  assign \A[3][242] [0] = 1'b1;
  assign \A[3][243] [1] = 1'b1;
  assign \A[3][244] [1] = 1'b1;
  assign \A[3][246] [4] = 1'b1;
  assign \A[3][246] [3] = 1'b1;
  assign \A[3][246] [2] = 1'b1;
  assign \A[3][246] [1] = 1'b1;
  assign \A[3][246] [0] = 1'b1;
  assign \A[3][247] [0] = 1'b1;
  assign \A[3][248] [4] = 1'b1;
  assign \A[3][248] [3] = 1'b1;
  assign \A[3][248] [2] = 1'b1;
  assign \A[3][248] [1] = 1'b1;
  assign \A[3][248] [0] = 1'b1;
  assign \A[3][249] [0] = 1'b1;
  assign \A[3][251] [4] = 1'b1;
  assign \A[3][251] [3] = 1'b1;
  assign \A[3][251] [2] = 1'b1;
  assign \A[3][251] [1] = 1'b1;
  assign \A[3][255] [4] = 1'b1;
  assign \A[3][255] [3] = 1'b1;
  assign \A[3][255] [2] = 1'b1;
  assign \A[3][255] [1] = 1'b1;
  assign \A[3][255] [0] = 1'b1;
  assign \A[4][0] [4] = 1'b1;
  assign \A[4][0] [3] = 1'b1;
  assign \A[4][0] [2] = 1'b1;
  assign \A[4][0] [1] = 1'b1;
  assign \A[4][0] [0] = 1'b1;
  assign \A[4][1] [4] = 1'b1;
  assign \A[4][1] [3] = 1'b1;
  assign \A[4][1] [2] = 1'b1;
  assign \A[4][1] [1] = 1'b1;
  assign \A[4][1] [0] = 1'b1;
  assign \A[4][3] [0] = 1'b1;
  assign \A[4][5] [4] = 1'b1;
  assign \A[4][5] [3] = 1'b1;
  assign \A[4][5] [2] = 1'b1;
  assign \A[4][5] [1] = 1'b1;
  assign \A[4][6] [4] = 1'b1;
  assign \A[4][6] [3] = 1'b1;
  assign \A[4][6] [2] = 1'b1;
  assign \A[4][6] [1] = 1'b1;
  assign \A[4][7] [4] = 1'b1;
  assign \A[4][7] [3] = 1'b1;
  assign \A[4][7] [2] = 1'b1;
  assign \A[4][7] [1] = 1'b1;
  assign \A[4][7] [0] = 1'b1;
  assign \A[4][8] [0] = 1'b1;
  assign \A[4][9] [4] = 1'b1;
  assign \A[4][9] [3] = 1'b1;
  assign \A[4][9] [2] = 1'b1;
  assign \A[4][9] [1] = 1'b1;
  assign \A[4][9] [0] = 1'b1;
  assign \A[4][10] [4] = 1'b1;
  assign \A[4][10] [3] = 1'b1;
  assign \A[4][10] [2] = 1'b1;
  assign \A[4][10] [1] = 1'b1;
  assign \A[4][10] [0] = 1'b1;
  assign \A[4][11] [4] = 1'b1;
  assign \A[4][11] [3] = 1'b1;
  assign \A[4][11] [2] = 1'b1;
  assign \A[4][11] [0] = 1'b1;
  assign \A[4][14] [0] = 1'b1;
  assign \A[4][15] [0] = 1'b1;
  assign \A[4][16] [4] = 1'b1;
  assign \A[4][16] [3] = 1'b1;
  assign \A[4][16] [2] = 1'b1;
  assign \A[4][16] [1] = 1'b1;
  assign \A[4][16] [0] = 1'b1;
  assign \A[4][19] [4] = 1'b1;
  assign \A[4][19] [3] = 1'b1;
  assign \A[4][19] [2] = 1'b1;
  assign \A[4][19] [1] = 1'b1;
  assign \A[4][19] [0] = 1'b1;
  assign \A[4][20] [4] = 1'b1;
  assign \A[4][20] [3] = 1'b1;
  assign \A[4][20] [2] = 1'b1;
  assign \A[4][20] [1] = 1'b1;
  assign \A[4][20] [0] = 1'b1;
  assign \A[4][21] [0] = 1'b1;
  assign \A[4][23] [4] = 1'b1;
  assign \A[4][23] [3] = 1'b1;
  assign \A[4][23] [2] = 1'b1;
  assign \A[4][23] [1] = 1'b1;
  assign \A[4][24] [0] = 1'b1;
  assign \A[4][25] [4] = 1'b1;
  assign \A[4][25] [3] = 1'b1;
  assign \A[4][25] [2] = 1'b1;
  assign \A[4][25] [1] = 1'b1;
  assign \A[4][25] [0] = 1'b1;
  assign \A[4][26] [4] = 1'b1;
  assign \A[4][26] [3] = 1'b1;
  assign \A[4][26] [2] = 1'b1;
  assign \A[4][26] [0] = 1'b1;
  assign \A[4][28] [4] = 1'b1;
  assign \A[4][28] [3] = 1'b1;
  assign \A[4][28] [2] = 1'b1;
  assign \A[4][28] [1] = 1'b1;
  assign \A[4][28] [0] = 1'b1;
  assign \A[4][29] [1] = 1'b1;
  assign \A[4][30] [1] = 1'b1;
  assign \A[4][30] [0] = 1'b1;
  assign \A[4][31] [4] = 1'b1;
  assign \A[4][31] [3] = 1'b1;
  assign \A[4][31] [2] = 1'b1;
  assign \A[4][31] [0] = 1'b1;
  assign \A[4][32] [4] = 1'b1;
  assign \A[4][32] [3] = 1'b1;
  assign \A[4][32] [2] = 1'b1;
  assign \A[4][32] [1] = 1'b1;
  assign \A[4][33] [4] = 1'b1;
  assign \A[4][33] [3] = 1'b1;
  assign \A[4][33] [2] = 1'b1;
  assign \A[4][33] [1] = 1'b1;
  assign \A[4][34] [4] = 1'b1;
  assign \A[4][34] [3] = 1'b1;
  assign \A[4][34] [2] = 1'b1;
  assign \A[4][34] [1] = 1'b1;
  assign \A[4][35] [4] = 1'b1;
  assign \A[4][35] [3] = 1'b1;
  assign \A[4][35] [2] = 1'b1;
  assign \A[4][35] [1] = 1'b1;
  assign \A[4][35] [0] = 1'b1;
  assign \A[4][37] [4] = 1'b1;
  assign \A[4][37] [3] = 1'b1;
  assign \A[4][37] [2] = 1'b1;
  assign \A[4][37] [0] = 1'b1;
  assign \A[4][39] [4] = 1'b1;
  assign \A[4][39] [3] = 1'b1;
  assign \A[4][39] [2] = 1'b1;
  assign \A[4][39] [1] = 1'b1;
  assign \A[4][39] [0] = 1'b1;
  assign \A[4][40] [4] = 1'b1;
  assign \A[4][40] [3] = 1'b1;
  assign \A[4][40] [2] = 1'b1;
  assign \A[4][40] [1] = 1'b1;
  assign \A[4][42] [4] = 1'b1;
  assign \A[4][42] [3] = 1'b1;
  assign \A[4][42] [2] = 1'b1;
  assign \A[4][42] [0] = 1'b1;
  assign \A[4][43] [4] = 1'b1;
  assign \A[4][43] [3] = 1'b1;
  assign \A[4][43] [2] = 1'b1;
  assign \A[4][43] [1] = 1'b1;
  assign \A[4][44] [2] = 1'b1;
  assign \A[4][46] [0] = 1'b1;
  assign \A[4][48] [4] = 1'b1;
  assign \A[4][48] [3] = 1'b1;
  assign \A[4][48] [2] = 1'b1;
  assign \A[4][48] [1] = 1'b1;
  assign \A[4][48] [0] = 1'b1;
  assign \A[4][49] [1] = 1'b1;
  assign \A[4][51] [4] = 1'b1;
  assign \A[4][51] [3] = 1'b1;
  assign \A[4][51] [2] = 1'b1;
  assign \A[4][51] [1] = 1'b1;
  assign \A[4][51] [0] = 1'b1;
  assign \A[4][52] [4] = 1'b1;
  assign \A[4][52] [3] = 1'b1;
  assign \A[4][52] [2] = 1'b1;
  assign \A[4][52] [1] = 1'b1;
  assign \A[4][53] [4] = 1'b1;
  assign \A[4][53] [3] = 1'b1;
  assign \A[4][53] [2] = 1'b1;
  assign \A[4][53] [1] = 1'b1;
  assign \A[4][53] [0] = 1'b1;
  assign \A[4][54] [4] = 1'b1;
  assign \A[4][54] [3] = 1'b1;
  assign \A[4][54] [2] = 1'b1;
  assign \A[4][54] [1] = 1'b1;
  assign \A[4][54] [0] = 1'b1;
  assign \A[4][55] [4] = 1'b1;
  assign \A[4][55] [3] = 1'b1;
  assign \A[4][55] [2] = 1'b1;
  assign \A[4][56] [1] = 1'b1;
  assign \A[4][56] [0] = 1'b1;
  assign \A[4][57] [0] = 1'b1;
  assign \A[4][58] [0] = 1'b1;
  assign \A[4][59] [4] = 1'b1;
  assign \A[4][59] [3] = 1'b1;
  assign \A[4][59] [2] = 1'b1;
  assign \A[4][59] [1] = 1'b1;
  assign \A[4][59] [0] = 1'b1;
  assign \A[4][60] [4] = 1'b1;
  assign \A[4][60] [3] = 1'b1;
  assign \A[4][60] [2] = 1'b1;
  assign \A[4][60] [1] = 1'b1;
  assign \A[4][60] [0] = 1'b1;
  assign \A[4][61] [1] = 1'b1;
  assign \A[4][62] [0] = 1'b1;
  assign \A[4][64] [1] = 1'b1;
  assign \A[4][65] [0] = 1'b1;
  assign \A[4][66] [4] = 1'b1;
  assign \A[4][66] [3] = 1'b1;
  assign \A[4][66] [2] = 1'b1;
  assign \A[4][66] [1] = 1'b1;
  assign \A[4][67] [4] = 1'b1;
  assign \A[4][67] [3] = 1'b1;
  assign \A[4][67] [2] = 1'b1;
  assign \A[4][67] [1] = 1'b1;
  assign \A[4][68] [4] = 1'b1;
  assign \A[4][68] [3] = 1'b1;
  assign \A[4][68] [2] = 1'b1;
  assign \A[4][68] [1] = 1'b1;
  assign \A[4][68] [0] = 1'b1;
  assign \A[4][69] [4] = 1'b1;
  assign \A[4][69] [3] = 1'b1;
  assign \A[4][69] [2] = 1'b1;
  assign \A[4][69] [1] = 1'b1;
  assign \A[4][69] [0] = 1'b1;
  assign \A[4][70] [4] = 1'b1;
  assign \A[4][70] [3] = 1'b1;
  assign \A[4][70] [2] = 1'b1;
  assign \A[4][71] [1] = 1'b1;
  assign \A[4][73] [4] = 1'b1;
  assign \A[4][73] [3] = 1'b1;
  assign \A[4][73] [2] = 1'b1;
  assign \A[4][73] [1] = 1'b1;
  assign \A[4][73] [0] = 1'b1;
  assign \A[4][74] [1] = 1'b1;
  assign \A[4][76] [4] = 1'b1;
  assign \A[4][76] [3] = 1'b1;
  assign \A[4][76] [2] = 1'b1;
  assign \A[4][76] [1] = 1'b1;
  assign \A[4][77] [0] = 1'b1;
  assign \A[4][78] [4] = 1'b1;
  assign \A[4][78] [3] = 1'b1;
  assign \A[4][78] [1] = 1'b1;
  assign \A[4][78] [0] = 1'b1;
  assign \A[4][79] [4] = 1'b1;
  assign \A[4][79] [3] = 1'b1;
  assign \A[4][79] [2] = 1'b1;
  assign \A[4][79] [1] = 1'b1;
  assign \A[4][79] [0] = 1'b1;
  assign \A[4][80] [4] = 1'b1;
  assign \A[4][80] [3] = 1'b1;
  assign \A[4][80] [2] = 1'b1;
  assign \A[4][80] [1] = 1'b1;
  assign \A[4][81] [1] = 1'b1;
  assign \A[4][82] [4] = 1'b1;
  assign \A[4][82] [3] = 1'b1;
  assign \A[4][82] [2] = 1'b1;
  assign \A[4][82] [1] = 1'b1;
  assign \A[4][82] [0] = 1'b1;
  assign \A[4][83] [4] = 1'b1;
  assign \A[4][83] [3] = 1'b1;
  assign \A[4][83] [2] = 1'b1;
  assign \A[4][83] [1] = 1'b1;
  assign \A[4][83] [0] = 1'b1;
  assign \A[4][84] [4] = 1'b1;
  assign \A[4][84] [3] = 1'b1;
  assign \A[4][84] [2] = 1'b1;
  assign \A[4][84] [1] = 1'b1;
  assign \A[4][84] [0] = 1'b1;
  assign \A[4][85] [1] = 1'b1;
  assign \A[4][86] [1] = 1'b1;
  assign \A[4][86] [0] = 1'b1;
  assign \A[4][87] [0] = 1'b1;
  assign \A[4][91] [4] = 1'b1;
  assign \A[4][91] [3] = 1'b1;
  assign \A[4][91] [2] = 1'b1;
  assign \A[4][91] [1] = 1'b1;
  assign \A[4][92] [0] = 1'b1;
  assign \A[4][94] [4] = 1'b1;
  assign \A[4][94] [3] = 1'b1;
  assign \A[4][94] [2] = 1'b1;
  assign \A[4][94] [1] = 1'b1;
  assign \A[4][95] [4] = 1'b1;
  assign \A[4][95] [3] = 1'b1;
  assign \A[4][95] [2] = 1'b1;
  assign \A[4][95] [1] = 1'b1;
  assign \A[4][95] [0] = 1'b1;
  assign \A[4][96] [4] = 1'b1;
  assign \A[4][96] [3] = 1'b1;
  assign \A[4][96] [2] = 1'b1;
  assign \A[4][96] [0] = 1'b1;
  assign \A[4][97] [0] = 1'b1;
  assign \A[4][98] [1] = 1'b1;
  assign \A[4][101] [1] = 1'b1;
  assign \A[4][102] [0] = 1'b1;
  assign \A[4][103] [4] = 1'b1;
  assign \A[4][103] [3] = 1'b1;
  assign \A[4][103] [2] = 1'b1;
  assign \A[4][103] [1] = 1'b1;
  assign \A[4][104] [0] = 1'b1;
  assign \A[4][106] [4] = 1'b1;
  assign \A[4][106] [3] = 1'b1;
  assign \A[4][106] [2] = 1'b1;
  assign \A[4][106] [1] = 1'b1;
  assign \A[4][110] [4] = 1'b1;
  assign \A[4][110] [3] = 1'b1;
  assign \A[4][110] [2] = 1'b1;
  assign \A[4][110] [0] = 1'b1;
  assign \A[4][111] [4] = 1'b1;
  assign \A[4][111] [3] = 1'b1;
  assign \A[4][111] [2] = 1'b1;
  assign \A[4][111] [1] = 1'b1;
  assign \A[4][111] [0] = 1'b1;
  assign \A[4][112] [4] = 1'b1;
  assign \A[4][112] [3] = 1'b1;
  assign \A[4][112] [2] = 1'b1;
  assign \A[4][112] [1] = 1'b1;
  assign \A[4][112] [0] = 1'b1;
  assign \A[4][113] [4] = 1'b1;
  assign \A[4][113] [3] = 1'b1;
  assign \A[4][113] [2] = 1'b1;
  assign \A[4][113] [1] = 1'b1;
  assign \A[4][113] [0] = 1'b1;
  assign \A[4][114] [1] = 1'b1;
  assign \A[4][116] [1] = 1'b1;
  assign \A[4][116] [0] = 1'b1;
  assign \A[4][117] [0] = 1'b1;
  assign \A[4][118] [4] = 1'b1;
  assign \A[4][118] [3] = 1'b1;
  assign \A[4][118] [2] = 1'b1;
  assign \A[4][118] [1] = 1'b1;
  assign \A[4][118] [0] = 1'b1;
  assign \A[4][119] [4] = 1'b1;
  assign \A[4][119] [3] = 1'b1;
  assign \A[4][119] [2] = 1'b1;
  assign \A[4][119] [1] = 1'b1;
  assign \A[4][119] [0] = 1'b1;
  assign \A[4][124] [4] = 1'b1;
  assign \A[4][124] [3] = 1'b1;
  assign \A[4][124] [2] = 1'b1;
  assign \A[4][124] [1] = 1'b1;
  assign \A[4][125] [4] = 1'b1;
  assign \A[4][125] [3] = 1'b1;
  assign \A[4][125] [2] = 1'b1;
  assign \A[4][125] [1] = 1'b1;
  assign \A[4][126] [4] = 1'b1;
  assign \A[4][126] [3] = 1'b1;
  assign \A[4][126] [2] = 1'b1;
  assign \A[4][126] [1] = 1'b1;
  assign \A[4][127] [4] = 1'b1;
  assign \A[4][127] [3] = 1'b1;
  assign \A[4][127] [2] = 1'b1;
  assign \A[4][127] [0] = 1'b1;
  assign \A[4][129] [4] = 1'b1;
  assign \A[4][129] [3] = 1'b1;
  assign \A[4][129] [2] = 1'b1;
  assign \A[4][129] [1] = 1'b1;
  assign \A[4][131] [2] = 1'b1;
  assign \A[4][132] [1] = 1'b1;
  assign \A[4][132] [0] = 1'b1;
  assign \A[4][133] [4] = 1'b1;
  assign \A[4][133] [3] = 1'b1;
  assign \A[4][133] [2] = 1'b1;
  assign \A[4][133] [1] = 1'b1;
  assign \A[4][133] [0] = 1'b1;
  assign \A[4][134] [4] = 1'b1;
  assign \A[4][134] [3] = 1'b1;
  assign \A[4][134] [2] = 1'b1;
  assign \A[4][134] [1] = 1'b1;
  assign \A[4][136] [4] = 1'b1;
  assign \A[4][136] [3] = 1'b1;
  assign \A[4][136] [2] = 1'b1;
  assign \A[4][136] [1] = 1'b1;
  assign \A[4][137] [1] = 1'b1;
  assign \A[4][138] [0] = 1'b1;
  assign \A[4][140] [4] = 1'b1;
  assign \A[4][140] [3] = 1'b1;
  assign \A[4][140] [2] = 1'b1;
  assign \A[4][140] [1] = 1'b1;
  assign \A[4][142] [0] = 1'b1;
  assign \A[4][143] [0] = 1'b1;
  assign \A[4][144] [4] = 1'b1;
  assign \A[4][144] [3] = 1'b1;
  assign \A[4][144] [2] = 1'b1;
  assign \A[4][144] [1] = 1'b1;
  assign \A[4][144] [0] = 1'b1;
  assign \A[4][145] [4] = 1'b1;
  assign \A[4][145] [3] = 1'b1;
  assign \A[4][145] [2] = 1'b1;
  assign \A[4][145] [1] = 1'b1;
  assign \A[4][145] [0] = 1'b1;
  assign \A[4][146] [0] = 1'b1;
  assign \A[4][148] [4] = 1'b1;
  assign \A[4][148] [3] = 1'b1;
  assign \A[4][148] [2] = 1'b1;
  assign \A[4][148] [1] = 1'b1;
  assign \A[4][149] [4] = 1'b1;
  assign \A[4][149] [3] = 1'b1;
  assign \A[4][149] [2] = 1'b1;
  assign \A[4][149] [1] = 1'b1;
  assign \A[4][149] [0] = 1'b1;
  assign \A[4][150] [4] = 1'b1;
  assign \A[4][150] [3] = 1'b1;
  assign \A[4][150] [2] = 1'b1;
  assign \A[4][150] [1] = 1'b1;
  assign \A[4][150] [0] = 1'b1;
  assign \A[4][154] [0] = 1'b1;
  assign \A[4][155] [4] = 1'b1;
  assign \A[4][155] [3] = 1'b1;
  assign \A[4][155] [2] = 1'b1;
  assign \A[4][155] [1] = 1'b1;
  assign \A[4][157] [4] = 1'b1;
  assign \A[4][157] [3] = 1'b1;
  assign \A[4][157] [2] = 1'b1;
  assign \A[4][157] [1] = 1'b1;
  assign \A[4][157] [0] = 1'b1;
  assign \A[4][158] [4] = 1'b1;
  assign \A[4][158] [3] = 1'b1;
  assign \A[4][158] [2] = 1'b1;
  assign \A[4][158] [1] = 1'b1;
  assign \A[4][159] [0] = 1'b1;
  assign \A[4][160] [1] = 1'b1;
  assign \A[4][161] [0] = 1'b1;
  assign \A[4][162] [1] = 1'b1;
  assign \A[4][163] [1] = 1'b1;
  assign \A[4][164] [4] = 1'b1;
  assign \A[4][164] [3] = 1'b1;
  assign \A[4][164] [2] = 1'b1;
  assign \A[4][164] [1] = 1'b1;
  assign \A[4][166] [4] = 1'b1;
  assign \A[4][166] [3] = 1'b1;
  assign \A[4][166] [2] = 1'b1;
  assign \A[4][166] [1] = 1'b1;
  assign \A[4][166] [0] = 1'b1;
  assign \A[4][167] [4] = 1'b1;
  assign \A[4][167] [3] = 1'b1;
  assign \A[4][167] [2] = 1'b1;
  assign \A[4][167] [1] = 1'b1;
  assign \A[4][168] [4] = 1'b1;
  assign \A[4][168] [3] = 1'b1;
  assign \A[4][168] [2] = 1'b1;
  assign \A[4][168] [1] = 1'b1;
  assign \A[4][168] [0] = 1'b1;
  assign \A[4][169] [4] = 1'b1;
  assign \A[4][169] [3] = 1'b1;
  assign \A[4][169] [2] = 1'b1;
  assign \A[4][169] [1] = 1'b1;
  assign \A[4][171] [0] = 1'b1;
  assign \A[4][172] [4] = 1'b1;
  assign \A[4][172] [3] = 1'b1;
  assign \A[4][172] [2] = 1'b1;
  assign \A[4][172] [1] = 1'b1;
  assign \A[4][172] [0] = 1'b1;
  assign \A[4][173] [1] = 1'b1;
  assign \A[4][174] [4] = 1'b1;
  assign \A[4][174] [3] = 1'b1;
  assign \A[4][174] [2] = 1'b1;
  assign \A[4][174] [1] = 1'b1;
  assign \A[4][174] [0] = 1'b1;
  assign \A[4][175] [0] = 1'b1;
  assign \A[4][176] [0] = 1'b1;
  assign \A[4][177] [1] = 1'b1;
  assign \A[4][177] [0] = 1'b1;
  assign \A[4][178] [4] = 1'b1;
  assign \A[4][178] [3] = 1'b1;
  assign \A[4][178] [2] = 1'b1;
  assign \A[4][178] [1] = 1'b1;
  assign \A[4][178] [0] = 1'b1;
  assign \A[4][179] [0] = 1'b1;
  assign \A[4][180] [4] = 1'b1;
  assign \A[4][180] [3] = 1'b1;
  assign \A[4][180] [2] = 1'b1;
  assign \A[4][180] [1] = 1'b1;
  assign \A[4][180] [0] = 1'b1;
  assign \A[4][182] [4] = 1'b1;
  assign \A[4][182] [3] = 1'b1;
  assign \A[4][182] [2] = 1'b1;
  assign \A[4][182] [0] = 1'b1;
  assign \A[4][183] [4] = 1'b1;
  assign \A[4][183] [3] = 1'b1;
  assign \A[4][183] [2] = 1'b1;
  assign \A[4][183] [1] = 1'b1;
  assign \A[4][183] [0] = 1'b1;
  assign \A[4][186] [0] = 1'b1;
  assign \A[4][187] [0] = 1'b1;
  assign \A[4][188] [1] = 1'b1;
  assign \A[4][188] [0] = 1'b1;
  assign \A[4][190] [1] = 1'b1;
  assign \A[4][191] [0] = 1'b1;
  assign \A[4][192] [4] = 1'b1;
  assign \A[4][192] [3] = 1'b1;
  assign \A[4][192] [2] = 1'b1;
  assign \A[4][192] [1] = 1'b1;
  assign \A[4][194] [0] = 1'b1;
  assign \A[4][195] [0] = 1'b1;
  assign \A[4][196] [4] = 1'b1;
  assign \A[4][196] [3] = 1'b1;
  assign \A[4][196] [2] = 1'b1;
  assign \A[4][196] [1] = 1'b1;
  assign \A[4][197] [4] = 1'b1;
  assign \A[4][197] [3] = 1'b1;
  assign \A[4][197] [2] = 1'b1;
  assign \A[4][197] [0] = 1'b1;
  assign \A[4][199] [1] = 1'b1;
  assign \A[4][202] [4] = 1'b1;
  assign \A[4][202] [3] = 1'b1;
  assign \A[4][202] [2] = 1'b1;
  assign \A[4][202] [1] = 1'b1;
  assign \A[4][202] [0] = 1'b1;
  assign \A[4][204] [4] = 1'b1;
  assign \A[4][204] [3] = 1'b1;
  assign \A[4][204] [2] = 1'b1;
  assign \A[4][204] [1] = 1'b1;
  assign \A[4][204] [0] = 1'b1;
  assign \A[4][205] [1] = 1'b1;
  assign \A[4][205] [0] = 1'b1;
  assign \A[4][207] [1] = 1'b1;
  assign \A[4][208] [0] = 1'b1;
  assign \A[4][209] [4] = 1'b1;
  assign \A[4][209] [3] = 1'b1;
  assign \A[4][209] [2] = 1'b1;
  assign \A[4][209] [0] = 1'b1;
  assign \A[4][210] [4] = 1'b1;
  assign \A[4][210] [3] = 1'b1;
  assign \A[4][210] [2] = 1'b1;
  assign \A[4][210] [1] = 1'b1;
  assign \A[4][210] [0] = 1'b1;
  assign \A[4][211] [0] = 1'b1;
  assign \A[4][212] [4] = 1'b1;
  assign \A[4][212] [3] = 1'b1;
  assign \A[4][212] [2] = 1'b1;
  assign \A[4][212] [1] = 1'b1;
  assign \A[4][212] [0] = 1'b1;
  assign \A[4][214] [4] = 1'b1;
  assign \A[4][214] [3] = 1'b1;
  assign \A[4][214] [2] = 1'b1;
  assign \A[4][214] [1] = 1'b1;
  assign \A[4][214] [0] = 1'b1;
  assign \A[4][215] [4] = 1'b1;
  assign \A[4][215] [3] = 1'b1;
  assign \A[4][215] [2] = 1'b1;
  assign \A[4][215] [1] = 1'b1;
  assign \A[4][215] [0] = 1'b1;
  assign \A[4][217] [1] = 1'b1;
  assign \A[4][217] [0] = 1'b1;
  assign \A[4][218] [4] = 1'b1;
  assign \A[4][218] [3] = 1'b1;
  assign \A[4][218] [2] = 1'b1;
  assign \A[4][218] [1] = 1'b1;
  assign \A[4][218] [0] = 1'b1;
  assign \A[4][219] [1] = 1'b1;
  assign \A[4][220] [1] = 1'b1;
  assign \A[4][221] [4] = 1'b1;
  assign \A[4][221] [3] = 1'b1;
  assign \A[4][221] [2] = 1'b1;
  assign \A[4][221] [1] = 1'b1;
  assign \A[4][221] [0] = 1'b1;
  assign \A[4][223] [1] = 1'b1;
  assign \A[4][224] [4] = 1'b1;
  assign \A[4][224] [3] = 1'b1;
  assign \A[4][224] [2] = 1'b1;
  assign \A[4][224] [1] = 1'b1;
  assign \A[4][224] [0] = 1'b1;
  assign \A[4][225] [4] = 1'b1;
  assign \A[4][225] [3] = 1'b1;
  assign \A[4][225] [2] = 1'b1;
  assign \A[4][225] [1] = 1'b1;
  assign \A[4][225] [0] = 1'b1;
  assign \A[4][226] [0] = 1'b1;
  assign \A[4][228] [1] = 1'b1;
  assign \A[4][229] [4] = 1'b1;
  assign \A[4][229] [3] = 1'b1;
  assign \A[4][229] [2] = 1'b1;
  assign \A[4][229] [1] = 1'b1;
  assign \A[4][229] [0] = 1'b1;
  assign \A[4][230] [4] = 1'b1;
  assign \A[4][230] [3] = 1'b1;
  assign \A[4][230] [2] = 1'b1;
  assign \A[4][230] [1] = 1'b1;
  assign \A[4][230] [0] = 1'b1;
  assign \A[4][232] [4] = 1'b1;
  assign \A[4][232] [3] = 1'b1;
  assign \A[4][232] [2] = 1'b1;
  assign \A[4][232] [1] = 1'b1;
  assign \A[4][232] [0] = 1'b1;
  assign \A[4][233] [4] = 1'b1;
  assign \A[4][233] [3] = 1'b1;
  assign \A[4][233] [2] = 1'b1;
  assign \A[4][233] [1] = 1'b1;
  assign \A[4][234] [4] = 1'b1;
  assign \A[4][234] [3] = 1'b1;
  assign \A[4][234] [2] = 1'b1;
  assign \A[4][234] [1] = 1'b1;
  assign \A[4][234] [0] = 1'b1;
  assign \A[4][235] [0] = 1'b1;
  assign \A[4][237] [0] = 1'b1;
  assign \A[4][238] [4] = 1'b1;
  assign \A[4][238] [3] = 1'b1;
  assign \A[4][238] [2] = 1'b1;
  assign \A[4][238] [1] = 1'b1;
  assign \A[4][239] [1] = 1'b1;
  assign \A[4][240] [1] = 1'b1;
  assign \A[4][240] [0] = 1'b1;
  assign \A[4][242] [0] = 1'b1;
  assign \A[4][243] [4] = 1'b1;
  assign \A[4][243] [3] = 1'b1;
  assign \A[4][243] [2] = 1'b1;
  assign \A[4][243] [1] = 1'b1;
  assign \A[4][243] [0] = 1'b1;
  assign \A[4][244] [4] = 1'b1;
  assign \A[4][244] [3] = 1'b1;
  assign \A[4][244] [2] = 1'b1;
  assign \A[4][244] [1] = 1'b1;
  assign \A[4][244] [0] = 1'b1;
  assign \A[4][245] [0] = 1'b1;
  assign \A[4][246] [0] = 1'b1;
  assign \A[4][247] [1] = 1'b1;
  assign \A[4][247] [0] = 1'b1;
  assign \A[4][248] [4] = 1'b1;
  assign \A[4][248] [3] = 1'b1;
  assign \A[4][248] [2] = 1'b1;
  assign \A[4][248] [1] = 1'b1;
  assign \A[4][248] [0] = 1'b1;
  assign \A[4][249] [4] = 1'b1;
  assign \A[4][249] [3] = 1'b1;
  assign \A[4][249] [2] = 1'b1;
  assign \A[4][249] [1] = 1'b1;
  assign \A[4][249] [0] = 1'b1;
  assign \A[4][251] [0] = 1'b1;
  assign \A[4][252] [0] = 1'b1;
  assign \A[4][253] [0] = 1'b1;
  assign \A[4][254] [4] = 1'b1;
  assign \A[4][254] [3] = 1'b1;
  assign \A[4][254] [2] = 1'b1;
  assign \A[4][254] [1] = 1'b1;
  assign \A[4][254] [0] = 1'b1;
  assign \A[4][255] [0] = 1'b1;
  assign \A[5][0] [4] = 1'b1;
  assign \A[5][0] [3] = 1'b1;
  assign \A[5][0] [2] = 1'b1;
  assign \A[5][0] [1] = 1'b1;
  assign \A[5][2] [4] = 1'b1;
  assign \A[5][2] [3] = 1'b1;
  assign \A[5][2] [2] = 1'b1;
  assign \A[5][2] [1] = 1'b1;
  assign \A[5][2] [0] = 1'b1;
  assign \A[5][3] [4] = 1'b1;
  assign \A[5][3] [3] = 1'b1;
  assign \A[5][3] [2] = 1'b1;
  assign \A[5][3] [1] = 1'b1;
  assign \A[5][3] [0] = 1'b1;
  assign \A[5][5] [4] = 1'b1;
  assign \A[5][5] [3] = 1'b1;
  assign \A[5][5] [2] = 1'b1;
  assign \A[5][5] [1] = 1'b1;
  assign \A[5][5] [0] = 1'b1;
  assign \A[5][6] [4] = 1'b1;
  assign \A[5][6] [3] = 1'b1;
  assign \A[5][6] [2] = 1'b1;
  assign \A[5][6] [1] = 1'b1;
  assign \A[5][6] [0] = 1'b1;
  assign \A[5][7] [4] = 1'b1;
  assign \A[5][7] [3] = 1'b1;
  assign \A[5][7] [2] = 1'b1;
  assign \A[5][7] [1] = 1'b1;
  assign \A[5][7] [0] = 1'b1;
  assign \A[5][8] [4] = 1'b1;
  assign \A[5][8] [3] = 1'b1;
  assign \A[5][8] [2] = 1'b1;
  assign \A[5][8] [1] = 1'b1;
  assign \A[5][8] [0] = 1'b1;
  assign \A[5][10] [4] = 1'b1;
  assign \A[5][10] [3] = 1'b1;
  assign \A[5][10] [2] = 1'b1;
  assign \A[5][10] [1] = 1'b1;
  assign \A[5][10] [0] = 1'b1;
  assign \A[5][11] [4] = 1'b1;
  assign \A[5][11] [3] = 1'b1;
  assign \A[5][11] [2] = 1'b1;
  assign \A[5][11] [1] = 1'b1;
  assign \A[5][11] [0] = 1'b1;
  assign \A[5][12] [4] = 1'b1;
  assign \A[5][12] [3] = 1'b1;
  assign \A[5][12] [2] = 1'b1;
  assign \A[5][12] [0] = 1'b1;
  assign \A[5][13] [4] = 1'b1;
  assign \A[5][13] [3] = 1'b1;
  assign \A[5][13] [2] = 1'b1;
  assign \A[5][13] [0] = 1'b1;
  assign \A[5][14] [4] = 1'b1;
  assign \A[5][14] [3] = 1'b1;
  assign \A[5][14] [2] = 1'b1;
  assign \A[5][14] [1] = 1'b1;
  assign \A[5][14] [0] = 1'b1;
  assign \A[5][15] [4] = 1'b1;
  assign \A[5][15] [3] = 1'b1;
  assign \A[5][15] [2] = 1'b1;
  assign \A[5][15] [1] = 1'b1;
  assign \A[5][16] [4] = 1'b1;
  assign \A[5][16] [3] = 1'b1;
  assign \A[5][16] [2] = 1'b1;
  assign \A[5][16] [1] = 1'b1;
  assign \A[5][16] [0] = 1'b1;
  assign \A[5][17] [0] = 1'b1;
  assign \A[5][18] [4] = 1'b1;
  assign \A[5][18] [3] = 1'b1;
  assign \A[5][18] [2] = 1'b1;
  assign \A[5][18] [1] = 1'b1;
  assign \A[5][18] [0] = 1'b1;
  assign \A[5][19] [1] = 1'b1;
  assign \A[5][20] [0] = 1'b1;
  assign \A[5][22] [1] = 1'b1;
  assign \A[5][23] [4] = 1'b1;
  assign \A[5][23] [3] = 1'b1;
  assign \A[5][23] [2] = 1'b1;
  assign \A[5][23] [1] = 1'b1;
  assign \A[5][23] [0] = 1'b1;
  assign \A[5][24] [4] = 1'b1;
  assign \A[5][24] [3] = 1'b1;
  assign \A[5][24] [2] = 1'b1;
  assign \A[5][24] [1] = 1'b1;
  assign \A[5][25] [4] = 1'b1;
  assign \A[5][25] [3] = 1'b1;
  assign \A[5][25] [2] = 1'b1;
  assign \A[5][25] [1] = 1'b1;
  assign \A[5][25] [0] = 1'b1;
  assign \A[5][26] [4] = 1'b1;
  assign \A[5][26] [3] = 1'b1;
  assign \A[5][26] [2] = 1'b1;
  assign \A[5][26] [1] = 1'b1;
  assign \A[5][26] [0] = 1'b1;
  assign \A[5][29] [4] = 1'b1;
  assign \A[5][29] [3] = 1'b1;
  assign \A[5][29] [2] = 1'b1;
  assign \A[5][29] [1] = 1'b1;
  assign \A[5][29] [0] = 1'b1;
  assign \A[5][30] [4] = 1'b1;
  assign \A[5][30] [3] = 1'b1;
  assign \A[5][30] [2] = 1'b1;
  assign \A[5][30] [1] = 1'b1;
  assign \A[5][30] [0] = 1'b1;
  assign \A[5][31] [4] = 1'b1;
  assign \A[5][31] [3] = 1'b1;
  assign \A[5][31] [2] = 1'b1;
  assign \A[5][31] [1] = 1'b1;
  assign \A[5][31] [0] = 1'b1;
  assign \A[5][34] [4] = 1'b1;
  assign \A[5][34] [3] = 1'b1;
  assign \A[5][34] [2] = 1'b1;
  assign \A[5][34] [1] = 1'b1;
  assign \A[5][34] [0] = 1'b1;
  assign \A[5][35] [0] = 1'b1;
  assign \A[5][37] [0] = 1'b1;
  assign \A[5][38] [1] = 1'b1;
  assign \A[5][39] [1] = 1'b1;
  assign \A[5][39] [0] = 1'b1;
  assign \A[5][40] [4] = 1'b1;
  assign \A[5][40] [3] = 1'b1;
  assign \A[5][40] [2] = 1'b1;
  assign \A[5][40] [1] = 1'b1;
  assign \A[5][40] [0] = 1'b1;
  assign \A[5][41] [4] = 1'b1;
  assign \A[5][41] [3] = 1'b1;
  assign \A[5][41] [2] = 1'b1;
  assign \A[5][41] [1] = 1'b1;
  assign \A[5][42] [4] = 1'b1;
  assign \A[5][42] [3] = 1'b1;
  assign \A[5][42] [1] = 1'b1;
  assign \A[5][42] [0] = 1'b1;
  assign \A[5][43] [4] = 1'b1;
  assign \A[5][43] [3] = 1'b1;
  assign \A[5][43] [2] = 1'b1;
  assign \A[5][43] [1] = 1'b1;
  assign \A[5][44] [4] = 1'b1;
  assign \A[5][44] [3] = 1'b1;
  assign \A[5][44] [2] = 1'b1;
  assign \A[5][44] [0] = 1'b1;
  assign \A[5][45] [4] = 1'b1;
  assign \A[5][45] [3] = 1'b1;
  assign \A[5][45] [2] = 1'b1;
  assign \A[5][45] [1] = 1'b1;
  assign \A[5][49] [4] = 1'b1;
  assign \A[5][49] [3] = 1'b1;
  assign \A[5][49] [2] = 1'b1;
  assign \A[5][49] [1] = 1'b1;
  assign \A[5][49] [0] = 1'b1;
  assign \A[5][50] [4] = 1'b1;
  assign \A[5][50] [3] = 1'b1;
  assign \A[5][50] [2] = 1'b1;
  assign \A[5][50] [1] = 1'b1;
  assign \A[5][50] [0] = 1'b1;
  assign \A[5][51] [1] = 1'b1;
  assign \A[5][52] [4] = 1'b1;
  assign \A[5][52] [3] = 1'b1;
  assign \A[5][52] [2] = 1'b1;
  assign \A[5][52] [1] = 1'b1;
  assign \A[5][52] [0] = 1'b1;
  assign \A[5][53] [0] = 1'b1;
  assign \A[5][54] [1] = 1'b1;
  assign \A[5][58] [4] = 1'b1;
  assign \A[5][58] [3] = 1'b1;
  assign \A[5][58] [2] = 1'b1;
  assign \A[5][58] [1] = 1'b1;
  assign \A[5][58] [0] = 1'b1;
  assign \A[5][59] [4] = 1'b1;
  assign \A[5][59] [3] = 1'b1;
  assign \A[5][59] [2] = 1'b1;
  assign \A[5][59] [1] = 1'b1;
  assign \A[5][59] [0] = 1'b1;
  assign \A[5][60] [4] = 1'b1;
  assign \A[5][60] [3] = 1'b1;
  assign \A[5][60] [2] = 1'b1;
  assign \A[5][60] [1] = 1'b1;
  assign \A[5][62] [0] = 1'b1;
  assign \A[5][63] [1] = 1'b1;
  assign \A[5][64] [1] = 1'b1;
  assign \A[5][65] [4] = 1'b1;
  assign \A[5][65] [3] = 1'b1;
  assign \A[5][65] [2] = 1'b1;
  assign \A[5][65] [1] = 1'b1;
  assign \A[5][65] [0] = 1'b1;
  assign \A[5][67] [0] = 1'b1;
  assign \A[5][68] [0] = 1'b1;
  assign \A[5][69] [0] = 1'b1;
  assign \A[5][70] [1] = 1'b1;
  assign \A[5][70] [0] = 1'b1;
  assign \A[5][71] [4] = 1'b1;
  assign \A[5][71] [3] = 1'b1;
  assign \A[5][71] [2] = 1'b1;
  assign \A[5][71] [1] = 1'b1;
  assign \A[5][72] [4] = 1'b1;
  assign \A[5][72] [3] = 1'b1;
  assign \A[5][72] [2] = 1'b1;
  assign \A[5][72] [1] = 1'b1;
  assign \A[5][72] [0] = 1'b1;
  assign \A[5][73] [4] = 1'b1;
  assign \A[5][73] [3] = 1'b1;
  assign \A[5][73] [2] = 1'b1;
  assign \A[5][73] [1] = 1'b1;
  assign \A[5][74] [1] = 1'b1;
  assign \A[5][74] [0] = 1'b1;
  assign \A[5][75] [4] = 1'b1;
  assign \A[5][75] [3] = 1'b1;
  assign \A[5][75] [2] = 1'b1;
  assign \A[5][75] [1] = 1'b1;
  assign \A[5][75] [0] = 1'b1;
  assign \A[5][76] [4] = 1'b1;
  assign \A[5][76] [3] = 1'b1;
  assign \A[5][76] [2] = 1'b1;
  assign \A[5][76] [1] = 1'b1;
  assign \A[5][76] [0] = 1'b1;
  assign \A[5][78] [4] = 1'b1;
  assign \A[5][78] [3] = 1'b1;
  assign \A[5][78] [2] = 1'b1;
  assign \A[5][78] [1] = 1'b1;
  assign \A[5][78] [0] = 1'b1;
  assign \A[5][82] [4] = 1'b1;
  assign \A[5][82] [3] = 1'b1;
  assign \A[5][82] [2] = 1'b1;
  assign \A[5][82] [1] = 1'b1;
  assign \A[5][83] [4] = 1'b1;
  assign \A[5][83] [3] = 1'b1;
  assign \A[5][83] [2] = 1'b1;
  assign \A[5][83] [1] = 1'b1;
  assign \A[5][83] [0] = 1'b1;
  assign \A[5][84] [1] = 1'b1;
  assign \A[5][85] [0] = 1'b1;
  assign \A[5][86] [0] = 1'b1;
  assign \A[5][87] [0] = 1'b1;
  assign \A[5][88] [0] = 1'b1;
  assign \A[5][89] [4] = 1'b1;
  assign \A[5][89] [3] = 1'b1;
  assign \A[5][89] [2] = 1'b1;
  assign \A[5][89] [1] = 1'b1;
  assign \A[5][90] [4] = 1'b1;
  assign \A[5][90] [3] = 1'b1;
  assign \A[5][90] [2] = 1'b1;
  assign \A[5][90] [1] = 1'b1;
  assign \A[5][91] [4] = 1'b1;
  assign \A[5][91] [3] = 1'b1;
  assign \A[5][91] [2] = 1'b1;
  assign \A[5][91] [1] = 1'b1;
  assign \A[5][92] [0] = 1'b1;
  assign \A[5][95] [4] = 1'b1;
  assign \A[5][95] [3] = 1'b1;
  assign \A[5][95] [2] = 1'b1;
  assign \A[5][95] [1] = 1'b1;
  assign \A[5][95] [0] = 1'b1;
  assign \A[5][96] [0] = 1'b1;
  assign \A[5][98] [4] = 1'b1;
  assign \A[5][98] [3] = 1'b1;
  assign \A[5][98] [2] = 1'b1;
  assign \A[5][98] [1] = 1'b1;
  assign \A[5][98] [0] = 1'b1;
  assign \A[5][99] [1] = 1'b1;
  assign \A[5][99] [0] = 1'b1;
  assign \A[5][100] [0] = 1'b1;
  assign \A[5][101] [4] = 1'b1;
  assign \A[5][101] [3] = 1'b1;
  assign \A[5][101] [2] = 1'b1;
  assign \A[5][101] [1] = 1'b1;
  assign \A[5][101] [0] = 1'b1;
  assign \A[5][102] [0] = 1'b1;
  assign \A[5][103] [1] = 1'b1;
  assign \A[5][107] [4] = 1'b1;
  assign \A[5][107] [3] = 1'b1;
  assign \A[5][107] [2] = 1'b1;
  assign \A[5][107] [1] = 1'b1;
  assign \A[5][108] [4] = 1'b1;
  assign \A[5][108] [3] = 1'b1;
  assign \A[5][108] [2] = 1'b1;
  assign \A[5][108] [0] = 1'b1;
  assign \A[5][110] [1] = 1'b1;
  assign \A[5][110] [0] = 1'b1;
  assign \A[5][111] [0] = 1'b1;
  assign \A[5][113] [4] = 1'b1;
  assign \A[5][113] [3] = 1'b1;
  assign \A[5][113] [2] = 1'b1;
  assign \A[5][113] [1] = 1'b1;
  assign \A[5][113] [0] = 1'b1;
  assign \A[5][114] [1] = 1'b1;
  assign \A[5][118] [1] = 1'b1;
  assign \A[5][118] [0] = 1'b1;
  assign \A[5][120] [4] = 1'b1;
  assign \A[5][120] [3] = 1'b1;
  assign \A[5][120] [2] = 1'b1;
  assign \A[5][120] [1] = 1'b1;
  assign \A[5][120] [0] = 1'b1;
  assign \A[5][121] [4] = 1'b1;
  assign \A[5][121] [3] = 1'b1;
  assign \A[5][121] [2] = 1'b1;
  assign \A[5][121] [0] = 1'b1;
  assign \A[5][124] [4] = 1'b1;
  assign \A[5][124] [3] = 1'b1;
  assign \A[5][124] [2] = 1'b1;
  assign \A[5][124] [1] = 1'b1;
  assign \A[5][125] [4] = 1'b1;
  assign \A[5][125] [3] = 1'b1;
  assign \A[5][125] [2] = 1'b1;
  assign \A[5][125] [1] = 1'b1;
  assign \A[5][125] [0] = 1'b1;
  assign \A[5][126] [4] = 1'b1;
  assign \A[5][126] [3] = 1'b1;
  assign \A[5][126] [2] = 1'b1;
  assign \A[5][126] [1] = 1'b1;
  assign \A[5][126] [0] = 1'b1;
  assign \A[5][127] [4] = 1'b1;
  assign \A[5][127] [3] = 1'b1;
  assign \A[5][127] [2] = 1'b1;
  assign \A[5][127] [1] = 1'b1;
  assign \A[5][127] [0] = 1'b1;
  assign \A[5][128] [0] = 1'b1;
  assign \A[5][129] [4] = 1'b1;
  assign \A[5][129] [3] = 1'b1;
  assign \A[5][129] [2] = 1'b1;
  assign \A[5][129] [1] = 1'b1;
  assign \A[5][129] [0] = 1'b1;
  assign \A[5][130] [1] = 1'b1;
  assign \A[5][132] [0] = 1'b1;
  assign \A[5][133] [4] = 1'b1;
  assign \A[5][133] [3] = 1'b1;
  assign \A[5][133] [2] = 1'b1;
  assign \A[5][133] [1] = 1'b1;
  assign \A[5][133] [0] = 1'b1;
  assign \A[5][134] [0] = 1'b1;
  assign \A[5][137] [4] = 1'b1;
  assign \A[5][137] [3] = 1'b1;
  assign \A[5][137] [2] = 1'b1;
  assign \A[5][137] [1] = 1'b1;
  assign \A[5][139] [4] = 1'b1;
  assign \A[5][139] [3] = 1'b1;
  assign \A[5][139] [2] = 1'b1;
  assign \A[5][139] [1] = 1'b1;
  assign \A[5][140] [4] = 1'b1;
  assign \A[5][140] [3] = 1'b1;
  assign \A[5][140] [2] = 1'b1;
  assign \A[5][140] [0] = 1'b1;
  assign \A[5][141] [4] = 1'b1;
  assign \A[5][141] [3] = 1'b1;
  assign \A[5][141] [2] = 1'b1;
  assign \A[5][141] [1] = 1'b1;
  assign \A[5][142] [4] = 1'b1;
  assign \A[5][142] [3] = 1'b1;
  assign \A[5][142] [2] = 1'b1;
  assign \A[5][142] [1] = 1'b1;
  assign \A[5][143] [0] = 1'b1;
  assign \A[5][144] [4] = 1'b1;
  assign \A[5][144] [3] = 1'b1;
  assign \A[5][144] [2] = 1'b1;
  assign \A[5][146] [4] = 1'b1;
  assign \A[5][146] [3] = 1'b1;
  assign \A[5][146] [2] = 1'b1;
  assign \A[5][146] [0] = 1'b1;
  assign \A[5][147] [4] = 1'b1;
  assign \A[5][147] [3] = 1'b1;
  assign \A[5][147] [2] = 1'b1;
  assign \A[5][147] [1] = 1'b1;
  assign \A[5][147] [0] = 1'b1;
  assign \A[5][149] [1] = 1'b1;
  assign \A[5][151] [0] = 1'b1;
  assign \A[5][152] [4] = 1'b1;
  assign \A[5][152] [3] = 1'b1;
  assign \A[5][152] [2] = 1'b1;
  assign \A[5][152] [0] = 1'b1;
  assign \A[5][153] [0] = 1'b1;
  assign \A[5][154] [4] = 1'b1;
  assign \A[5][154] [3] = 1'b1;
  assign \A[5][154] [2] = 1'b1;
  assign \A[5][154] [0] = 1'b1;
  assign \A[5][155] [4] = 1'b1;
  assign \A[5][155] [3] = 1'b1;
  assign \A[5][155] [2] = 1'b1;
  assign \A[5][155] [1] = 1'b1;
  assign \A[5][156] [4] = 1'b1;
  assign \A[5][156] [3] = 1'b1;
  assign \A[5][156] [2] = 1'b1;
  assign \A[5][156] [1] = 1'b1;
  assign \A[5][156] [0] = 1'b1;
  assign \A[5][157] [4] = 1'b1;
  assign \A[5][157] [3] = 1'b1;
  assign \A[5][157] [2] = 1'b1;
  assign \A[5][157] [1] = 1'b1;
  assign \A[5][157] [0] = 1'b1;
  assign \A[5][159] [4] = 1'b1;
  assign \A[5][159] [3] = 1'b1;
  assign \A[5][159] [2] = 1'b1;
  assign \A[5][159] [1] = 1'b1;
  assign \A[5][159] [0] = 1'b1;
  assign \A[5][160] [4] = 1'b1;
  assign \A[5][160] [3] = 1'b1;
  assign \A[5][160] [2] = 1'b1;
  assign \A[5][160] [1] = 1'b1;
  assign \A[5][161] [4] = 1'b1;
  assign \A[5][161] [3] = 1'b1;
  assign \A[5][161] [2] = 1'b1;
  assign \A[5][161] [1] = 1'b1;
  assign \A[5][161] [0] = 1'b1;
  assign \A[5][162] [4] = 1'b1;
  assign \A[5][162] [3] = 1'b1;
  assign \A[5][162] [2] = 1'b1;
  assign \A[5][162] [1] = 1'b1;
  assign \A[5][163] [4] = 1'b1;
  assign \A[5][163] [3] = 1'b1;
  assign \A[5][163] [2] = 1'b1;
  assign \A[5][163] [1] = 1'b1;
  assign \A[5][163] [0] = 1'b1;
  assign \A[5][165] [0] = 1'b1;
  assign \A[5][166] [1] = 1'b1;
  assign \A[5][167] [4] = 1'b1;
  assign \A[5][167] [3] = 1'b1;
  assign \A[5][167] [2] = 1'b1;
  assign \A[5][167] [1] = 1'b1;
  assign \A[5][169] [1] = 1'b1;
  assign \A[5][169] [0] = 1'b1;
  assign \A[5][170] [4] = 1'b1;
  assign \A[5][170] [3] = 1'b1;
  assign \A[5][170] [2] = 1'b1;
  assign \A[5][170] [1] = 1'b1;
  assign \A[5][170] [0] = 1'b1;
  assign \A[5][171] [4] = 1'b1;
  assign \A[5][171] [3] = 1'b1;
  assign \A[5][171] [2] = 1'b1;
  assign \A[5][171] [1] = 1'b1;
  assign \A[5][171] [0] = 1'b1;
  assign \A[5][173] [0] = 1'b1;
  assign \A[5][174] [4] = 1'b1;
  assign \A[5][174] [3] = 1'b1;
  assign \A[5][174] [2] = 1'b1;
  assign \A[5][174] [1] = 1'b1;
  assign \A[5][174] [0] = 1'b1;
  assign \A[5][175] [4] = 1'b1;
  assign \A[5][175] [3] = 1'b1;
  assign \A[5][175] [2] = 1'b1;
  assign \A[5][175] [0] = 1'b1;
  assign \A[5][176] [4] = 1'b1;
  assign \A[5][176] [3] = 1'b1;
  assign \A[5][176] [2] = 1'b1;
  assign \A[5][176] [1] = 1'b1;
  assign \A[5][176] [0] = 1'b1;
  assign \A[5][177] [4] = 1'b1;
  assign \A[5][177] [3] = 1'b1;
  assign \A[5][177] [2] = 1'b1;
  assign \A[5][177] [1] = 1'b1;
  assign \A[5][178] [0] = 1'b1;
  assign \A[5][179] [0] = 1'b1;
  assign \A[5][180] [4] = 1'b1;
  assign \A[5][180] [3] = 1'b1;
  assign \A[5][180] [2] = 1'b1;
  assign \A[5][180] [1] = 1'b1;
  assign \A[5][181] [1] = 1'b1;
  assign \A[5][182] [1] = 1'b1;
  assign \A[5][183] [0] = 1'b1;
  assign \A[5][184] [4] = 1'b1;
  assign \A[5][184] [3] = 1'b1;
  assign \A[5][184] [2] = 1'b1;
  assign \A[5][184] [1] = 1'b1;
  assign \A[5][184] [0] = 1'b1;
  assign \A[5][185] [0] = 1'b1;
  assign \A[5][187] [1] = 1'b1;
  assign \A[5][188] [0] = 1'b1;
  assign \A[5][189] [1] = 1'b1;
  assign \A[5][190] [0] = 1'b1;
  assign \A[5][191] [4] = 1'b1;
  assign \A[5][191] [3] = 1'b1;
  assign \A[5][191] [2] = 1'b1;
  assign \A[5][191] [0] = 1'b1;
  assign \A[5][192] [4] = 1'b1;
  assign \A[5][192] [3] = 1'b1;
  assign \A[5][192] [2] = 1'b1;
  assign \A[5][193] [0] = 1'b1;
  assign \A[5][196] [1] = 1'b1;
  assign \A[5][196] [0] = 1'b1;
  assign \A[5][197] [0] = 1'b1;
  assign \A[5][198] [0] = 1'b1;
  assign \A[5][200] [0] = 1'b1;
  assign \A[5][201] [0] = 1'b1;
  assign \A[5][202] [4] = 1'b1;
  assign \A[5][202] [3] = 1'b1;
  assign \A[5][202] [2] = 1'b1;
  assign \A[5][202] [1] = 1'b1;
  assign \A[5][203] [0] = 1'b1;
  assign \A[5][205] [4] = 1'b1;
  assign \A[5][205] [3] = 1'b1;
  assign \A[5][205] [2] = 1'b1;
  assign \A[5][205] [1] = 1'b1;
  assign \A[5][205] [0] = 1'b1;
  assign \A[5][206] [4] = 1'b1;
  assign \A[5][206] [3] = 1'b1;
  assign \A[5][206] [2] = 1'b1;
  assign \A[5][206] [1] = 1'b1;
  assign \A[5][208] [4] = 1'b1;
  assign \A[5][208] [3] = 1'b1;
  assign \A[5][208] [2] = 1'b1;
  assign \A[5][208] [1] = 1'b1;
  assign \A[5][208] [0] = 1'b1;
  assign \A[5][209] [4] = 1'b1;
  assign \A[5][209] [3] = 1'b1;
  assign \A[5][209] [2] = 1'b1;
  assign \A[5][209] [1] = 1'b1;
  assign \A[5][210] [4] = 1'b1;
  assign \A[5][210] [3] = 1'b1;
  assign \A[5][210] [2] = 1'b1;
  assign \A[5][210] [1] = 1'b1;
  assign \A[5][212] [2] = 1'b1;
  assign \A[5][214] [4] = 1'b1;
  assign \A[5][214] [3] = 1'b1;
  assign \A[5][214] [2] = 1'b1;
  assign \A[5][214] [1] = 1'b1;
  assign \A[5][214] [0] = 1'b1;
  assign \A[5][215] [0] = 1'b1;
  assign \A[5][216] [4] = 1'b1;
  assign \A[5][216] [3] = 1'b1;
  assign \A[5][216] [2] = 1'b1;
  assign \A[5][216] [1] = 1'b1;
  assign \A[5][217] [0] = 1'b1;
  assign \A[5][219] [1] = 1'b1;
  assign \A[5][221] [4] = 1'b1;
  assign \A[5][221] [3] = 1'b1;
  assign \A[5][221] [2] = 1'b1;
  assign \A[5][221] [1] = 1'b1;
  assign \A[5][222] [0] = 1'b1;
  assign \A[5][223] [4] = 1'b1;
  assign \A[5][223] [3] = 1'b1;
  assign \A[5][223] [2] = 1'b1;
  assign \A[5][223] [1] = 1'b1;
  assign \A[5][224] [0] = 1'b1;
  assign \A[5][225] [0] = 1'b1;
  assign \A[5][226] [4] = 1'b1;
  assign \A[5][226] [3] = 1'b1;
  assign \A[5][226] [2] = 1'b1;
  assign \A[5][226] [1] = 1'b1;
  assign \A[5][226] [0] = 1'b1;
  assign \A[5][227] [4] = 1'b1;
  assign \A[5][227] [3] = 1'b1;
  assign \A[5][227] [2] = 1'b1;
  assign \A[5][227] [1] = 1'b1;
  assign \A[5][227] [0] = 1'b1;
  assign \A[5][228] [4] = 1'b1;
  assign \A[5][228] [3] = 1'b1;
  assign \A[5][228] [2] = 1'b1;
  assign \A[5][228] [1] = 1'b1;
  assign \A[5][228] [0] = 1'b1;
  assign \A[5][230] [4] = 1'b1;
  assign \A[5][230] [3] = 1'b1;
  assign \A[5][230] [2] = 1'b1;
  assign \A[5][230] [1] = 1'b1;
  assign \A[5][230] [0] = 1'b1;
  assign \A[5][231] [4] = 1'b1;
  assign \A[5][231] [3] = 1'b1;
  assign \A[5][231] [2] = 1'b1;
  assign \A[5][231] [1] = 1'b1;
  assign \A[5][231] [0] = 1'b1;
  assign \A[5][232] [0] = 1'b1;
  assign \A[5][233] [1] = 1'b1;
  assign \A[5][233] [0] = 1'b1;
  assign \A[5][234] [1] = 1'b1;
  assign \A[5][235] [4] = 1'b1;
  assign \A[5][235] [3] = 1'b1;
  assign \A[5][235] [2] = 1'b1;
  assign \A[5][235] [1] = 1'b1;
  assign \A[5][236] [4] = 1'b1;
  assign \A[5][236] [3] = 1'b1;
  assign \A[5][236] [2] = 1'b1;
  assign \A[5][236] [1] = 1'b1;
  assign \A[5][237] [4] = 1'b1;
  assign \A[5][237] [3] = 1'b1;
  assign \A[5][237] [2] = 1'b1;
  assign \A[5][237] [0] = 1'b1;
  assign \A[5][238] [4] = 1'b1;
  assign \A[5][238] [3] = 1'b1;
  assign \A[5][238] [2] = 1'b1;
  assign \A[5][238] [1] = 1'b1;
  assign \A[5][238] [0] = 1'b1;
  assign \A[5][240] [4] = 1'b1;
  assign \A[5][240] [3] = 1'b1;
  assign \A[5][240] [2] = 1'b1;
  assign \A[5][240] [0] = 1'b1;
  assign \A[5][241] [4] = 1'b1;
  assign \A[5][241] [3] = 1'b1;
  assign \A[5][241] [2] = 1'b1;
  assign \A[5][241] [1] = 1'b1;
  assign \A[5][242] [4] = 1'b1;
  assign \A[5][242] [3] = 1'b1;
  assign \A[5][242] [2] = 1'b1;
  assign \A[5][242] [1] = 1'b1;
  assign \A[5][243] [4] = 1'b1;
  assign \A[5][243] [3] = 1'b1;
  assign \A[5][243] [2] = 1'b1;
  assign \A[5][243] [1] = 1'b1;
  assign \A[5][244] [0] = 1'b1;
  assign \A[5][245] [4] = 1'b1;
  assign \A[5][245] [3] = 1'b1;
  assign \A[5][245] [2] = 1'b1;
  assign \A[5][245] [1] = 1'b1;
  assign \A[5][245] [0] = 1'b1;
  assign \A[5][246] [0] = 1'b1;
  assign \A[5][248] [4] = 1'b1;
  assign \A[5][248] [3] = 1'b1;
  assign \A[5][248] [2] = 1'b1;
  assign \A[5][248] [1] = 1'b1;
  assign \A[5][248] [0] = 1'b1;
  assign \A[5][250] [0] = 1'b1;
  assign \A[5][251] [0] = 1'b1;
  assign \A[5][252] [0] = 1'b1;
  assign \A[5][254] [4] = 1'b1;
  assign \A[5][254] [3] = 1'b1;
  assign \A[5][254] [2] = 1'b1;
  assign \A[5][254] [1] = 1'b1;
  assign \A[5][254] [0] = 1'b1;
  assign \A[5][255] [4] = 1'b1;
  assign \A[5][255] [3] = 1'b1;
  assign \A[5][255] [2] = 1'b1;
  assign \A[5][255] [1] = 1'b1;
  assign \A[5][255] [0] = 1'b1;
  assign \A[6][0] [1] = 1'b1;
  assign \A[6][1] [0] = 1'b1;
  assign \A[6][2] [4] = 1'b1;
  assign \A[6][2] [3] = 1'b1;
  assign \A[6][2] [2] = 1'b1;
  assign \A[6][2] [1] = 1'b1;
  assign \A[6][2] [0] = 1'b1;
  assign \A[6][7] [4] = 1'b1;
  assign \A[6][7] [3] = 1'b1;
  assign \A[6][7] [2] = 1'b1;
  assign \A[6][7] [0] = 1'b1;
  assign \A[6][8] [1] = 1'b1;
  assign \A[6][8] [0] = 1'b1;
  assign \A[6][9] [0] = 1'b1;
  assign \A[6][10] [1] = 1'b1;
  assign \A[6][10] [0] = 1'b1;
  assign \A[6][11] [1] = 1'b1;
  assign \A[6][11] [0] = 1'b1;
  assign \A[6][12] [1] = 1'b1;
  assign \A[6][13] [4] = 1'b1;
  assign \A[6][13] [3] = 1'b1;
  assign \A[6][13] [2] = 1'b1;
  assign \A[6][13] [1] = 1'b1;
  assign \A[6][14] [4] = 1'b1;
  assign \A[6][14] [3] = 1'b1;
  assign \A[6][14] [2] = 1'b1;
  assign \A[6][14] [1] = 1'b1;
  assign \A[6][15] [4] = 1'b1;
  assign \A[6][15] [3] = 1'b1;
  assign \A[6][15] [2] = 1'b1;
  assign \A[6][15] [1] = 1'b1;
  assign \A[6][16] [4] = 1'b1;
  assign \A[6][16] [3] = 1'b1;
  assign \A[6][16] [2] = 1'b1;
  assign \A[6][16] [1] = 1'b1;
  assign \A[6][16] [0] = 1'b1;
  assign \A[6][17] [0] = 1'b1;
  assign \A[6][21] [0] = 1'b1;
  assign \A[6][23] [1] = 1'b1;
  assign \A[6][24] [0] = 1'b1;
  assign \A[6][25] [4] = 1'b1;
  assign \A[6][25] [3] = 1'b1;
  assign \A[6][25] [2] = 1'b1;
  assign \A[6][25] [1] = 1'b1;
  assign \A[6][26] [2] = 1'b1;
  assign \A[6][28] [4] = 1'b1;
  assign \A[6][28] [3] = 1'b1;
  assign \A[6][28] [2] = 1'b1;
  assign \A[6][28] [0] = 1'b1;
  assign \A[6][30] [4] = 1'b1;
  assign \A[6][30] [3] = 1'b1;
  assign \A[6][30] [2] = 1'b1;
  assign \A[6][30] [1] = 1'b1;
  assign \A[6][30] [0] = 1'b1;
  assign \A[6][31] [0] = 1'b1;
  assign \A[6][32] [4] = 1'b1;
  assign \A[6][32] [3] = 1'b1;
  assign \A[6][32] [2] = 1'b1;
  assign \A[6][32] [1] = 1'b1;
  assign \A[6][32] [0] = 1'b1;
  assign \A[6][33] [1] = 1'b1;
  assign \A[6][34] [0] = 1'b1;
  assign \A[6][35] [0] = 1'b1;
  assign \A[6][37] [0] = 1'b1;
  assign \A[6][40] [0] = 1'b1;
  assign \A[6][41] [4] = 1'b1;
  assign \A[6][41] [3] = 1'b1;
  assign \A[6][41] [2] = 1'b1;
  assign \A[6][41] [0] = 1'b1;
  assign \A[6][43] [0] = 1'b1;
  assign \A[6][45] [4] = 1'b1;
  assign \A[6][45] [3] = 1'b1;
  assign \A[6][45] [2] = 1'b1;
  assign \A[6][45] [1] = 1'b1;
  assign \A[6][45] [0] = 1'b1;
  assign \A[6][46] [1] = 1'b1;
  assign \A[6][46] [0] = 1'b1;
  assign \A[6][47] [4] = 1'b1;
  assign \A[6][47] [3] = 1'b1;
  assign \A[6][47] [2] = 1'b1;
  assign \A[6][47] [1] = 1'b1;
  assign \A[6][47] [0] = 1'b1;
  assign \A[6][48] [4] = 1'b1;
  assign \A[6][48] [3] = 1'b1;
  assign \A[6][48] [2] = 1'b1;
  assign \A[6][48] [1] = 1'b1;
  assign \A[6][48] [0] = 1'b1;
  assign \A[6][49] [1] = 1'b1;
  assign \A[6][49] [0] = 1'b1;
  assign \A[6][51] [1] = 1'b1;
  assign \A[6][52] [0] = 1'b1;
  assign \A[6][53] [0] = 1'b1;
  assign \A[6][56] [0] = 1'b1;
  assign \A[6][57] [4] = 1'b1;
  assign \A[6][57] [3] = 1'b1;
  assign \A[6][57] [2] = 1'b1;
  assign \A[6][57] [1] = 1'b1;
  assign \A[6][57] [0] = 1'b1;
  assign \A[6][58] [4] = 1'b1;
  assign \A[6][58] [3] = 1'b1;
  assign \A[6][58] [2] = 1'b1;
  assign \A[6][58] [1] = 1'b1;
  assign \A[6][58] [0] = 1'b1;
  assign \A[6][59] [4] = 1'b1;
  assign \A[6][59] [3] = 1'b1;
  assign \A[6][59] [2] = 1'b1;
  assign \A[6][59] [1] = 1'b1;
  assign \A[6][59] [0] = 1'b1;
  assign \A[6][60] [1] = 1'b1;
  assign \A[6][60] [0] = 1'b1;
  assign \A[6][61] [0] = 1'b1;
  assign \A[6][63] [1] = 1'b1;
  assign \A[6][64] [0] = 1'b1;
  assign \A[6][65] [1] = 1'b1;
  assign \A[6][65] [0] = 1'b1;
  assign \A[6][66] [1] = 1'b1;
  assign \A[6][66] [0] = 1'b1;
  assign \A[6][67] [0] = 1'b1;
  assign \A[6][69] [0] = 1'b1;
  assign \A[6][71] [1] = 1'b1;
  assign \A[6][71] [0] = 1'b1;
  assign \A[6][73] [4] = 1'b1;
  assign \A[6][73] [3] = 1'b1;
  assign \A[6][73] [2] = 1'b1;
  assign \A[6][73] [1] = 1'b1;
  assign \A[6][73] [0] = 1'b1;
  assign \A[6][75] [0] = 1'b1;
  assign \A[6][76] [0] = 1'b1;
  assign \A[6][77] [0] = 1'b1;
  assign \A[6][79] [2] = 1'b1;
  assign \A[6][81] [1] = 1'b1;
  assign \A[6][81] [0] = 1'b1;
  assign \A[6][82] [1] = 1'b1;
  assign \A[6][83] [0] = 1'b1;
  assign \A[6][84] [1] = 1'b1;
  assign \A[6][85] [1] = 1'b1;
  assign \A[6][85] [0] = 1'b1;
  assign \A[6][86] [1] = 1'b1;
  assign \A[6][86] [0] = 1'b1;
  assign \A[6][87] [4] = 1'b1;
  assign \A[6][87] [3] = 1'b1;
  assign \A[6][87] [2] = 1'b1;
  assign \A[6][87] [1] = 1'b1;
  assign \A[6][90] [4] = 1'b1;
  assign \A[6][90] [3] = 1'b1;
  assign \A[6][90] [2] = 1'b1;
  assign \A[6][90] [1] = 1'b1;
  assign \A[6][91] [4] = 1'b1;
  assign \A[6][91] [3] = 1'b1;
  assign \A[6][91] [2] = 1'b1;
  assign \A[6][91] [0] = 1'b1;
  assign \A[6][92] [0] = 1'b1;
  assign \A[6][93] [1] = 1'b1;
  assign \A[6][94] [4] = 1'b1;
  assign \A[6][94] [3] = 1'b1;
  assign \A[6][94] [2] = 1'b1;
  assign \A[6][94] [1] = 1'b1;
  assign \A[6][94] [0] = 1'b1;
  assign \A[6][96] [1] = 1'b1;
  assign \A[6][97] [0] = 1'b1;
  assign \A[6][98] [1] = 1'b1;
  assign \A[6][99] [4] = 1'b1;
  assign \A[6][99] [3] = 1'b1;
  assign \A[6][99] [2] = 1'b1;
  assign \A[6][99] [1] = 1'b1;
  assign \A[6][99] [0] = 1'b1;
  assign \A[6][100] [1] = 1'b1;
  assign \A[6][101] [0] = 1'b1;
  assign \A[6][102] [0] = 1'b1;
  assign \A[6][105] [1] = 1'b1;
  assign \A[6][105] [0] = 1'b1;
  assign \A[6][106] [0] = 1'b1;
  assign \A[6][107] [1] = 1'b1;
  assign \A[6][109] [1] = 1'b1;
  assign \A[6][110] [1] = 1'b1;
  assign \A[6][111] [0] = 1'b1;
  assign \A[6][112] [0] = 1'b1;
  assign \A[6][113] [1] = 1'b1;
  assign \A[6][114] [1] = 1'b1;
  assign \A[6][114] [0] = 1'b1;
  assign \A[6][115] [0] = 1'b1;
  assign \A[6][117] [1] = 1'b1;
  assign \A[6][118] [4] = 1'b1;
  assign \A[6][118] [3] = 1'b1;
  assign \A[6][118] [2] = 1'b1;
  assign \A[6][118] [1] = 1'b1;
  assign \A[6][118] [0] = 1'b1;
  assign \A[6][119] [0] = 1'b1;
  assign \A[6][120] [4] = 1'b1;
  assign \A[6][120] [3] = 1'b1;
  assign \A[6][120] [2] = 1'b1;
  assign \A[6][120] [1] = 1'b1;
  assign \A[6][120] [0] = 1'b1;
  assign \A[6][121] [1] = 1'b1;
  assign \A[6][121] [0] = 1'b1;
  assign \A[6][122] [4] = 1'b1;
  assign \A[6][122] [3] = 1'b1;
  assign \A[6][122] [2] = 1'b1;
  assign \A[6][122] [1] = 1'b1;
  assign \A[6][125] [4] = 1'b1;
  assign \A[6][125] [3] = 1'b1;
  assign \A[6][125] [2] = 1'b1;
  assign \A[6][125] [1] = 1'b1;
  assign \A[6][125] [0] = 1'b1;
  assign \A[6][126] [4] = 1'b1;
  assign \A[6][126] [3] = 1'b1;
  assign \A[6][126] [2] = 1'b1;
  assign \A[6][126] [1] = 1'b1;
  assign \A[6][126] [0] = 1'b1;
  assign \A[6][127] [1] = 1'b1;
  assign \A[6][128] [4] = 1'b1;
  assign \A[6][128] [3] = 1'b1;
  assign \A[6][128] [2] = 1'b1;
  assign \A[6][128] [1] = 1'b1;
  assign \A[6][128] [0] = 1'b1;
  assign \A[6][129] [1] = 1'b1;
  assign \A[6][131] [0] = 1'b1;
  assign \A[6][132] [1] = 1'b1;
  assign \A[6][133] [4] = 1'b1;
  assign \A[6][133] [3] = 1'b1;
  assign \A[6][133] [2] = 1'b1;
  assign \A[6][133] [1] = 1'b1;
  assign \A[6][133] [0] = 1'b1;
  assign \A[6][135] [4] = 1'b1;
  assign \A[6][135] [3] = 1'b1;
  assign \A[6][135] [2] = 1'b1;
  assign \A[6][135] [1] = 1'b1;
  assign \A[6][136] [0] = 1'b1;
  assign \A[6][138] [4] = 1'b1;
  assign \A[6][138] [3] = 1'b1;
  assign \A[6][138] [2] = 1'b1;
  assign \A[6][138] [1] = 1'b1;
  assign \A[6][139] [1] = 1'b1;
  assign \A[6][140] [4] = 1'b1;
  assign \A[6][140] [3] = 1'b1;
  assign \A[6][140] [2] = 1'b1;
  assign \A[6][140] [1] = 1'b1;
  assign \A[6][142] [0] = 1'b1;
  assign \A[6][143] [1] = 1'b1;
  assign \A[6][144] [1] = 1'b1;
  assign \A[6][144] [0] = 1'b1;
  assign \A[6][145] [4] = 1'b1;
  assign \A[6][145] [3] = 1'b1;
  assign \A[6][145] [2] = 1'b1;
  assign \A[6][145] [1] = 1'b1;
  assign \A[6][145] [0] = 1'b1;
  assign \A[6][146] [0] = 1'b1;
  assign \A[6][148] [4] = 1'b1;
  assign \A[6][148] [3] = 1'b1;
  assign \A[6][148] [2] = 1'b1;
  assign \A[6][148] [1] = 1'b1;
  assign \A[6][148] [0] = 1'b1;
  assign \A[6][150] [4] = 1'b1;
  assign \A[6][150] [3] = 1'b1;
  assign \A[6][150] [2] = 1'b1;
  assign \A[6][150] [1] = 1'b1;
  assign \A[6][150] [0] = 1'b1;
  assign \A[6][151] [4] = 1'b1;
  assign \A[6][151] [3] = 1'b1;
  assign \A[6][151] [2] = 1'b1;
  assign \A[6][151] [1] = 1'b1;
  assign \A[6][151] [0] = 1'b1;
  assign \A[6][153] [4] = 1'b1;
  assign \A[6][153] [3] = 1'b1;
  assign \A[6][153] [2] = 1'b1;
  assign \A[6][153] [1] = 1'b1;
  assign \A[6][154] [0] = 1'b1;
  assign \A[6][155] [1] = 1'b1;
  assign \A[6][156] [0] = 1'b1;
  assign \A[6][157] [4] = 1'b1;
  assign \A[6][157] [3] = 1'b1;
  assign \A[6][157] [2] = 1'b1;
  assign \A[6][157] [1] = 1'b1;
  assign \A[6][158] [4] = 1'b1;
  assign \A[6][158] [3] = 1'b1;
  assign \A[6][158] [2] = 1'b1;
  assign \A[6][158] [1] = 1'b1;
  assign \A[6][158] [0] = 1'b1;
  assign \A[6][159] [0] = 1'b1;
  assign \A[6][160] [0] = 1'b1;
  assign \A[6][161] [4] = 1'b1;
  assign \A[6][161] [3] = 1'b1;
  assign \A[6][161] [2] = 1'b1;
  assign \A[6][161] [1] = 1'b1;
  assign \A[6][161] [0] = 1'b1;
  assign \A[6][163] [4] = 1'b1;
  assign \A[6][163] [3] = 1'b1;
  assign \A[6][163] [2] = 1'b1;
  assign \A[6][163] [1] = 1'b1;
  assign \A[6][163] [0] = 1'b1;
  assign \A[6][164] [4] = 1'b1;
  assign \A[6][164] [3] = 1'b1;
  assign \A[6][164] [2] = 1'b1;
  assign \A[6][164] [1] = 1'b1;
  assign \A[6][165] [0] = 1'b1;
  assign \A[6][167] [0] = 1'b1;
  assign \A[6][168] [0] = 1'b1;
  assign \A[6][170] [4] = 1'b1;
  assign \A[6][170] [3] = 1'b1;
  assign \A[6][170] [2] = 1'b1;
  assign \A[6][170] [0] = 1'b1;
  assign \A[6][171] [1] = 1'b1;
  assign \A[6][171] [0] = 1'b1;
  assign \A[6][172] [1] = 1'b1;
  assign \A[6][172] [0] = 1'b1;
  assign \A[6][173] [1] = 1'b1;
  assign \A[6][175] [4] = 1'b1;
  assign \A[6][175] [3] = 1'b1;
  assign \A[6][175] [2] = 1'b1;
  assign \A[6][175] [1] = 1'b1;
  assign \A[6][175] [0] = 1'b1;
  assign \A[6][177] [4] = 1'b1;
  assign \A[6][177] [3] = 1'b1;
  assign \A[6][177] [2] = 1'b1;
  assign \A[6][177] [1] = 1'b1;
  assign \A[6][177] [0] = 1'b1;
  assign \A[6][178] [4] = 1'b1;
  assign \A[6][178] [3] = 1'b1;
  assign \A[6][178] [2] = 1'b1;
  assign \A[6][178] [1] = 1'b1;
  assign \A[6][178] [0] = 1'b1;
  assign \A[6][179] [4] = 1'b1;
  assign \A[6][179] [3] = 1'b1;
  assign \A[6][179] [2] = 1'b1;
  assign \A[6][180] [4] = 1'b1;
  assign \A[6][180] [3] = 1'b1;
  assign \A[6][180] [2] = 1'b1;
  assign \A[6][182] [4] = 1'b1;
  assign \A[6][182] [3] = 1'b1;
  assign \A[6][182] [2] = 1'b1;
  assign \A[6][182] [1] = 1'b1;
  assign \A[6][183] [4] = 1'b1;
  assign \A[6][183] [3] = 1'b1;
  assign \A[6][183] [2] = 1'b1;
  assign \A[6][184] [0] = 1'b1;
  assign \A[6][185] [1] = 1'b1;
  assign \A[6][187] [4] = 1'b1;
  assign \A[6][187] [3] = 1'b1;
  assign \A[6][187] [2] = 1'b1;
  assign \A[6][187] [1] = 1'b1;
  assign \A[6][188] [4] = 1'b1;
  assign \A[6][188] [3] = 1'b1;
  assign \A[6][188] [2] = 1'b1;
  assign \A[6][188] [1] = 1'b1;
  assign \A[6][189] [0] = 1'b1;
  assign \A[6][190] [4] = 1'b1;
  assign \A[6][190] [3] = 1'b1;
  assign \A[6][190] [2] = 1'b1;
  assign \A[6][190] [1] = 1'b1;
  assign \A[6][190] [0] = 1'b1;
  assign \A[6][191] [0] = 1'b1;
  assign \A[6][193] [4] = 1'b1;
  assign \A[6][193] [3] = 1'b1;
  assign \A[6][193] [2] = 1'b1;
  assign \A[6][193] [1] = 1'b1;
  assign \A[6][193] [0] = 1'b1;
  assign \A[6][194] [4] = 1'b1;
  assign \A[6][194] [3] = 1'b1;
  assign \A[6][194] [2] = 1'b1;
  assign \A[6][194] [0] = 1'b1;
  assign \A[6][195] [0] = 1'b1;
  assign \A[6][196] [4] = 1'b1;
  assign \A[6][196] [3] = 1'b1;
  assign \A[6][196] [2] = 1'b1;
  assign \A[6][196] [1] = 1'b1;
  assign \A[6][197] [4] = 1'b1;
  assign \A[6][197] [3] = 1'b1;
  assign \A[6][197] [2] = 1'b1;
  assign \A[6][197] [1] = 1'b1;
  assign \A[6][198] [4] = 1'b1;
  assign \A[6][198] [3] = 1'b1;
  assign \A[6][198] [2] = 1'b1;
  assign \A[6][198] [1] = 1'b1;
  assign \A[6][200] [0] = 1'b1;
  assign \A[6][201] [4] = 1'b1;
  assign \A[6][201] [3] = 1'b1;
  assign \A[6][201] [2] = 1'b1;
  assign \A[6][201] [1] = 1'b1;
  assign \A[6][201] [0] = 1'b1;
  assign \A[6][203] [4] = 1'b1;
  assign \A[6][203] [3] = 1'b1;
  assign \A[6][203] [2] = 1'b1;
  assign \A[6][203] [1] = 1'b1;
  assign \A[6][203] [0] = 1'b1;
  assign \A[6][204] [4] = 1'b1;
  assign \A[6][204] [3] = 1'b1;
  assign \A[6][204] [2] = 1'b1;
  assign \A[6][204] [1] = 1'b1;
  assign \A[6][204] [0] = 1'b1;
  assign \A[6][205] [4] = 1'b1;
  assign \A[6][205] [3] = 1'b1;
  assign \A[6][205] [2] = 1'b1;
  assign \A[6][205] [1] = 1'b1;
  assign \A[6][206] [0] = 1'b1;
  assign \A[6][207] [1] = 1'b1;
  assign \A[6][208] [0] = 1'b1;
  assign \A[6][209] [0] = 1'b1;
  assign \A[6][210] [4] = 1'b1;
  assign \A[6][210] [3] = 1'b1;
  assign \A[6][210] [2] = 1'b1;
  assign \A[6][210] [1] = 1'b1;
  assign \A[6][210] [0] = 1'b1;
  assign \A[6][211] [1] = 1'b1;
  assign \A[6][213] [1] = 1'b1;
  assign \A[6][215] [4] = 1'b1;
  assign \A[6][215] [3] = 1'b1;
  assign \A[6][215] [2] = 1'b1;
  assign \A[6][215] [1] = 1'b1;
  assign \A[6][217] [4] = 1'b1;
  assign \A[6][217] [3] = 1'b1;
  assign \A[6][217] [2] = 1'b1;
  assign \A[6][217] [1] = 1'b1;
  assign \A[6][217] [0] = 1'b1;
  assign \A[6][218] [4] = 1'b1;
  assign \A[6][218] [3] = 1'b1;
  assign \A[6][218] [2] = 1'b1;
  assign \A[6][218] [1] = 1'b1;
  assign \A[6][218] [0] = 1'b1;
  assign \A[6][220] [0] = 1'b1;
  assign \A[6][221] [4] = 1'b1;
  assign \A[6][221] [3] = 1'b1;
  assign \A[6][221] [2] = 1'b1;
  assign \A[6][221] [1] = 1'b1;
  assign \A[6][222] [4] = 1'b1;
  assign \A[6][222] [3] = 1'b1;
  assign \A[6][222] [2] = 1'b1;
  assign \A[6][222] [0] = 1'b1;
  assign \A[6][223] [4] = 1'b1;
  assign \A[6][223] [3] = 1'b1;
  assign \A[6][223] [2] = 1'b1;
  assign \A[6][223] [1] = 1'b1;
  assign \A[6][223] [0] = 1'b1;
  assign \A[6][225] [0] = 1'b1;
  assign \A[6][226] [4] = 1'b1;
  assign \A[6][226] [3] = 1'b1;
  assign \A[6][226] [2] = 1'b1;
  assign \A[6][226] [1] = 1'b1;
  assign \A[6][226] [0] = 1'b1;
  assign \A[6][227] [4] = 1'b1;
  assign \A[6][227] [3] = 1'b1;
  assign \A[6][227] [2] = 1'b1;
  assign \A[6][227] [1] = 1'b1;
  assign \A[6][227] [0] = 1'b1;
  assign \A[6][228] [4] = 1'b1;
  assign \A[6][228] [3] = 1'b1;
  assign \A[6][228] [2] = 1'b1;
  assign \A[6][228] [1] = 1'b1;
  assign \A[6][228] [0] = 1'b1;
  assign \A[6][229] [4] = 1'b1;
  assign \A[6][229] [3] = 1'b1;
  assign \A[6][229] [2] = 1'b1;
  assign \A[6][229] [0] = 1'b1;
  assign \A[6][230] [0] = 1'b1;
  assign \A[6][231] [4] = 1'b1;
  assign \A[6][231] [3] = 1'b1;
  assign \A[6][231] [2] = 1'b1;
  assign \A[6][231] [0] = 1'b1;
  assign \A[6][233] [4] = 1'b1;
  assign \A[6][233] [3] = 1'b1;
  assign \A[6][233] [2] = 1'b1;
  assign \A[6][233] [1] = 1'b1;
  assign \A[6][233] [0] = 1'b1;
  assign \A[6][234] [4] = 1'b1;
  assign \A[6][234] [3] = 1'b1;
  assign \A[6][234] [2] = 1'b1;
  assign \A[6][234] [0] = 1'b1;
  assign \A[6][237] [4] = 1'b1;
  assign \A[6][237] [3] = 1'b1;
  assign \A[6][237] [2] = 1'b1;
  assign \A[6][237] [1] = 1'b1;
  assign \A[6][238] [4] = 1'b1;
  assign \A[6][238] [3] = 1'b1;
  assign \A[6][238] [2] = 1'b1;
  assign \A[6][238] [0] = 1'b1;
  assign \A[6][239] [4] = 1'b1;
  assign \A[6][239] [3] = 1'b1;
  assign \A[6][239] [2] = 1'b1;
  assign \A[6][239] [1] = 1'b1;
  assign \A[6][240] [0] = 1'b1;
  assign \A[6][241] [0] = 1'b1;
  assign \A[6][242] [0] = 1'b1;
  assign \A[6][243] [0] = 1'b1;
  assign \A[6][244] [4] = 1'b1;
  assign \A[6][244] [3] = 1'b1;
  assign \A[6][244] [2] = 1'b1;
  assign \A[6][244] [1] = 1'b1;
  assign \A[6][244] [0] = 1'b1;
  assign \A[6][246] [1] = 1'b1;
  assign \A[6][246] [0] = 1'b1;
  assign \A[6][247] [4] = 1'b1;
  assign \A[6][247] [3] = 1'b1;
  assign \A[6][247] [2] = 1'b1;
  assign \A[6][247] [1] = 1'b1;
  assign \A[6][247] [0] = 1'b1;
  assign \A[6][250] [0] = 1'b1;
  assign \A[6][251] [1] = 1'b1;
  assign \A[6][252] [4] = 1'b1;
  assign \A[6][252] [3] = 1'b1;
  assign \A[6][252] [2] = 1'b1;
  assign \A[6][252] [1] = 1'b1;
  assign \A[6][253] [1] = 1'b1;
  assign \A[6][254] [4] = 1'b1;
  assign \A[6][254] [3] = 1'b1;
  assign \A[6][254] [2] = 1'b1;
  assign \A[6][254] [1] = 1'b1;
  assign \A[6][254] [0] = 1'b1;
  assign \A[6][255] [4] = 1'b1;
  assign \A[6][255] [3] = 1'b1;
  assign \A[6][255] [2] = 1'b1;
  assign \A[6][255] [0] = 1'b1;
  assign \A[7][0] [4] = 1'b1;
  assign \A[7][0] [3] = 1'b1;
  assign \A[7][0] [2] = 1'b1;
  assign \A[7][0] [1] = 1'b1;
  assign \A[7][0] [0] = 1'b1;
  assign \A[7][1] [4] = 1'b1;
  assign \A[7][1] [3] = 1'b1;
  assign \A[7][1] [2] = 1'b1;
  assign \A[7][1] [1] = 1'b1;
  assign \A[7][1] [0] = 1'b1;
  assign \A[7][4] [4] = 1'b1;
  assign \A[7][4] [3] = 1'b1;
  assign \A[7][4] [2] = 1'b1;
  assign \A[7][4] [1] = 1'b1;
  assign \A[7][6] [1] = 1'b1;
  assign \A[7][7] [0] = 1'b1;
  assign \A[7][8] [4] = 1'b1;
  assign \A[7][8] [3] = 1'b1;
  assign \A[7][8] [2] = 1'b1;
  assign \A[7][8] [1] = 1'b1;
  assign \A[7][9] [4] = 1'b1;
  assign \A[7][9] [3] = 1'b1;
  assign \A[7][9] [2] = 1'b1;
  assign \A[7][9] [1] = 1'b1;
  assign \A[7][9] [0] = 1'b1;
  assign \A[7][10] [0] = 1'b1;
  assign \A[7][11] [4] = 1'b1;
  assign \A[7][11] [3] = 1'b1;
  assign \A[7][11] [2] = 1'b1;
  assign \A[7][11] [1] = 1'b1;
  assign \A[7][11] [0] = 1'b1;
  assign \A[7][12] [1] = 1'b1;
  assign \A[7][13] [4] = 1'b1;
  assign \A[7][13] [3] = 1'b1;
  assign \A[7][13] [2] = 1'b1;
  assign \A[7][13] [1] = 1'b1;
  assign \A[7][13] [0] = 1'b1;
  assign \A[7][14] [4] = 1'b1;
  assign \A[7][14] [3] = 1'b1;
  assign \A[7][14] [2] = 1'b1;
  assign \A[7][14] [1] = 1'b1;
  assign \A[7][14] [0] = 1'b1;
  assign \A[7][15] [1] = 1'b1;
  assign \A[7][16] [0] = 1'b1;
  assign \A[7][17] [0] = 1'b1;
  assign \A[7][18] [4] = 1'b1;
  assign \A[7][18] [3] = 1'b1;
  assign \A[7][18] [2] = 1'b1;
  assign \A[7][18] [1] = 1'b1;
  assign \A[7][21] [4] = 1'b1;
  assign \A[7][21] [3] = 1'b1;
  assign \A[7][21] [2] = 1'b1;
  assign \A[7][21] [1] = 1'b1;
  assign \A[7][22] [4] = 1'b1;
  assign \A[7][22] [3] = 1'b1;
  assign \A[7][22] [2] = 1'b1;
  assign \A[7][22] [1] = 1'b1;
  assign \A[7][22] [0] = 1'b1;
  assign \A[7][23] [0] = 1'b1;
  assign \A[7][24] [0] = 1'b1;
  assign \A[7][25] [2] = 1'b1;
  assign \A[7][26] [4] = 1'b1;
  assign \A[7][26] [3] = 1'b1;
  assign \A[7][26] [2] = 1'b1;
  assign \A[7][26] [0] = 1'b1;
  assign \A[7][28] [0] = 1'b1;
  assign \A[7][29] [4] = 1'b1;
  assign \A[7][29] [3] = 1'b1;
  assign \A[7][29] [2] = 1'b1;
  assign \A[7][29] [0] = 1'b1;
  assign \A[7][31] [1] = 1'b1;
  assign \A[7][35] [0] = 1'b1;
  assign \A[7][38] [4] = 1'b1;
  assign \A[7][38] [3] = 1'b1;
  assign \A[7][38] [2] = 1'b1;
  assign \A[7][38] [1] = 1'b1;
  assign \A[7][39] [4] = 1'b1;
  assign \A[7][39] [3] = 1'b1;
  assign \A[7][39] [2] = 1'b1;
  assign \A[7][39] [0] = 1'b1;
  assign \A[7][40] [4] = 1'b1;
  assign \A[7][40] [3] = 1'b1;
  assign \A[7][40] [2] = 1'b1;
  assign \A[7][40] [1] = 1'b1;
  assign \A[7][40] [0] = 1'b1;
  assign \A[7][41] [4] = 1'b1;
  assign \A[7][41] [3] = 1'b1;
  assign \A[7][41] [2] = 1'b1;
  assign \A[7][41] [1] = 1'b1;
  assign \A[7][42] [4] = 1'b1;
  assign \A[7][42] [3] = 1'b1;
  assign \A[7][42] [2] = 1'b1;
  assign \A[7][42] [1] = 1'b1;
  assign \A[7][43] [4] = 1'b1;
  assign \A[7][43] [3] = 1'b1;
  assign \A[7][43] [2] = 1'b1;
  assign \A[7][43] [1] = 1'b1;
  assign \A[7][43] [0] = 1'b1;
  assign \A[7][44] [0] = 1'b1;
  assign \A[7][45] [0] = 1'b1;
  assign \A[7][46] [4] = 1'b1;
  assign \A[7][46] [3] = 1'b1;
  assign \A[7][46] [2] = 1'b1;
  assign \A[7][46] [1] = 1'b1;
  assign \A[7][46] [0] = 1'b1;
  assign \A[7][47] [0] = 1'b1;
  assign \A[7][48] [0] = 1'b1;
  assign \A[7][49] [4] = 1'b1;
  assign \A[7][49] [3] = 1'b1;
  assign \A[7][49] [2] = 1'b1;
  assign \A[7][49] [1] = 1'b1;
  assign \A[7][50] [1] = 1'b1;
  assign \A[7][51] [4] = 1'b1;
  assign \A[7][51] [3] = 1'b1;
  assign \A[7][51] [2] = 1'b1;
  assign \A[7][51] [0] = 1'b1;
  assign \A[7][52] [0] = 1'b1;
  assign \A[7][55] [0] = 1'b1;
  assign \A[7][56] [4] = 1'b1;
  assign \A[7][56] [3] = 1'b1;
  assign \A[7][56] [2] = 1'b1;
  assign \A[7][56] [1] = 1'b1;
  assign \A[7][56] [0] = 1'b1;
  assign \A[7][57] [4] = 1'b1;
  assign \A[7][57] [3] = 1'b1;
  assign \A[7][57] [2] = 1'b1;
  assign \A[7][58] [4] = 1'b1;
  assign \A[7][58] [3] = 1'b1;
  assign \A[7][58] [1] = 1'b1;
  assign \A[7][58] [0] = 1'b1;
  assign \A[7][59] [4] = 1'b1;
  assign \A[7][59] [3] = 1'b1;
  assign \A[7][59] [2] = 1'b1;
  assign \A[7][59] [1] = 1'b1;
  assign \A[7][62] [4] = 1'b1;
  assign \A[7][62] [3] = 1'b1;
  assign \A[7][62] [2] = 1'b1;
  assign \A[7][62] [0] = 1'b1;
  assign \A[7][63] [4] = 1'b1;
  assign \A[7][63] [3] = 1'b1;
  assign \A[7][63] [2] = 1'b1;
  assign \A[7][63] [1] = 1'b1;
  assign \A[7][64] [4] = 1'b1;
  assign \A[7][64] [3] = 1'b1;
  assign \A[7][64] [2] = 1'b1;
  assign \A[7][64] [1] = 1'b1;
  assign \A[7][65] [1] = 1'b1;
  assign \A[7][66] [0] = 1'b1;
  assign \A[7][67] [4] = 1'b1;
  assign \A[7][67] [3] = 1'b1;
  assign \A[7][67] [2] = 1'b1;
  assign \A[7][67] [1] = 1'b1;
  assign \A[7][67] [0] = 1'b1;
  assign \A[7][68] [0] = 1'b1;
  assign \A[7][69] [4] = 1'b1;
  assign \A[7][69] [3] = 1'b1;
  assign \A[7][69] [2] = 1'b1;
  assign \A[7][69] [1] = 1'b1;
  assign \A[7][69] [0] = 1'b1;
  assign \A[7][70] [4] = 1'b1;
  assign \A[7][70] [3] = 1'b1;
  assign \A[7][70] [2] = 1'b1;
  assign \A[7][70] [1] = 1'b1;
  assign \A[7][71] [0] = 1'b1;
  assign \A[7][72] [0] = 1'b1;
  assign \A[7][73] [4] = 1'b1;
  assign \A[7][73] [3] = 1'b1;
  assign \A[7][73] [2] = 1'b1;
  assign \A[7][73] [0] = 1'b1;
  assign \A[7][74] [4] = 1'b1;
  assign \A[7][74] [3] = 1'b1;
  assign \A[7][74] [1] = 1'b1;
  assign \A[7][74] [0] = 1'b1;
  assign \A[7][75] [4] = 1'b1;
  assign \A[7][75] [3] = 1'b1;
  assign \A[7][75] [2] = 1'b1;
  assign \A[7][75] [0] = 1'b1;
  assign \A[7][76] [4] = 1'b1;
  assign \A[7][76] [3] = 1'b1;
  assign \A[7][76] [2] = 1'b1;
  assign \A[7][76] [1] = 1'b1;
  assign \A[7][77] [4] = 1'b1;
  assign \A[7][77] [3] = 1'b1;
  assign \A[7][77] [2] = 1'b1;
  assign \A[7][77] [0] = 1'b1;
  assign \A[7][78] [4] = 1'b1;
  assign \A[7][78] [3] = 1'b1;
  assign \A[7][78] [2] = 1'b1;
  assign \A[7][78] [1] = 1'b1;
  assign \A[7][80] [4] = 1'b1;
  assign \A[7][80] [3] = 1'b1;
  assign \A[7][80] [2] = 1'b1;
  assign \A[7][80] [1] = 1'b1;
  assign \A[7][80] [0] = 1'b1;
  assign \A[7][81] [4] = 1'b1;
  assign \A[7][81] [3] = 1'b1;
  assign \A[7][81] [2] = 1'b1;
  assign \A[7][81] [1] = 1'b1;
  assign \A[7][82] [4] = 1'b1;
  assign \A[7][82] [3] = 1'b1;
  assign \A[7][82] [2] = 1'b1;
  assign \A[7][82] [1] = 1'b1;
  assign \A[7][82] [0] = 1'b1;
  assign \A[7][83] [4] = 1'b1;
  assign \A[7][83] [3] = 1'b1;
  assign \A[7][83] [2] = 1'b1;
  assign \A[7][83] [1] = 1'b1;
  assign \A[7][84] [4] = 1'b1;
  assign \A[7][84] [3] = 1'b1;
  assign \A[7][84] [2] = 1'b1;
  assign \A[7][84] [1] = 1'b1;
  assign \A[7][85] [0] = 1'b1;
  assign \A[7][86] [2] = 1'b1;
  assign \A[7][86] [0] = 1'b1;
  assign \A[7][87] [0] = 1'b1;
  assign \A[7][88] [0] = 1'b1;
  assign \A[7][92] [4] = 1'b1;
  assign \A[7][92] [3] = 1'b1;
  assign \A[7][92] [2] = 1'b1;
  assign \A[7][92] [1] = 1'b1;
  assign \A[7][92] [0] = 1'b1;
  assign \A[7][93] [4] = 1'b1;
  assign \A[7][93] [3] = 1'b1;
  assign \A[7][93] [2] = 1'b1;
  assign \A[7][93] [1] = 1'b1;
  assign \A[7][94] [4] = 1'b1;
  assign \A[7][94] [3] = 1'b1;
  assign \A[7][94] [2] = 1'b1;
  assign \A[7][95] [4] = 1'b1;
  assign \A[7][95] [3] = 1'b1;
  assign \A[7][95] [2] = 1'b1;
  assign \A[7][95] [0] = 1'b1;
  assign \A[7][97] [4] = 1'b1;
  assign \A[7][97] [3] = 1'b1;
  assign \A[7][97] [2] = 1'b1;
  assign \A[7][97] [1] = 1'b1;
  assign \A[7][97] [0] = 1'b1;
  assign \A[7][98] [4] = 1'b1;
  assign \A[7][98] [3] = 1'b1;
  assign \A[7][98] [2] = 1'b1;
  assign \A[7][98] [1] = 1'b1;
  assign \A[7][99] [4] = 1'b1;
  assign \A[7][99] [3] = 1'b1;
  assign \A[7][99] [2] = 1'b1;
  assign \A[7][99] [1] = 1'b1;
  assign \A[7][99] [0] = 1'b1;
  assign \A[7][100] [0] = 1'b1;
  assign \A[7][101] [0] = 1'b1;
  assign \A[7][102] [2] = 1'b1;
  assign \A[7][102] [0] = 1'b1;
  assign \A[7][103] [4] = 1'b1;
  assign \A[7][103] [3] = 1'b1;
  assign \A[7][103] [2] = 1'b1;
  assign \A[7][103] [1] = 1'b1;
  assign \A[7][103] [0] = 1'b1;
  assign \A[7][104] [0] = 1'b1;
  assign \A[7][107] [1] = 1'b1;
  assign \A[7][109] [4] = 1'b1;
  assign \A[7][109] [3] = 1'b1;
  assign \A[7][109] [2] = 1'b1;
  assign \A[7][109] [1] = 1'b1;
  assign \A[7][111] [4] = 1'b1;
  assign \A[7][111] [3] = 1'b1;
  assign \A[7][111] [1] = 1'b1;
  assign \A[7][111] [0] = 1'b1;
  assign \A[7][113] [4] = 1'b1;
  assign \A[7][113] [3] = 1'b1;
  assign \A[7][113] [2] = 1'b1;
  assign \A[7][113] [1] = 1'b1;
  assign \A[7][113] [0] = 1'b1;
  assign \A[7][114] [0] = 1'b1;
  assign \A[7][117] [0] = 1'b1;
  assign \A[7][118] [0] = 1'b1;
  assign \A[7][120] [0] = 1'b1;
  assign \A[7][121] [4] = 1'b1;
  assign \A[7][121] [3] = 1'b1;
  assign \A[7][121] [2] = 1'b1;
  assign \A[7][121] [1] = 1'b1;
  assign \A[7][121] [0] = 1'b1;
  assign \A[7][124] [2] = 1'b1;
  assign \A[7][126] [4] = 1'b1;
  assign \A[7][126] [3] = 1'b1;
  assign \A[7][126] [2] = 1'b1;
  assign \A[7][126] [1] = 1'b1;
  assign \A[7][127] [4] = 1'b1;
  assign \A[7][127] [3] = 1'b1;
  assign \A[7][127] [2] = 1'b1;
  assign \A[7][127] [1] = 1'b1;
  assign \A[7][127] [0] = 1'b1;
  assign \A[7][128] [1] = 1'b1;
  assign \A[7][129] [4] = 1'b1;
  assign \A[7][129] [3] = 1'b1;
  assign \A[7][129] [2] = 1'b1;
  assign \A[7][129] [1] = 1'b1;
  assign \A[7][130] [1] = 1'b1;
  assign \A[7][130] [0] = 1'b1;
  assign \A[7][133] [0] = 1'b1;
  assign \A[7][134] [0] = 1'b1;
  assign \A[7][135] [1] = 1'b1;
  assign \A[7][135] [0] = 1'b1;
  assign \A[7][136] [0] = 1'b1;
  assign \A[7][138] [1] = 1'b1;
  assign \A[7][142] [4] = 1'b1;
  assign \A[7][142] [3] = 1'b1;
  assign \A[7][142] [2] = 1'b1;
  assign \A[7][142] [1] = 1'b1;
  assign \A[7][142] [0] = 1'b1;
  assign \A[7][143] [4] = 1'b1;
  assign \A[7][143] [3] = 1'b1;
  assign \A[7][143] [2] = 1'b1;
  assign \A[7][143] [1] = 1'b1;
  assign \A[7][143] [0] = 1'b1;
  assign \A[7][144] [0] = 1'b1;
  assign \A[7][145] [1] = 1'b1;
  assign \A[7][146] [4] = 1'b1;
  assign \A[7][146] [3] = 1'b1;
  assign \A[7][146] [2] = 1'b1;
  assign \A[7][146] [0] = 1'b1;
  assign \A[7][149] [0] = 1'b1;
  assign \A[7][150] [0] = 1'b1;
  assign \A[7][151] [0] = 1'b1;
  assign \A[7][152] [0] = 1'b1;
  assign \A[7][153] [0] = 1'b1;
  assign \A[7][154] [1] = 1'b1;
  assign \A[7][156] [0] = 1'b1;
  assign \A[7][157] [0] = 1'b1;
  assign \A[7][158] [4] = 1'b1;
  assign \A[7][158] [3] = 1'b1;
  assign \A[7][158] [2] = 1'b1;
  assign \A[7][158] [1] = 1'b1;
  assign \A[7][158] [0] = 1'b1;
  assign \A[7][159] [0] = 1'b1;
  assign \A[7][161] [0] = 1'b1;
  assign \A[7][162] [0] = 1'b1;
  assign \A[7][163] [1] = 1'b1;
  assign \A[7][165] [1] = 1'b1;
  assign \A[7][166] [1] = 1'b1;
  assign \A[7][167] [4] = 1'b1;
  assign \A[7][167] [3] = 1'b1;
  assign \A[7][167] [2] = 1'b1;
  assign \A[7][167] [1] = 1'b1;
  assign \A[7][167] [0] = 1'b1;
  assign \A[7][168] [1] = 1'b1;
  assign \A[7][169] [1] = 1'b1;
  assign \A[7][170] [4] = 1'b1;
  assign \A[7][170] [3] = 1'b1;
  assign \A[7][170] [2] = 1'b1;
  assign \A[7][170] [1] = 1'b1;
  assign \A[7][170] [0] = 1'b1;
  assign \A[7][171] [0] = 1'b1;
  assign \A[7][173] [1] = 1'b1;
  assign \A[7][173] [0] = 1'b1;
  assign \A[7][174] [0] = 1'b1;
  assign \A[7][176] [0] = 1'b1;
  assign \A[7][177] [2] = 1'b1;
  assign \A[7][177] [0] = 1'b1;
  assign \A[7][178] [0] = 1'b1;
  assign \A[7][179] [0] = 1'b1;
  assign \A[7][180] [4] = 1'b1;
  assign \A[7][180] [3] = 1'b1;
  assign \A[7][180] [2] = 1'b1;
  assign \A[7][180] [1] = 1'b1;
  assign \A[7][180] [0] = 1'b1;
  assign \A[7][181] [4] = 1'b1;
  assign \A[7][181] [3] = 1'b1;
  assign \A[7][181] [2] = 1'b1;
  assign \A[7][181] [1] = 1'b1;
  assign \A[7][181] [0] = 1'b1;
  assign \A[7][183] [0] = 1'b1;
  assign \A[7][184] [0] = 1'b1;
  assign \A[7][185] [0] = 1'b1;
  assign \A[7][186] [0] = 1'b1;
  assign \A[7][188] [1] = 1'b1;
  assign \A[7][190] [1] = 1'b1;
  assign \A[7][190] [0] = 1'b1;
  assign \A[7][191] [0] = 1'b1;
  assign \A[7][192] [1] = 1'b1;
  assign \A[7][192] [0] = 1'b1;
  assign \A[7][193] [2] = 1'b1;
  assign \A[7][193] [0] = 1'b1;
  assign \A[7][194] [0] = 1'b1;
  assign \A[7][196] [1] = 1'b1;
  assign \A[7][196] [0] = 1'b1;
  assign \A[7][197] [4] = 1'b1;
  assign \A[7][197] [3] = 1'b1;
  assign \A[7][197] [2] = 1'b1;
  assign \A[7][197] [1] = 1'b1;
  assign \A[7][197] [0] = 1'b1;
  assign \A[7][198] [4] = 1'b1;
  assign \A[7][198] [3] = 1'b1;
  assign \A[7][198] [2] = 1'b1;
  assign \A[7][198] [1] = 1'b1;
  assign \A[7][199] [0] = 1'b1;
  assign \A[7][201] [4] = 1'b1;
  assign \A[7][201] [3] = 1'b1;
  assign \A[7][201] [2] = 1'b1;
  assign \A[7][201] [0] = 1'b1;
  assign \A[7][202] [0] = 1'b1;
  assign \A[7][203] [1] = 1'b1;
  assign \A[7][205] [0] = 1'b1;
  assign \A[7][206] [0] = 1'b1;
  assign \A[7][207] [2] = 1'b1;
  assign \A[7][208] [0] = 1'b1;
  assign \A[7][210] [4] = 1'b1;
  assign \A[7][210] [3] = 1'b1;
  assign \A[7][210] [2] = 1'b1;
  assign \A[7][210] [1] = 1'b1;
  assign \A[7][210] [0] = 1'b1;
  assign \A[7][211] [4] = 1'b1;
  assign \A[7][211] [3] = 1'b1;
  assign \A[7][211] [2] = 1'b1;
  assign \A[7][211] [1] = 1'b1;
  assign \A[7][211] [0] = 1'b1;
  assign \A[7][212] [4] = 1'b1;
  assign \A[7][212] [3] = 1'b1;
  assign \A[7][212] [2] = 1'b1;
  assign \A[7][212] [1] = 1'b1;
  assign \A[7][212] [0] = 1'b1;
  assign \A[7][214] [4] = 1'b1;
  assign \A[7][214] [3] = 1'b1;
  assign \A[7][214] [2] = 1'b1;
  assign \A[7][214] [1] = 1'b1;
  assign \A[7][214] [0] = 1'b1;
  assign \A[7][215] [4] = 1'b1;
  assign \A[7][215] [3] = 1'b1;
  assign \A[7][215] [2] = 1'b1;
  assign \A[7][215] [1] = 1'b1;
  assign \A[7][216] [0] = 1'b1;
  assign \A[7][218] [4] = 1'b1;
  assign \A[7][218] [3] = 1'b1;
  assign \A[7][218] [2] = 1'b1;
  assign \A[7][218] [0] = 1'b1;
  assign \A[7][219] [4] = 1'b1;
  assign \A[7][219] [3] = 1'b1;
  assign \A[7][219] [2] = 1'b1;
  assign \A[7][219] [1] = 1'b1;
  assign \A[7][219] [0] = 1'b1;
  assign \A[7][220] [0] = 1'b1;
  assign \A[7][221] [4] = 1'b1;
  assign \A[7][221] [3] = 1'b1;
  assign \A[7][221] [1] = 1'b1;
  assign \A[7][221] [0] = 1'b1;
  assign \A[7][222] [0] = 1'b1;
  assign \A[7][224] [4] = 1'b1;
  assign \A[7][224] [3] = 1'b1;
  assign \A[7][224] [2] = 1'b1;
  assign \A[7][224] [1] = 1'b1;
  assign \A[7][225] [4] = 1'b1;
  assign \A[7][225] [3] = 1'b1;
  assign \A[7][225] [2] = 1'b1;
  assign \A[7][225] [1] = 1'b1;
  assign \A[7][225] [0] = 1'b1;
  assign \A[7][226] [4] = 1'b1;
  assign \A[7][226] [3] = 1'b1;
  assign \A[7][226] [2] = 1'b1;
  assign \A[7][226] [1] = 1'b1;
  assign \A[7][227] [1] = 1'b1;
  assign \A[7][228] [1] = 1'b1;
  assign \A[7][228] [0] = 1'b1;
  assign \A[7][229] [0] = 1'b1;
  assign \A[7][231] [2] = 1'b1;
  assign \A[7][233] [4] = 1'b1;
  assign \A[7][233] [3] = 1'b1;
  assign \A[7][233] [2] = 1'b1;
  assign \A[7][233] [1] = 1'b1;
  assign \A[7][233] [0] = 1'b1;
  assign \A[7][234] [1] = 1'b1;
  assign \A[7][238] [4] = 1'b1;
  assign \A[7][238] [3] = 1'b1;
  assign \A[7][238] [2] = 1'b1;
  assign \A[7][238] [0] = 1'b1;
  assign \A[7][239] [4] = 1'b1;
  assign \A[7][239] [3] = 1'b1;
  assign \A[7][239] [2] = 1'b1;
  assign \A[7][239] [0] = 1'b1;
  assign \A[7][240] [4] = 1'b1;
  assign \A[7][240] [3] = 1'b1;
  assign \A[7][240] [2] = 1'b1;
  assign \A[7][240] [1] = 1'b1;
  assign \A[7][241] [1] = 1'b1;
  assign \A[7][243] [1] = 1'b1;
  assign \A[7][244] [0] = 1'b1;
  assign \A[7][246] [0] = 1'b1;
  assign \A[7][247] [0] = 1'b1;
  assign \A[7][248] [0] = 1'b1;
  assign \A[7][249] [4] = 1'b1;
  assign \A[7][249] [3] = 1'b1;
  assign \A[7][249] [2] = 1'b1;
  assign \A[7][249] [1] = 1'b1;
  assign \A[7][250] [1] = 1'b1;
  assign \A[7][251] [1] = 1'b1;
  assign \A[7][253] [4] = 1'b1;
  assign \A[7][253] [3] = 1'b1;
  assign \A[7][253] [2] = 1'b1;
  assign \A[7][253] [1] = 1'b1;
  assign \A[7][253] [0] = 1'b1;
  assign \A[7][254] [4] = 1'b1;
  assign \A[7][254] [3] = 1'b1;
  assign \A[7][254] [2] = 1'b1;
  assign \A[7][254] [0] = 1'b1;
  assign \A[7][255] [4] = 1'b1;
  assign \A[7][255] [3] = 1'b1;
  assign \A[7][255] [2] = 1'b1;
  assign \A[7][255] [0] = 1'b1;
  assign \A[8][0] [1] = 1'b1;
  assign \A[8][0] [0] = 1'b1;
  assign \A[8][1] [0] = 1'b1;
  assign \A[8][2] [1] = 1'b1;
  assign \A[8][3] [4] = 1'b1;
  assign \A[8][3] [3] = 1'b1;
  assign \A[8][3] [2] = 1'b1;
  assign \A[8][3] [1] = 1'b1;
  assign \A[8][3] [0] = 1'b1;
  assign \A[8][4] [0] = 1'b1;
  assign \A[8][7] [4] = 1'b1;
  assign \A[8][7] [3] = 1'b1;
  assign \A[8][7] [2] = 1'b1;
  assign \A[8][7] [1] = 1'b1;
  assign \A[8][8] [0] = 1'b1;
  assign \A[8][9] [0] = 1'b1;
  assign \A[8][10] [4] = 1'b1;
  assign \A[8][10] [3] = 1'b1;
  assign \A[8][10] [2] = 1'b1;
  assign \A[8][10] [1] = 1'b1;
  assign \A[8][11] [0] = 1'b1;
  assign \A[8][13] [1] = 1'b1;
  assign \A[8][14] [4] = 1'b1;
  assign \A[8][14] [3] = 1'b1;
  assign \A[8][14] [2] = 1'b1;
  assign \A[8][14] [1] = 1'b1;
  assign \A[8][14] [0] = 1'b1;
  assign \A[8][16] [4] = 1'b1;
  assign \A[8][16] [3] = 1'b1;
  assign \A[8][16] [2] = 1'b1;
  assign \A[8][16] [1] = 1'b1;
  assign \A[8][16] [0] = 1'b1;
  assign \A[8][19] [1] = 1'b1;
  assign \A[8][20] [1] = 1'b1;
  assign \A[8][21] [4] = 1'b1;
  assign \A[8][21] [3] = 1'b1;
  assign \A[8][21] [2] = 1'b1;
  assign \A[8][21] [1] = 1'b1;
  assign \A[8][22] [4] = 1'b1;
  assign \A[8][22] [3] = 1'b1;
  assign \A[8][22] [2] = 1'b1;
  assign \A[8][22] [1] = 1'b1;
  assign \A[8][23] [4] = 1'b1;
  assign \A[8][23] [3] = 1'b1;
  assign \A[8][23] [2] = 1'b1;
  assign \A[8][23] [1] = 1'b1;
  assign \A[8][23] [0] = 1'b1;
  assign \A[8][24] [0] = 1'b1;
  assign \A[8][25] [4] = 1'b1;
  assign \A[8][25] [3] = 1'b1;
  assign \A[8][25] [2] = 1'b1;
  assign \A[8][25] [1] = 1'b1;
  assign \A[8][25] [0] = 1'b1;
  assign \A[8][27] [4] = 1'b1;
  assign \A[8][27] [3] = 1'b1;
  assign \A[8][27] [2] = 1'b1;
  assign \A[8][27] [1] = 1'b1;
  assign \A[8][27] [0] = 1'b1;
  assign \A[8][28] [1] = 1'b1;
  assign \A[8][29] [4] = 1'b1;
  assign \A[8][29] [3] = 1'b1;
  assign \A[8][29] [2] = 1'b1;
  assign \A[8][29] [1] = 1'b1;
  assign \A[8][30] [4] = 1'b1;
  assign \A[8][30] [3] = 1'b1;
  assign \A[8][30] [2] = 1'b1;
  assign \A[8][30] [0] = 1'b1;
  assign \A[8][32] [1] = 1'b1;
  assign \A[8][34] [4] = 1'b1;
  assign \A[8][34] [3] = 1'b1;
  assign \A[8][34] [2] = 1'b1;
  assign \A[8][34] [1] = 1'b1;
  assign \A[8][34] [0] = 1'b1;
  assign \A[8][36] [0] = 1'b1;
  assign \A[8][37] [0] = 1'b1;
  assign \A[8][38] [0] = 1'b1;
  assign \A[8][39] [0] = 1'b1;
  assign \A[8][40] [0] = 1'b1;
  assign \A[8][41] [4] = 1'b1;
  assign \A[8][41] [3] = 1'b1;
  assign \A[8][41] [2] = 1'b1;
  assign \A[8][41] [1] = 1'b1;
  assign \A[8][41] [0] = 1'b1;
  assign \A[8][42] [4] = 1'b1;
  assign \A[8][42] [3] = 1'b1;
  assign \A[8][42] [2] = 1'b1;
  assign \A[8][42] [1] = 1'b1;
  assign \A[8][42] [0] = 1'b1;
  assign \A[8][44] [4] = 1'b1;
  assign \A[8][44] [3] = 1'b1;
  assign \A[8][44] [2] = 1'b1;
  assign \A[8][44] [0] = 1'b1;
  assign \A[8][45] [4] = 1'b1;
  assign \A[8][45] [3] = 1'b1;
  assign \A[8][45] [2] = 1'b1;
  assign \A[8][45] [0] = 1'b1;
  assign \A[8][46] [0] = 1'b1;
  assign \A[8][47] [4] = 1'b1;
  assign \A[8][47] [3] = 1'b1;
  assign \A[8][47] [2] = 1'b1;
  assign \A[8][47] [1] = 1'b1;
  assign \A[8][47] [0] = 1'b1;
  assign \A[8][48] [1] = 1'b1;
  assign \A[8][48] [0] = 1'b1;
  assign \A[8][49] [1] = 1'b1;
  assign \A[8][51] [1] = 1'b1;
  assign \A[8][53] [1] = 1'b1;
  assign \A[8][54] [0] = 1'b1;
  assign \A[8][55] [4] = 1'b1;
  assign \A[8][55] [3] = 1'b1;
  assign \A[8][55] [2] = 1'b1;
  assign \A[8][55] [0] = 1'b1;
  assign \A[8][56] [4] = 1'b1;
  assign \A[8][56] [3] = 1'b1;
  assign \A[8][56] [2] = 1'b1;
  assign \A[8][56] [1] = 1'b1;
  assign \A[8][56] [0] = 1'b1;
  assign \A[8][57] [4] = 1'b1;
  assign \A[8][57] [3] = 1'b1;
  assign \A[8][57] [2] = 1'b1;
  assign \A[8][57] [1] = 1'b1;
  assign \A[8][58] [4] = 1'b1;
  assign \A[8][58] [3] = 1'b1;
  assign \A[8][58] [2] = 1'b1;
  assign \A[8][58] [1] = 1'b1;
  assign \A[8][58] [0] = 1'b1;
  assign \A[8][59] [4] = 1'b1;
  assign \A[8][59] [3] = 1'b1;
  assign \A[8][59] [2] = 1'b1;
  assign \A[8][59] [1] = 1'b1;
  assign \A[8][61] [4] = 1'b1;
  assign \A[8][61] [3] = 1'b1;
  assign \A[8][61] [2] = 1'b1;
  assign \A[8][61] [1] = 1'b1;
  assign \A[8][61] [0] = 1'b1;
  assign \A[8][62] [4] = 1'b1;
  assign \A[8][62] [3] = 1'b1;
  assign \A[8][62] [2] = 1'b1;
  assign \A[8][62] [1] = 1'b1;
  assign \A[8][63] [4] = 1'b1;
  assign \A[8][63] [3] = 1'b1;
  assign \A[8][63] [2] = 1'b1;
  assign \A[8][63] [1] = 1'b1;
  assign \A[8][64] [4] = 1'b1;
  assign \A[8][64] [3] = 1'b1;
  assign \A[8][64] [2] = 1'b1;
  assign \A[8][64] [0] = 1'b1;
  assign \A[8][65] [1] = 1'b1;
  assign \A[8][65] [0] = 1'b1;
  assign \A[8][67] [4] = 1'b1;
  assign \A[8][67] [3] = 1'b1;
  assign \A[8][67] [2] = 1'b1;
  assign \A[8][67] [1] = 1'b1;
  assign \A[8][67] [0] = 1'b1;
  assign \A[8][68] [0] = 1'b1;
  assign \A[8][69] [0] = 1'b1;
  assign \A[8][71] [4] = 1'b1;
  assign \A[8][71] [3] = 1'b1;
  assign \A[8][71] [2] = 1'b1;
  assign \A[8][71] [0] = 1'b1;
  assign \A[8][72] [4] = 1'b1;
  assign \A[8][72] [3] = 1'b1;
  assign \A[8][72] [2] = 1'b1;
  assign \A[8][73] [4] = 1'b1;
  assign \A[8][73] [3] = 1'b1;
  assign \A[8][73] [2] = 1'b1;
  assign \A[8][75] [4] = 1'b1;
  assign \A[8][75] [3] = 1'b1;
  assign \A[8][75] [2] = 1'b1;
  assign \A[8][75] [1] = 1'b1;
  assign \A[8][75] [0] = 1'b1;
  assign \A[8][76] [4] = 1'b1;
  assign \A[8][76] [3] = 1'b1;
  assign \A[8][76] [2] = 1'b1;
  assign \A[8][76] [0] = 1'b1;
  assign \A[8][77] [4] = 1'b1;
  assign \A[8][77] [3] = 1'b1;
  assign \A[8][77] [2] = 1'b1;
  assign \A[8][77] [1] = 1'b1;
  assign \A[8][78] [4] = 1'b1;
  assign \A[8][78] [3] = 1'b1;
  assign \A[8][78] [2] = 1'b1;
  assign \A[8][78] [1] = 1'b1;
  assign \A[8][79] [0] = 1'b1;
  assign \A[8][80] [4] = 1'b1;
  assign \A[8][80] [3] = 1'b1;
  assign \A[8][80] [2] = 1'b1;
  assign \A[8][80] [1] = 1'b1;
  assign \A[8][81] [4] = 1'b1;
  assign \A[8][81] [3] = 1'b1;
  assign \A[8][81] [2] = 1'b1;
  assign \A[8][81] [1] = 1'b1;
  assign \A[8][82] [4] = 1'b1;
  assign \A[8][82] [3] = 1'b1;
  assign \A[8][82] [2] = 1'b1;
  assign \A[8][82] [1] = 1'b1;
  assign \A[8][83] [4] = 1'b1;
  assign \A[8][83] [3] = 1'b1;
  assign \A[8][83] [2] = 1'b1;
  assign \A[8][83] [1] = 1'b1;
  assign \A[8][84] [4] = 1'b1;
  assign \A[8][84] [3] = 1'b1;
  assign \A[8][84] [2] = 1'b1;
  assign \A[8][84] [0] = 1'b1;
  assign \A[8][86] [4] = 1'b1;
  assign \A[8][86] [3] = 1'b1;
  assign \A[8][86] [2] = 1'b1;
  assign \A[8][86] [1] = 1'b1;
  assign \A[8][88] [0] = 1'b1;
  assign \A[8][89] [4] = 1'b1;
  assign \A[8][89] [3] = 1'b1;
  assign \A[8][89] [2] = 1'b1;
  assign \A[8][89] [1] = 1'b1;
  assign \A[8][89] [0] = 1'b1;
  assign \A[8][90] [0] = 1'b1;
  assign \A[8][91] [4] = 1'b1;
  assign \A[8][91] [3] = 1'b1;
  assign \A[8][91] [2] = 1'b1;
  assign \A[8][91] [0] = 1'b1;
  assign \A[8][92] [4] = 1'b1;
  assign \A[8][92] [3] = 1'b1;
  assign \A[8][92] [2] = 1'b1;
  assign \A[8][92] [1] = 1'b1;
  assign \A[8][93] [1] = 1'b1;
  assign \A[8][94] [4] = 1'b1;
  assign \A[8][94] [3] = 1'b1;
  assign \A[8][94] [1] = 1'b1;
  assign \A[8][94] [0] = 1'b1;
  assign \A[8][95] [0] = 1'b1;
  assign \A[8][96] [4] = 1'b1;
  assign \A[8][96] [3] = 1'b1;
  assign \A[8][96] [2] = 1'b1;
  assign \A[8][96] [1] = 1'b1;
  assign \A[8][97] [4] = 1'b1;
  assign \A[8][97] [3] = 1'b1;
  assign \A[8][97] [2] = 1'b1;
  assign \A[8][97] [1] = 1'b1;
  assign \A[8][98] [4] = 1'b1;
  assign \A[8][98] [3] = 1'b1;
  assign \A[8][98] [2] = 1'b1;
  assign \A[8][98] [1] = 1'b1;
  assign \A[8][98] [0] = 1'b1;
  assign \A[8][100] [4] = 1'b1;
  assign \A[8][100] [3] = 1'b1;
  assign \A[8][100] [2] = 1'b1;
  assign \A[8][100] [0] = 1'b1;
  assign \A[8][103] [4] = 1'b1;
  assign \A[8][103] [3] = 1'b1;
  assign \A[8][103] [2] = 1'b1;
  assign \A[8][103] [1] = 1'b1;
  assign \A[8][103] [0] = 1'b1;
  assign \A[8][104] [4] = 1'b1;
  assign \A[8][104] [3] = 1'b1;
  assign \A[8][104] [2] = 1'b1;
  assign \A[8][104] [1] = 1'b1;
  assign \A[8][105] [4] = 1'b1;
  assign \A[8][105] [3] = 1'b1;
  assign \A[8][105] [2] = 1'b1;
  assign \A[8][105] [1] = 1'b1;
  assign \A[8][105] [0] = 1'b1;
  assign \A[8][106] [4] = 1'b1;
  assign \A[8][106] [3] = 1'b1;
  assign \A[8][106] [2] = 1'b1;
  assign \A[8][106] [1] = 1'b1;
  assign \A[8][106] [0] = 1'b1;
  assign \A[8][109] [0] = 1'b1;
  assign \A[8][110] [4] = 1'b1;
  assign \A[8][110] [3] = 1'b1;
  assign \A[8][110] [2] = 1'b1;
  assign \A[8][110] [1] = 1'b1;
  assign \A[8][110] [0] = 1'b1;
  assign \A[8][111] [4] = 1'b1;
  assign \A[8][111] [3] = 1'b1;
  assign \A[8][111] [2] = 1'b1;
  assign \A[8][111] [0] = 1'b1;
  assign \A[8][112] [0] = 1'b1;
  assign \A[8][113] [4] = 1'b1;
  assign \A[8][113] [3] = 1'b1;
  assign \A[8][113] [2] = 1'b1;
  assign \A[8][113] [1] = 1'b1;
  assign \A[8][114] [4] = 1'b1;
  assign \A[8][114] [3] = 1'b1;
  assign \A[8][114] [2] = 1'b1;
  assign \A[8][114] [1] = 1'b1;
  assign \A[8][115] [0] = 1'b1;
  assign \A[8][117] [0] = 1'b1;
  assign \A[8][118] [4] = 1'b1;
  assign \A[8][118] [3] = 1'b1;
  assign \A[8][118] [2] = 1'b1;
  assign \A[8][118] [1] = 1'b1;
  assign \A[8][119] [0] = 1'b1;
  assign \A[8][120] [4] = 1'b1;
  assign \A[8][120] [3] = 1'b1;
  assign \A[8][120] [2] = 1'b1;
  assign \A[8][120] [1] = 1'b1;
  assign \A[8][121] [4] = 1'b1;
  assign \A[8][121] [3] = 1'b1;
  assign \A[8][121] [2] = 1'b1;
  assign \A[8][121] [1] = 1'b1;
  assign \A[8][121] [0] = 1'b1;
  assign \A[8][122] [0] = 1'b1;
  assign \A[8][124] [0] = 1'b1;
  assign \A[8][125] [4] = 1'b1;
  assign \A[8][125] [3] = 1'b1;
  assign \A[8][125] [2] = 1'b1;
  assign \A[8][125] [1] = 1'b1;
  assign \A[8][126] [4] = 1'b1;
  assign \A[8][126] [3] = 1'b1;
  assign \A[8][126] [2] = 1'b1;
  assign \A[8][126] [1] = 1'b1;
  assign \A[8][126] [0] = 1'b1;
  assign \A[8][128] [1] = 1'b1;
  assign \A[8][129] [0] = 1'b1;
  assign \A[8][130] [0] = 1'b1;
  assign \A[8][131] [1] = 1'b1;
  assign \A[8][131] [0] = 1'b1;
  assign \A[8][132] [4] = 1'b1;
  assign \A[8][132] [3] = 1'b1;
  assign \A[8][132] [2] = 1'b1;
  assign \A[8][132] [1] = 1'b1;
  assign \A[8][134] [0] = 1'b1;
  assign \A[8][136] [0] = 1'b1;
  assign \A[8][137] [4] = 1'b1;
  assign \A[8][137] [3] = 1'b1;
  assign \A[8][137] [2] = 1'b1;
  assign \A[8][137] [0] = 1'b1;
  assign \A[8][138] [0] = 1'b1;
  assign \A[8][139] [4] = 1'b1;
  assign \A[8][139] [3] = 1'b1;
  assign \A[8][139] [2] = 1'b1;
  assign \A[8][139] [1] = 1'b1;
  assign \A[8][139] [0] = 1'b1;
  assign \A[8][140] [4] = 1'b1;
  assign \A[8][140] [3] = 1'b1;
  assign \A[8][140] [2] = 1'b1;
  assign \A[8][140] [1] = 1'b1;
  assign \A[8][141] [0] = 1'b1;
  assign \A[8][142] [4] = 1'b1;
  assign \A[8][142] [3] = 1'b1;
  assign \A[8][142] [2] = 1'b1;
  assign \A[8][142] [1] = 1'b1;
  assign \A[8][143] [1] = 1'b1;
  assign \A[8][144] [0] = 1'b1;
  assign \A[8][145] [1] = 1'b1;
  assign \A[8][146] [0] = 1'b1;
  assign \A[8][147] [1] = 1'b1;
  assign \A[8][148] [1] = 1'b1;
  assign \A[8][148] [0] = 1'b1;
  assign \A[8][149] [0] = 1'b1;
  assign \A[8][150] [4] = 1'b1;
  assign \A[8][150] [3] = 1'b1;
  assign \A[8][150] [2] = 1'b1;
  assign \A[8][150] [1] = 1'b1;
  assign \A[8][151] [4] = 1'b1;
  assign \A[8][151] [3] = 1'b1;
  assign \A[8][151] [2] = 1'b1;
  assign \A[8][151] [1] = 1'b1;
  assign \A[8][151] [0] = 1'b1;
  assign \A[8][152] [1] = 1'b1;
  assign \A[8][154] [1] = 1'b1;
  assign \A[8][156] [0] = 1'b1;
  assign \A[8][157] [0] = 1'b1;
  assign \A[8][158] [4] = 1'b1;
  assign \A[8][158] [3] = 1'b1;
  assign \A[8][158] [2] = 1'b1;
  assign \A[8][159] [4] = 1'b1;
  assign \A[8][159] [3] = 1'b1;
  assign \A[8][159] [2] = 1'b1;
  assign \A[8][159] [1] = 1'b1;
  assign \A[8][159] [0] = 1'b1;
  assign \A[8][160] [1] = 1'b1;
  assign \A[8][161] [2] = 1'b1;
  assign \A[8][162] [1] = 1'b1;
  assign \A[8][162] [0] = 1'b1;
  assign \A[8][163] [0] = 1'b1;
  assign \A[8][164] [1] = 1'b1;
  assign \A[8][164] [0] = 1'b1;
  assign \A[8][165] [0] = 1'b1;
  assign \A[8][166] [2] = 1'b1;
  assign \A[8][168] [0] = 1'b1;
  assign \A[8][169] [1] = 1'b1;
  assign \A[8][170] [4] = 1'b1;
  assign \A[8][170] [3] = 1'b1;
  assign \A[8][170] [2] = 1'b1;
  assign \A[8][170] [1] = 1'b1;
  assign \A[8][170] [0] = 1'b1;
  assign \A[8][171] [4] = 1'b1;
  assign \A[8][171] [3] = 1'b1;
  assign \A[8][171] [2] = 1'b1;
  assign \A[8][171] [1] = 1'b1;
  assign \A[8][171] [0] = 1'b1;
  assign \A[8][172] [4] = 1'b1;
  assign \A[8][172] [3] = 1'b1;
  assign \A[8][172] [2] = 1'b1;
  assign \A[8][172] [1] = 1'b1;
  assign \A[8][172] [0] = 1'b1;
  assign \A[8][173] [4] = 1'b1;
  assign \A[8][173] [3] = 1'b1;
  assign \A[8][173] [2] = 1'b1;
  assign \A[8][173] [1] = 1'b1;
  assign \A[8][175] [0] = 1'b1;
  assign \A[8][176] [4] = 1'b1;
  assign \A[8][176] [3] = 1'b1;
  assign \A[8][176] [2] = 1'b1;
  assign \A[8][176] [1] = 1'b1;
  assign \A[8][176] [0] = 1'b1;
  assign \A[8][177] [2] = 1'b1;
  assign \A[8][178] [0] = 1'b1;
  assign \A[8][179] [1] = 1'b1;
  assign \A[8][180] [1] = 1'b1;
  assign \A[8][180] [0] = 1'b1;
  assign \A[8][181] [1] = 1'b1;
  assign \A[8][181] [0] = 1'b1;
  assign \A[8][182] [1] = 1'b1;
  assign \A[8][182] [0] = 1'b1;
  assign \A[8][184] [4] = 1'b1;
  assign \A[8][184] [3] = 1'b1;
  assign \A[8][184] [2] = 1'b1;
  assign \A[8][184] [1] = 1'b1;
  assign \A[8][186] [4] = 1'b1;
  assign \A[8][186] [3] = 1'b1;
  assign \A[8][186] [2] = 1'b1;
  assign \A[8][186] [1] = 1'b1;
  assign \A[8][186] [0] = 1'b1;
  assign \A[8][187] [4] = 1'b1;
  assign \A[8][187] [3] = 1'b1;
  assign \A[8][187] [2] = 1'b1;
  assign \A[8][187] [1] = 1'b1;
  assign \A[8][188] [4] = 1'b1;
  assign \A[8][188] [3] = 1'b1;
  assign \A[8][188] [2] = 1'b1;
  assign \A[8][190] [4] = 1'b1;
  assign \A[8][190] [3] = 1'b1;
  assign \A[8][190] [2] = 1'b1;
  assign \A[8][190] [1] = 1'b1;
  assign \A[8][191] [4] = 1'b1;
  assign \A[8][191] [3] = 1'b1;
  assign \A[8][191] [2] = 1'b1;
  assign \A[8][191] [0] = 1'b1;
  assign \A[8][192] [0] = 1'b1;
  assign \A[8][193] [2] = 1'b1;
  assign \A[8][195] [1] = 1'b1;
  assign \A[8][195] [0] = 1'b1;
  assign \A[8][196] [0] = 1'b1;
  assign \A[8][197] [0] = 1'b1;
  assign \A[8][198] [1] = 1'b1;
  assign \A[8][198] [0] = 1'b1;
  assign \A[8][199] [4] = 1'b1;
  assign \A[8][199] [3] = 1'b1;
  assign \A[8][199] [2] = 1'b1;
  assign \A[8][199] [1] = 1'b1;
  assign \A[8][199] [0] = 1'b1;
  assign \A[8][200] [1] = 1'b1;
  assign \A[8][201] [0] = 1'b1;
  assign \A[8][203] [4] = 1'b1;
  assign \A[8][203] [3] = 1'b1;
  assign \A[8][203] [2] = 1'b1;
  assign \A[8][203] [1] = 1'b1;
  assign \A[8][203] [0] = 1'b1;
  assign \A[8][204] [1] = 1'b1;
  assign \A[8][205] [4] = 1'b1;
  assign \A[8][205] [3] = 1'b1;
  assign \A[8][205] [2] = 1'b1;
  assign \A[8][205] [1] = 1'b1;
  assign \A[8][206] [4] = 1'b1;
  assign \A[8][206] [3] = 1'b1;
  assign \A[8][206] [2] = 1'b1;
  assign \A[8][206] [1] = 1'b1;
  assign \A[8][206] [0] = 1'b1;
  assign \A[8][207] [0] = 1'b1;
  assign \A[8][208] [2] = 1'b1;
  assign \A[8][209] [0] = 1'b1;
  assign \A[8][210] [4] = 1'b1;
  assign \A[8][210] [3] = 1'b1;
  assign \A[8][210] [2] = 1'b1;
  assign \A[8][210] [1] = 1'b1;
  assign \A[8][210] [0] = 1'b1;
  assign \A[8][211] [0] = 1'b1;
  assign \A[8][215] [4] = 1'b1;
  assign \A[8][215] [3] = 1'b1;
  assign \A[8][215] [2] = 1'b1;
  assign \A[8][215] [1] = 1'b1;
  assign \A[8][215] [0] = 1'b1;
  assign \A[8][216] [0] = 1'b1;
  assign \A[8][218] [0] = 1'b1;
  assign \A[8][220] [4] = 1'b1;
  assign \A[8][220] [3] = 1'b1;
  assign \A[8][220] [2] = 1'b1;
  assign \A[8][220] [1] = 1'b1;
  assign \A[8][220] [0] = 1'b1;
  assign \A[8][221] [4] = 1'b1;
  assign \A[8][221] [3] = 1'b1;
  assign \A[8][221] [2] = 1'b1;
  assign \A[8][221] [1] = 1'b1;
  assign \A[8][221] [0] = 1'b1;
  assign \A[8][222] [4] = 1'b1;
  assign \A[8][222] [3] = 1'b1;
  assign \A[8][222] [2] = 1'b1;
  assign \A[8][222] [1] = 1'b1;
  assign \A[8][222] [0] = 1'b1;
  assign \A[8][223] [4] = 1'b1;
  assign \A[8][223] [3] = 1'b1;
  assign \A[8][223] [2] = 1'b1;
  assign \A[8][223] [0] = 1'b1;
  assign \A[8][224] [0] = 1'b1;
  assign \A[8][225] [4] = 1'b1;
  assign \A[8][225] [3] = 1'b1;
  assign \A[8][225] [2] = 1'b1;
  assign \A[8][225] [1] = 1'b1;
  assign \A[8][225] [0] = 1'b1;
  assign \A[8][226] [0] = 1'b1;
  assign \A[8][227] [0] = 1'b1;
  assign \A[8][228] [4] = 1'b1;
  assign \A[8][228] [3] = 1'b1;
  assign \A[8][228] [2] = 1'b1;
  assign \A[8][228] [1] = 1'b1;
  assign \A[8][228] [0] = 1'b1;
  assign \A[8][229] [0] = 1'b1;
  assign \A[8][230] [1] = 1'b1;
  assign \A[8][230] [0] = 1'b1;
  assign \A[8][231] [4] = 1'b1;
  assign \A[8][231] [3] = 1'b1;
  assign \A[8][231] [2] = 1'b1;
  assign \A[8][231] [1] = 1'b1;
  assign \A[8][232] [4] = 1'b1;
  assign \A[8][232] [3] = 1'b1;
  assign \A[8][232] [2] = 1'b1;
  assign \A[8][232] [1] = 1'b1;
  assign \A[8][232] [0] = 1'b1;
  assign \A[8][233] [0] = 1'b1;
  assign \A[8][234] [0] = 1'b1;
  assign \A[8][235] [4] = 1'b1;
  assign \A[8][235] [3] = 1'b1;
  assign \A[8][235] [2] = 1'b1;
  assign \A[8][235] [1] = 1'b1;
  assign \A[8][236] [0] = 1'b1;
  assign \A[8][237] [4] = 1'b1;
  assign \A[8][237] [3] = 1'b1;
  assign \A[8][237] [2] = 1'b1;
  assign \A[8][237] [1] = 1'b1;
  assign \A[8][237] [0] = 1'b1;
  assign \A[8][238] [4] = 1'b1;
  assign \A[8][238] [3] = 1'b1;
  assign \A[8][238] [2] = 1'b1;
  assign \A[8][238] [1] = 1'b1;
  assign \A[8][239] [1] = 1'b1;
  assign \A[8][240] [4] = 1'b1;
  assign \A[8][240] [3] = 1'b1;
  assign \A[8][240] [2] = 1'b1;
  assign \A[8][240] [0] = 1'b1;
  assign \A[8][241] [0] = 1'b1;
  assign \A[8][243] [4] = 1'b1;
  assign \A[8][243] [3] = 1'b1;
  assign \A[8][243] [2] = 1'b1;
  assign \A[8][243] [1] = 1'b1;
  assign \A[8][247] [1] = 1'b1;
  assign \A[8][250] [1] = 1'b1;
  assign \A[8][251] [0] = 1'b1;
  assign \A[8][252] [4] = 1'b1;
  assign \A[8][252] [3] = 1'b1;
  assign \A[8][252] [2] = 1'b1;
  assign \A[8][252] [1] = 1'b1;
  assign \A[8][252] [0] = 1'b1;
  assign \A[8][253] [2] = 1'b1;
  assign \A[9][0] [2] = 1'b1;
  assign \A[9][2] [1] = 1'b1;
  assign \A[9][3] [1] = 1'b1;
  assign \A[9][3] [0] = 1'b1;
  assign \A[9][4] [4] = 1'b1;
  assign \A[9][4] [3] = 1'b1;
  assign \A[9][4] [2] = 1'b1;
  assign \A[9][4] [1] = 1'b1;
  assign \A[9][4] [0] = 1'b1;
  assign \A[9][5] [1] = 1'b1;
  assign \A[9][6] [4] = 1'b1;
  assign \A[9][6] [3] = 1'b1;
  assign \A[9][6] [2] = 1'b1;
  assign \A[9][6] [1] = 1'b1;
  assign \A[9][7] [2] = 1'b1;
  assign \A[9][7] [0] = 1'b1;
  assign \A[9][8] [0] = 1'b1;
  assign \A[9][10] [0] = 1'b1;
  assign \A[9][11] [4] = 1'b1;
  assign \A[9][11] [3] = 1'b1;
  assign \A[9][11] [2] = 1'b1;
  assign \A[9][11] [1] = 1'b1;
  assign \A[9][11] [0] = 1'b1;
  assign \A[9][14] [4] = 1'b1;
  assign \A[9][14] [3] = 1'b1;
  assign \A[9][14] [2] = 1'b1;
  assign \A[9][14] [1] = 1'b1;
  assign \A[9][14] [0] = 1'b1;
  assign \A[9][16] [1] = 1'b1;
  assign \A[9][17] [1] = 1'b1;
  assign \A[9][18] [4] = 1'b1;
  assign \A[9][18] [3] = 1'b1;
  assign \A[9][18] [2] = 1'b1;
  assign \A[9][18] [1] = 1'b1;
  assign \A[9][19] [1] = 1'b1;
  assign \A[9][21] [0] = 1'b1;
  assign \A[9][22] [0] = 1'b1;
  assign \A[9][25] [4] = 1'b1;
  assign \A[9][25] [3] = 1'b1;
  assign \A[9][25] [2] = 1'b1;
  assign \A[9][25] [1] = 1'b1;
  assign \A[9][26] [4] = 1'b1;
  assign \A[9][26] [3] = 1'b1;
  assign \A[9][26] [2] = 1'b1;
  assign \A[9][26] [1] = 1'b1;
  assign \A[9][26] [0] = 1'b1;
  assign \A[9][29] [4] = 1'b1;
  assign \A[9][29] [3] = 1'b1;
  assign \A[9][29] [2] = 1'b1;
  assign \A[9][29] [1] = 1'b1;
  assign \A[9][30] [2] = 1'b1;
  assign \A[9][32] [4] = 1'b1;
  assign \A[9][32] [3] = 1'b1;
  assign \A[9][32] [2] = 1'b1;
  assign \A[9][32] [1] = 1'b1;
  assign \A[9][32] [0] = 1'b1;
  assign \A[9][33] [1] = 1'b1;
  assign \A[9][34] [0] = 1'b1;
  assign \A[9][36] [0] = 1'b1;
  assign \A[9][38] [1] = 1'b1;
  assign \A[9][39] [1] = 1'b1;
  assign \A[9][42] [4] = 1'b1;
  assign \A[9][42] [3] = 1'b1;
  assign \A[9][42] [2] = 1'b1;
  assign \A[9][42] [1] = 1'b1;
  assign \A[9][42] [0] = 1'b1;
  assign \A[9][43] [1] = 1'b1;
  assign \A[9][45] [1] = 1'b1;
  assign \A[9][46] [1] = 1'b1;
  assign \A[9][47] [1] = 1'b1;
  assign \A[9][48] [4] = 1'b1;
  assign \A[9][48] [3] = 1'b1;
  assign \A[9][48] [2] = 1'b1;
  assign \A[9][48] [1] = 1'b1;
  assign \A[9][48] [0] = 1'b1;
  assign \A[9][49] [4] = 1'b1;
  assign \A[9][49] [3] = 1'b1;
  assign \A[9][49] [2] = 1'b1;
  assign \A[9][49] [1] = 1'b1;
  assign \A[9][50] [1] = 1'b1;
  assign \A[9][52] [4] = 1'b1;
  assign \A[9][52] [3] = 1'b1;
  assign \A[9][52] [2] = 1'b1;
  assign \A[9][52] [1] = 1'b1;
  assign \A[9][54] [4] = 1'b1;
  assign \A[9][54] [3] = 1'b1;
  assign \A[9][54] [2] = 1'b1;
  assign \A[9][54] [1] = 1'b1;
  assign \A[9][54] [0] = 1'b1;
  assign \A[9][55] [0] = 1'b1;
  assign \A[9][56] [1] = 1'b1;
  assign \A[9][57] [1] = 1'b1;
  assign \A[9][58] [4] = 1'b1;
  assign \A[9][58] [3] = 1'b1;
  assign \A[9][58] [2] = 1'b1;
  assign \A[9][58] [1] = 1'b1;
  assign \A[9][58] [0] = 1'b1;
  assign \A[9][60] [1] = 1'b1;
  assign \A[9][61] [0] = 1'b1;
  assign \A[9][62] [1] = 1'b1;
  assign \A[9][64] [4] = 1'b1;
  assign \A[9][64] [3] = 1'b1;
  assign \A[9][64] [2] = 1'b1;
  assign \A[9][64] [1] = 1'b1;
  assign \A[9][64] [0] = 1'b1;
  assign \A[9][65] [4] = 1'b1;
  assign \A[9][65] [3] = 1'b1;
  assign \A[9][65] [2] = 1'b1;
  assign \A[9][65] [0] = 1'b1;
  assign \A[9][66] [4] = 1'b1;
  assign \A[9][66] [3] = 1'b1;
  assign \A[9][66] [2] = 1'b1;
  assign \A[9][66] [1] = 1'b1;
  assign \A[9][68] [4] = 1'b1;
  assign \A[9][68] [3] = 1'b1;
  assign \A[9][68] [2] = 1'b1;
  assign \A[9][68] [1] = 1'b1;
  assign \A[9][68] [0] = 1'b1;
  assign \A[9][69] [0] = 1'b1;
  assign \A[9][70] [4] = 1'b1;
  assign \A[9][70] [3] = 1'b1;
  assign \A[9][70] [2] = 1'b1;
  assign \A[9][70] [1] = 1'b1;
  assign \A[9][71] [1] = 1'b1;
  assign \A[9][72] [1] = 1'b1;
  assign \A[9][72] [0] = 1'b1;
  assign \A[9][74] [1] = 1'b1;
  assign \A[9][74] [0] = 1'b1;
  assign \A[9][75] [0] = 1'b1;
  assign \A[9][76] [1] = 1'b1;
  assign \A[9][76] [0] = 1'b1;
  assign \A[9][77] [1] = 1'b1;
  assign \A[9][79] [0] = 1'b1;
  assign \A[9][80] [4] = 1'b1;
  assign \A[9][80] [3] = 1'b1;
  assign \A[9][80] [2] = 1'b1;
  assign \A[9][80] [1] = 1'b1;
  assign \A[9][81] [4] = 1'b1;
  assign \A[9][81] [3] = 1'b1;
  assign \A[9][81] [2] = 1'b1;
  assign \A[9][81] [1] = 1'b1;
  assign \A[9][82] [1] = 1'b1;
  assign \A[9][82] [0] = 1'b1;
  assign \A[9][84] [4] = 1'b1;
  assign \A[9][84] [3] = 1'b1;
  assign \A[9][84] [2] = 1'b1;
  assign \A[9][84] [1] = 1'b1;
  assign \A[9][86] [1] = 1'b1;
  assign \A[9][87] [0] = 1'b1;
  assign \A[9][88] [0] = 1'b1;
  assign \A[9][91] [4] = 1'b1;
  assign \A[9][91] [3] = 1'b1;
  assign \A[9][91] [2] = 1'b1;
  assign \A[9][91] [1] = 1'b1;
  assign \A[9][91] [0] = 1'b1;
  assign \A[9][93] [4] = 1'b1;
  assign \A[9][93] [3] = 1'b1;
  assign \A[9][93] [2] = 1'b1;
  assign \A[9][93] [1] = 1'b1;
  assign \A[9][94] [4] = 1'b1;
  assign \A[9][94] [3] = 1'b1;
  assign \A[9][94] [2] = 1'b1;
  assign \A[9][94] [1] = 1'b1;
  assign \A[9][95] [0] = 1'b1;
  assign \A[9][97] [4] = 1'b1;
  assign \A[9][97] [3] = 1'b1;
  assign \A[9][97] [2] = 1'b1;
  assign \A[9][97] [1] = 1'b1;
  assign \A[9][98] [4] = 1'b1;
  assign \A[9][98] [3] = 1'b1;
  assign \A[9][98] [2] = 1'b1;
  assign \A[9][98] [0] = 1'b1;
  assign \A[9][100] [1] = 1'b1;
  assign \A[9][101] [1] = 1'b1;
  assign \A[9][102] [0] = 1'b1;
  assign \A[9][103] [0] = 1'b1;
  assign \A[9][105] [0] = 1'b1;
  assign \A[9][106] [0] = 1'b1;
  assign \A[9][108] [1] = 1'b1;
  assign \A[9][110] [4] = 1'b1;
  assign \A[9][110] [3] = 1'b1;
  assign \A[9][110] [2] = 1'b1;
  assign \A[9][110] [1] = 1'b1;
  assign \A[9][113] [1] = 1'b1;
  assign \A[9][114] [0] = 1'b1;
  assign \A[9][116] [0] = 1'b1;
  assign \A[9][118] [0] = 1'b1;
  assign \A[9][119] [0] = 1'b1;
  assign \A[9][120] [1] = 1'b1;
  assign \A[9][121] [0] = 1'b1;
  assign \A[9][123] [1] = 1'b1;
  assign \A[9][124] [1] = 1'b1;
  assign \A[9][124] [0] = 1'b1;
  assign \A[9][126] [4] = 1'b1;
  assign \A[9][126] [3] = 1'b1;
  assign \A[9][126] [2] = 1'b1;
  assign \A[9][126] [1] = 1'b1;
  assign \A[9][127] [0] = 1'b1;
  assign \A[9][128] [4] = 1'b1;
  assign \A[9][128] [3] = 1'b1;
  assign \A[9][128] [2] = 1'b1;
  assign \A[9][128] [1] = 1'b1;
  assign \A[9][129] [4] = 1'b1;
  assign \A[9][129] [3] = 1'b1;
  assign \A[9][129] [2] = 1'b1;
  assign \A[9][129] [1] = 1'b1;
  assign \A[9][130] [0] = 1'b1;
  assign \A[9][131] [0] = 1'b1;
  assign \A[9][133] [4] = 1'b1;
  assign \A[9][133] [3] = 1'b1;
  assign \A[9][133] [2] = 1'b1;
  assign \A[9][133] [1] = 1'b1;
  assign \A[9][133] [0] = 1'b1;
  assign \A[9][134] [1] = 1'b1;
  assign \A[9][135] [4] = 1'b1;
  assign \A[9][135] [3] = 1'b1;
  assign \A[9][135] [2] = 1'b1;
  assign \A[9][135] [1] = 1'b1;
  assign \A[9][135] [0] = 1'b1;
  assign \A[9][137] [1] = 1'b1;
  assign \A[9][138] [0] = 1'b1;
  assign \A[9][139] [0] = 1'b1;
  assign \A[9][140] [4] = 1'b1;
  assign \A[9][140] [3] = 1'b1;
  assign \A[9][140] [2] = 1'b1;
  assign \A[9][140] [1] = 1'b1;
  assign \A[9][140] [0] = 1'b1;
  assign \A[9][141] [0] = 1'b1;
  assign \A[9][143] [1] = 1'b1;
  assign \A[9][143] [0] = 1'b1;
  assign \A[9][146] [4] = 1'b1;
  assign \A[9][146] [3] = 1'b1;
  assign \A[9][146] [2] = 1'b1;
  assign \A[9][146] [0] = 1'b1;
  assign \A[9][148] [4] = 1'b1;
  assign \A[9][148] [3] = 1'b1;
  assign \A[9][148] [2] = 1'b1;
  assign \A[9][148] [1] = 1'b1;
  assign \A[9][149] [1] = 1'b1;
  assign \A[9][150] [0] = 1'b1;
  assign \A[9][151] [0] = 1'b1;
  assign \A[9][152] [4] = 1'b1;
  assign \A[9][152] [3] = 1'b1;
  assign \A[9][152] [2] = 1'b1;
  assign \A[9][152] [1] = 1'b1;
  assign \A[9][152] [0] = 1'b1;
  assign \A[9][153] [1] = 1'b1;
  assign \A[9][154] [0] = 1'b1;
  assign \A[9][155] [0] = 1'b1;
  assign \A[9][156] [1] = 1'b1;
  assign \A[9][156] [0] = 1'b1;
  assign \A[9][157] [4] = 1'b1;
  assign \A[9][157] [3] = 1'b1;
  assign \A[9][157] [2] = 1'b1;
  assign \A[9][157] [1] = 1'b1;
  assign \A[9][157] [0] = 1'b1;
  assign \A[9][159] [1] = 1'b1;
  assign \A[9][159] [0] = 1'b1;
  assign \A[9][161] [4] = 1'b1;
  assign \A[9][161] [3] = 1'b1;
  assign \A[9][161] [2] = 1'b1;
  assign \A[9][161] [1] = 1'b1;
  assign \A[9][161] [0] = 1'b1;
  assign \A[9][163] [4] = 1'b1;
  assign \A[9][163] [3] = 1'b1;
  assign \A[9][163] [2] = 1'b1;
  assign \A[9][163] [0] = 1'b1;
  assign \A[9][164] [4] = 1'b1;
  assign \A[9][164] [3] = 1'b1;
  assign \A[9][164] [2] = 1'b1;
  assign \A[9][164] [1] = 1'b1;
  assign \A[9][164] [0] = 1'b1;
  assign \A[9][166] [0] = 1'b1;
  assign \A[9][168] [1] = 1'b1;
  assign \A[9][169] [4] = 1'b1;
  assign \A[9][169] [3] = 1'b1;
  assign \A[9][169] [2] = 1'b1;
  assign \A[9][169] [1] = 1'b1;
  assign \A[9][170] [0] = 1'b1;
  assign \A[9][172] [0] = 1'b1;
  assign \A[9][173] [1] = 1'b1;
  assign \A[9][174] [0] = 1'b1;
  assign \A[9][175] [1] = 1'b1;
  assign \A[9][176] [4] = 1'b1;
  assign \A[9][176] [3] = 1'b1;
  assign \A[9][176] [2] = 1'b1;
  assign \A[9][176] [0] = 1'b1;
  assign \A[9][177] [4] = 1'b1;
  assign \A[9][177] [3] = 1'b1;
  assign \A[9][177] [2] = 1'b1;
  assign \A[9][177] [1] = 1'b1;
  assign \A[9][178] [4] = 1'b1;
  assign \A[9][178] [3] = 1'b1;
  assign \A[9][178] [2] = 1'b1;
  assign \A[9][178] [1] = 1'b1;
  assign \A[9][178] [0] = 1'b1;
  assign \A[9][179] [4] = 1'b1;
  assign \A[9][179] [3] = 1'b1;
  assign \A[9][179] [2] = 1'b1;
  assign \A[9][179] [1] = 1'b1;
  assign \A[9][179] [0] = 1'b1;
  assign \A[9][180] [0] = 1'b1;
  assign \A[9][181] [4] = 1'b1;
  assign \A[9][181] [3] = 1'b1;
  assign \A[9][181] [2] = 1'b1;
  assign \A[9][181] [1] = 1'b1;
  assign \A[9][182] [4] = 1'b1;
  assign \A[9][182] [3] = 1'b1;
  assign \A[9][182] [2] = 1'b1;
  assign \A[9][183] [1] = 1'b1;
  assign \A[9][184] [1] = 1'b1;
  assign \A[9][185] [0] = 1'b1;
  assign \A[9][187] [4] = 1'b1;
  assign \A[9][187] [3] = 1'b1;
  assign \A[9][187] [2] = 1'b1;
  assign \A[9][187] [1] = 1'b1;
  assign \A[9][188] [4] = 1'b1;
  assign \A[9][188] [3] = 1'b1;
  assign \A[9][188] [2] = 1'b1;
  assign \A[9][188] [1] = 1'b1;
  assign \A[9][188] [0] = 1'b1;
  assign \A[9][190] [4] = 1'b1;
  assign \A[9][190] [3] = 1'b1;
  assign \A[9][190] [2] = 1'b1;
  assign \A[9][190] [1] = 1'b1;
  assign \A[9][190] [0] = 1'b1;
  assign \A[9][191] [0] = 1'b1;
  assign \A[9][192] [4] = 1'b1;
  assign \A[9][192] [3] = 1'b1;
  assign \A[9][192] [2] = 1'b1;
  assign \A[9][192] [1] = 1'b1;
  assign \A[9][193] [4] = 1'b1;
  assign \A[9][193] [3] = 1'b1;
  assign \A[9][193] [2] = 1'b1;
  assign \A[9][193] [1] = 1'b1;
  assign \A[9][195] [4] = 1'b1;
  assign \A[9][195] [3] = 1'b1;
  assign \A[9][195] [2] = 1'b1;
  assign \A[9][195] [1] = 1'b1;
  assign \A[9][195] [0] = 1'b1;
  assign \A[9][196] [4] = 1'b1;
  assign \A[9][196] [3] = 1'b1;
  assign \A[9][196] [2] = 1'b1;
  assign \A[9][196] [1] = 1'b1;
  assign \A[9][196] [0] = 1'b1;
  assign \A[9][197] [1] = 1'b1;
  assign \A[9][197] [0] = 1'b1;
  assign \A[9][198] [4] = 1'b1;
  assign \A[9][198] [3] = 1'b1;
  assign \A[9][198] [2] = 1'b1;
  assign \A[9][198] [1] = 1'b1;
  assign \A[9][198] [0] = 1'b1;
  assign \A[9][199] [4] = 1'b1;
  assign \A[9][199] [3] = 1'b1;
  assign \A[9][199] [2] = 1'b1;
  assign \A[9][199] [1] = 1'b1;
  assign \A[9][200] [4] = 1'b1;
  assign \A[9][200] [3] = 1'b1;
  assign \A[9][200] [2] = 1'b1;
  assign \A[9][200] [1] = 1'b1;
  assign \A[9][201] [4] = 1'b1;
  assign \A[9][201] [3] = 1'b1;
  assign \A[9][201] [2] = 1'b1;
  assign \A[9][201] [1] = 1'b1;
  assign \A[9][201] [0] = 1'b1;
  assign \A[9][202] [4] = 1'b1;
  assign \A[9][202] [3] = 1'b1;
  assign \A[9][202] [2] = 1'b1;
  assign \A[9][202] [1] = 1'b1;
  assign \A[9][203] [0] = 1'b1;
  assign \A[9][204] [4] = 1'b1;
  assign \A[9][204] [3] = 1'b1;
  assign \A[9][204] [2] = 1'b1;
  assign \A[9][204] [1] = 1'b1;
  assign \A[9][204] [0] = 1'b1;
  assign \A[9][205] [0] = 1'b1;
  assign \A[9][206] [4] = 1'b1;
  assign \A[9][206] [3] = 1'b1;
  assign \A[9][206] [2] = 1'b1;
  assign \A[9][206] [1] = 1'b1;
  assign \A[9][206] [0] = 1'b1;
  assign \A[9][208] [4] = 1'b1;
  assign \A[9][208] [3] = 1'b1;
  assign \A[9][208] [2] = 1'b1;
  assign \A[9][208] [1] = 1'b1;
  assign \A[9][208] [0] = 1'b1;
  assign \A[9][209] [1] = 1'b1;
  assign \A[9][209] [0] = 1'b1;
  assign \A[9][210] [4] = 1'b1;
  assign \A[9][210] [3] = 1'b1;
  assign \A[9][210] [2] = 1'b1;
  assign \A[9][210] [1] = 1'b1;
  assign \A[9][211] [4] = 1'b1;
  assign \A[9][211] [3] = 1'b1;
  assign \A[9][211] [2] = 1'b1;
  assign \A[9][211] [1] = 1'b1;
  assign \A[9][212] [4] = 1'b1;
  assign \A[9][212] [3] = 1'b1;
  assign \A[9][212] [2] = 1'b1;
  assign \A[9][212] [1] = 1'b1;
  assign \A[9][213] [4] = 1'b1;
  assign \A[9][213] [3] = 1'b1;
  assign \A[9][213] [2] = 1'b1;
  assign \A[9][213] [1] = 1'b1;
  assign \A[9][214] [4] = 1'b1;
  assign \A[9][214] [3] = 1'b1;
  assign \A[9][214] [2] = 1'b1;
  assign \A[9][214] [1] = 1'b1;
  assign \A[9][215] [4] = 1'b1;
  assign \A[9][215] [3] = 1'b1;
  assign \A[9][215] [2] = 1'b1;
  assign \A[9][215] [1] = 1'b1;
  assign \A[9][216] [4] = 1'b1;
  assign \A[9][216] [3] = 1'b1;
  assign \A[9][216] [2] = 1'b1;
  assign \A[9][216] [1] = 1'b1;
  assign \A[9][216] [0] = 1'b1;
  assign \A[9][217] [4] = 1'b1;
  assign \A[9][217] [3] = 1'b1;
  assign \A[9][217] [2] = 1'b1;
  assign \A[9][217] [0] = 1'b1;
  assign \A[9][218] [4] = 1'b1;
  assign \A[9][218] [3] = 1'b1;
  assign \A[9][218] [2] = 1'b1;
  assign \A[9][218] [1] = 1'b1;
  assign \A[9][218] [0] = 1'b1;
  assign \A[9][219] [1] = 1'b1;
  assign \A[9][220] [4] = 1'b1;
  assign \A[9][220] [3] = 1'b1;
  assign \A[9][220] [2] = 1'b1;
  assign \A[9][220] [1] = 1'b1;
  assign \A[9][220] [0] = 1'b1;
  assign \A[9][221] [4] = 1'b1;
  assign \A[9][221] [3] = 1'b1;
  assign \A[9][221] [2] = 1'b1;
  assign \A[9][221] [0] = 1'b1;
  assign \A[9][222] [0] = 1'b1;
  assign \A[9][223] [4] = 1'b1;
  assign \A[9][223] [3] = 1'b1;
  assign \A[9][223] [2] = 1'b1;
  assign \A[9][223] [1] = 1'b1;
  assign \A[9][223] [0] = 1'b1;
  assign \A[9][224] [0] = 1'b1;
  assign \A[9][225] [4] = 1'b1;
  assign \A[9][225] [3] = 1'b1;
  assign \A[9][225] [2] = 1'b1;
  assign \A[9][225] [1] = 1'b1;
  assign \A[9][225] [0] = 1'b1;
  assign \A[9][226] [4] = 1'b1;
  assign \A[9][226] [3] = 1'b1;
  assign \A[9][226] [2] = 1'b1;
  assign \A[9][226] [0] = 1'b1;
  assign \A[9][227] [4] = 1'b1;
  assign \A[9][227] [3] = 1'b1;
  assign \A[9][227] [2] = 1'b1;
  assign \A[9][227] [0] = 1'b1;
  assign \A[9][228] [4] = 1'b1;
  assign \A[9][228] [3] = 1'b1;
  assign \A[9][228] [2] = 1'b1;
  assign \A[9][228] [1] = 1'b1;
  assign \A[9][228] [0] = 1'b1;
  assign \A[9][229] [4] = 1'b1;
  assign \A[9][229] [3] = 1'b1;
  assign \A[9][229] [2] = 1'b1;
  assign \A[9][229] [1] = 1'b1;
  assign \A[9][229] [0] = 1'b1;
  assign \A[9][230] [4] = 1'b1;
  assign \A[9][230] [3] = 1'b1;
  assign \A[9][230] [2] = 1'b1;
  assign \A[9][230] [0] = 1'b1;
  assign \A[9][231] [4] = 1'b1;
  assign \A[9][231] [3] = 1'b1;
  assign \A[9][231] [2] = 1'b1;
  assign \A[9][231] [1] = 1'b1;
  assign \A[9][231] [0] = 1'b1;
  assign \A[9][232] [4] = 1'b1;
  assign \A[9][232] [3] = 1'b1;
  assign \A[9][232] [2] = 1'b1;
  assign \A[9][232] [1] = 1'b1;
  assign \A[9][233] [4] = 1'b1;
  assign \A[9][233] [3] = 1'b1;
  assign \A[9][233] [2] = 1'b1;
  assign \A[9][233] [1] = 1'b1;
  assign \A[9][234] [4] = 1'b1;
  assign \A[9][234] [3] = 1'b1;
  assign \A[9][234] [2] = 1'b1;
  assign \A[9][235] [4] = 1'b1;
  assign \A[9][235] [3] = 1'b1;
  assign \A[9][235] [2] = 1'b1;
  assign \A[9][235] [1] = 1'b1;
  assign \A[9][235] [0] = 1'b1;
  assign \A[9][236] [0] = 1'b1;
  assign \A[9][238] [4] = 1'b1;
  assign \A[9][238] [3] = 1'b1;
  assign \A[9][238] [2] = 1'b1;
  assign \A[9][238] [1] = 1'b1;
  assign \A[9][239] [4] = 1'b1;
  assign \A[9][239] [3] = 1'b1;
  assign \A[9][239] [2] = 1'b1;
  assign \A[9][239] [1] = 1'b1;
  assign \A[9][239] [0] = 1'b1;
  assign \A[9][240] [4] = 1'b1;
  assign \A[9][240] [3] = 1'b1;
  assign \A[9][240] [2] = 1'b1;
  assign \A[9][240] [1] = 1'b1;
  assign \A[9][240] [0] = 1'b1;
  assign \A[9][241] [4] = 1'b1;
  assign \A[9][241] [3] = 1'b1;
  assign \A[9][241] [2] = 1'b1;
  assign \A[9][241] [0] = 1'b1;
  assign \A[9][242] [1] = 1'b1;
  assign \A[9][244] [4] = 1'b1;
  assign \A[9][244] [3] = 1'b1;
  assign \A[9][244] [2] = 1'b1;
  assign \A[9][244] [1] = 1'b1;
  assign \A[9][245] [4] = 1'b1;
  assign \A[9][245] [3] = 1'b1;
  assign \A[9][245] [1] = 1'b1;
  assign \A[9][245] [0] = 1'b1;
  assign \A[9][246] [4] = 1'b1;
  assign \A[9][246] [3] = 1'b1;
  assign \A[9][246] [2] = 1'b1;
  assign \A[9][246] [1] = 1'b1;
  assign \A[9][246] [0] = 1'b1;
  assign \A[9][247] [4] = 1'b1;
  assign \A[9][247] [3] = 1'b1;
  assign \A[9][247] [2] = 1'b1;
  assign \A[9][247] [1] = 1'b1;
  assign \A[9][247] [0] = 1'b1;
  assign \A[9][248] [4] = 1'b1;
  assign \A[9][248] [3] = 1'b1;
  assign \A[9][248] [2] = 1'b1;
  assign \A[9][248] [1] = 1'b1;
  assign \A[9][248] [0] = 1'b1;
  assign \A[9][250] [4] = 1'b1;
  assign \A[9][250] [3] = 1'b1;
  assign \A[9][250] [2] = 1'b1;
  assign \A[9][250] [1] = 1'b1;
  assign \A[9][251] [4] = 1'b1;
  assign \A[9][251] [3] = 1'b1;
  assign \A[9][251] [2] = 1'b1;
  assign \A[9][251] [1] = 1'b1;
  assign \A[9][251] [0] = 1'b1;
  assign \A[9][252] [4] = 1'b1;
  assign \A[9][252] [3] = 1'b1;
  assign \A[9][252] [2] = 1'b1;
  assign \A[9][252] [1] = 1'b1;
  assign \A[9][252] [0] = 1'b1;
  assign \A[9][253] [4] = 1'b1;
  assign \A[9][253] [3] = 1'b1;
  assign \A[9][253] [1] = 1'b1;
  assign \A[9][253] [0] = 1'b1;
  assign \A[9][254] [4] = 1'b1;
  assign \A[9][254] [3] = 1'b1;
  assign \A[9][254] [2] = 1'b1;
  assign \A[9][254] [0] = 1'b1;
  assign \A[9][255] [1] = 1'b1;
  assign \A[10][0] [4] = 1'b1;
  assign \A[10][0] [3] = 1'b1;
  assign \A[10][0] [2] = 1'b1;
  assign \A[10][0] [1] = 1'b1;
  assign \A[10][1] [0] = 1'b1;
  assign \A[10][2] [4] = 1'b1;
  assign \A[10][2] [3] = 1'b1;
  assign \A[10][2] [2] = 1'b1;
  assign \A[10][2] [1] = 1'b1;
  assign \A[10][2] [0] = 1'b1;
  assign \A[10][3] [4] = 1'b1;
  assign \A[10][3] [3] = 1'b1;
  assign \A[10][3] [2] = 1'b1;
  assign \A[10][3] [1] = 1'b1;
  assign \A[10][3] [0] = 1'b1;
  assign \A[10][4] [4] = 1'b1;
  assign \A[10][4] [3] = 1'b1;
  assign \A[10][4] [2] = 1'b1;
  assign \A[10][4] [1] = 1'b1;
  assign \A[10][5] [4] = 1'b1;
  assign \A[10][5] [3] = 1'b1;
  assign \A[10][5] [2] = 1'b1;
  assign \A[10][5] [0] = 1'b1;
  assign \A[10][6] [4] = 1'b1;
  assign \A[10][6] [3] = 1'b1;
  assign \A[10][6] [2] = 1'b1;
  assign \A[10][6] [1] = 1'b1;
  assign \A[10][6] [0] = 1'b1;
  assign \A[10][7] [0] = 1'b1;
  assign \A[10][8] [4] = 1'b1;
  assign \A[10][8] [3] = 1'b1;
  assign \A[10][8] [2] = 1'b1;
  assign \A[10][8] [1] = 1'b1;
  assign \A[10][10] [4] = 1'b1;
  assign \A[10][10] [3] = 1'b1;
  assign \A[10][10] [2] = 1'b1;
  assign \A[10][10] [1] = 1'b1;
  assign \A[10][10] [0] = 1'b1;
  assign \A[10][12] [4] = 1'b1;
  assign \A[10][12] [3] = 1'b1;
  assign \A[10][12] [2] = 1'b1;
  assign \A[10][12] [1] = 1'b1;
  assign \A[10][12] [0] = 1'b1;
  assign \A[10][15] [0] = 1'b1;
  assign \A[10][16] [4] = 1'b1;
  assign \A[10][16] [3] = 1'b1;
  assign \A[10][16] [2] = 1'b1;
  assign \A[10][16] [1] = 1'b1;
  assign \A[10][16] [0] = 1'b1;
  assign \A[10][17] [0] = 1'b1;
  assign \A[10][18] [4] = 1'b1;
  assign \A[10][18] [3] = 1'b1;
  assign \A[10][18] [2] = 1'b1;
  assign \A[10][18] [1] = 1'b1;
  assign \A[10][19] [4] = 1'b1;
  assign \A[10][19] [3] = 1'b1;
  assign \A[10][19] [2] = 1'b1;
  assign \A[10][19] [1] = 1'b1;
  assign \A[10][19] [0] = 1'b1;
  assign \A[10][20] [1] = 1'b1;
  assign \A[10][21] [0] = 1'b1;
  assign \A[10][23] [4] = 1'b1;
  assign \A[10][23] [3] = 1'b1;
  assign \A[10][23] [2] = 1'b1;
  assign \A[10][23] [1] = 1'b1;
  assign \A[10][23] [0] = 1'b1;
  assign \A[10][24] [4] = 1'b1;
  assign \A[10][24] [3] = 1'b1;
  assign \A[10][24] [2] = 1'b1;
  assign \A[10][24] [1] = 1'b1;
  assign \A[10][24] [0] = 1'b1;
  assign \A[10][25] [4] = 1'b1;
  assign \A[10][25] [3] = 1'b1;
  assign \A[10][25] [2] = 1'b1;
  assign \A[10][25] [1] = 1'b1;
  assign \A[10][27] [4] = 1'b1;
  assign \A[10][27] [3] = 1'b1;
  assign \A[10][27] [2] = 1'b1;
  assign \A[10][27] [1] = 1'b1;
  assign \A[10][27] [0] = 1'b1;
  assign \A[10][28] [0] = 1'b1;
  assign \A[10][29] [4] = 1'b1;
  assign \A[10][29] [3] = 1'b1;
  assign \A[10][29] [2] = 1'b1;
  assign \A[10][29] [1] = 1'b1;
  assign \A[10][29] [0] = 1'b1;
  assign \A[10][30] [0] = 1'b1;
  assign \A[10][32] [4] = 1'b1;
  assign \A[10][32] [3] = 1'b1;
  assign \A[10][32] [2] = 1'b1;
  assign \A[10][32] [1] = 1'b1;
  assign \A[10][33] [0] = 1'b1;
  assign \A[10][35] [4] = 1'b1;
  assign \A[10][35] [3] = 1'b1;
  assign \A[10][35] [2] = 1'b1;
  assign \A[10][35] [1] = 1'b1;
  assign \A[10][37] [1] = 1'b1;
  assign \A[10][38] [4] = 1'b1;
  assign \A[10][38] [3] = 1'b1;
  assign \A[10][38] [2] = 1'b1;
  assign \A[10][38] [1] = 1'b1;
  assign \A[10][39] [4] = 1'b1;
  assign \A[10][39] [3] = 1'b1;
  assign \A[10][39] [2] = 1'b1;
  assign \A[10][39] [1] = 1'b1;
  assign \A[10][40] [0] = 1'b1;
  assign \A[10][41] [0] = 1'b1;
  assign \A[10][42] [4] = 1'b1;
  assign \A[10][42] [3] = 1'b1;
  assign \A[10][42] [2] = 1'b1;
  assign \A[10][42] [1] = 1'b1;
  assign \A[10][43] [4] = 1'b1;
  assign \A[10][43] [3] = 1'b1;
  assign \A[10][43] [2] = 1'b1;
  assign \A[10][43] [1] = 1'b1;
  assign \A[10][43] [0] = 1'b1;
  assign \A[10][44] [4] = 1'b1;
  assign \A[10][44] [3] = 1'b1;
  assign \A[10][44] [2] = 1'b1;
  assign \A[10][44] [1] = 1'b1;
  assign \A[10][44] [0] = 1'b1;
  assign \A[10][46] [4] = 1'b1;
  assign \A[10][46] [3] = 1'b1;
  assign \A[10][46] [2] = 1'b1;
  assign \A[10][46] [1] = 1'b1;
  assign \A[10][46] [0] = 1'b1;
  assign \A[10][48] [4] = 1'b1;
  assign \A[10][48] [3] = 1'b1;
  assign \A[10][48] [2] = 1'b1;
  assign \A[10][48] [1] = 1'b1;
  assign \A[10][48] [0] = 1'b1;
  assign \A[10][49] [4] = 1'b1;
  assign \A[10][49] [3] = 1'b1;
  assign \A[10][49] [2] = 1'b1;
  assign \A[10][49] [1] = 1'b1;
  assign \A[10][49] [0] = 1'b1;
  assign \A[10][51] [1] = 1'b1;
  assign \A[10][52] [1] = 1'b1;
  assign \A[10][53] [1] = 1'b1;
  assign \A[10][55] [4] = 1'b1;
  assign \A[10][55] [3] = 1'b1;
  assign \A[10][55] [2] = 1'b1;
  assign \A[10][55] [1] = 1'b1;
  assign \A[10][56] [0] = 1'b1;
  assign \A[10][57] [4] = 1'b1;
  assign \A[10][57] [3] = 1'b1;
  assign \A[10][57] [2] = 1'b1;
  assign \A[10][57] [0] = 1'b1;
  assign \A[10][60] [0] = 1'b1;
  assign \A[10][61] [4] = 1'b1;
  assign \A[10][61] [3] = 1'b1;
  assign \A[10][61] [2] = 1'b1;
  assign \A[10][61] [1] = 1'b1;
  assign \A[10][61] [0] = 1'b1;
  assign \A[10][63] [4] = 1'b1;
  assign \A[10][63] [3] = 1'b1;
  assign \A[10][63] [2] = 1'b1;
  assign \A[10][63] [1] = 1'b1;
  assign \A[10][65] [0] = 1'b1;
  assign \A[10][66] [0] = 1'b1;
  assign \A[10][67] [4] = 1'b1;
  assign \A[10][67] [3] = 1'b1;
  assign \A[10][67] [2] = 1'b1;
  assign \A[10][67] [1] = 1'b1;
  assign \A[10][67] [0] = 1'b1;
  assign \A[10][70] [0] = 1'b1;
  assign \A[10][72] [4] = 1'b1;
  assign \A[10][72] [3] = 1'b1;
  assign \A[10][72] [2] = 1'b1;
  assign \A[10][72] [1] = 1'b1;
  assign \A[10][72] [0] = 1'b1;
  assign \A[10][73] [4] = 1'b1;
  assign \A[10][73] [3] = 1'b1;
  assign \A[10][73] [2] = 1'b1;
  assign \A[10][73] [1] = 1'b1;
  assign \A[10][75] [1] = 1'b1;
  assign \A[10][76] [4] = 1'b1;
  assign \A[10][76] [3] = 1'b1;
  assign \A[10][76] [2] = 1'b1;
  assign \A[10][76] [1] = 1'b1;
  assign \A[10][76] [0] = 1'b1;
  assign \A[10][78] [1] = 1'b1;
  assign \A[10][79] [0] = 1'b1;
  assign \A[10][80] [0] = 1'b1;
  assign \A[10][82] [0] = 1'b1;
  assign \A[10][83] [4] = 1'b1;
  assign \A[10][83] [3] = 1'b1;
  assign \A[10][83] [2] = 1'b1;
  assign \A[10][83] [1] = 1'b1;
  assign \A[10][83] [0] = 1'b1;
  assign \A[10][84] [4] = 1'b1;
  assign \A[10][84] [3] = 1'b1;
  assign \A[10][84] [2] = 1'b1;
  assign \A[10][84] [1] = 1'b1;
  assign \A[10][84] [0] = 1'b1;
  assign \A[10][85] [4] = 1'b1;
  assign \A[10][85] [3] = 1'b1;
  assign \A[10][85] [2] = 1'b1;
  assign \A[10][85] [1] = 1'b1;
  assign \A[10][86] [0] = 1'b1;
  assign \A[10][91] [0] = 1'b1;
  assign \A[10][92] [4] = 1'b1;
  assign \A[10][92] [3] = 1'b1;
  assign \A[10][92] [2] = 1'b1;
  assign \A[10][92] [1] = 1'b1;
  assign \A[10][92] [0] = 1'b1;
  assign \A[10][94] [0] = 1'b1;
  assign \A[10][95] [0] = 1'b1;
  assign \A[10][96] [1] = 1'b1;
  assign \A[10][97] [4] = 1'b1;
  assign \A[10][97] [3] = 1'b1;
  assign \A[10][97] [2] = 1'b1;
  assign \A[10][97] [1] = 1'b1;
  assign \A[10][97] [0] = 1'b1;
  assign \A[10][98] [0] = 1'b1;
  assign \A[10][101] [1] = 1'b1;
  assign \A[10][101] [0] = 1'b1;
  assign \A[10][102] [1] = 1'b1;
  assign \A[10][102] [0] = 1'b1;
  assign \A[10][103] [4] = 1'b1;
  assign \A[10][103] [3] = 1'b1;
  assign \A[10][103] [2] = 1'b1;
  assign \A[10][103] [1] = 1'b1;
  assign \A[10][103] [0] = 1'b1;
  assign \A[10][106] [4] = 1'b1;
  assign \A[10][106] [3] = 1'b1;
  assign \A[10][106] [2] = 1'b1;
  assign \A[10][106] [1] = 1'b1;
  assign \A[10][107] [4] = 1'b1;
  assign \A[10][107] [3] = 1'b1;
  assign \A[10][107] [2] = 1'b1;
  assign \A[10][107] [0] = 1'b1;
  assign \A[10][108] [4] = 1'b1;
  assign \A[10][108] [3] = 1'b1;
  assign \A[10][108] [2] = 1'b1;
  assign \A[10][108] [1] = 1'b1;
  assign \A[10][108] [0] = 1'b1;
  assign \A[10][109] [4] = 1'b1;
  assign \A[10][109] [3] = 1'b1;
  assign \A[10][109] [2] = 1'b1;
  assign \A[10][109] [1] = 1'b1;
  assign \A[10][109] [0] = 1'b1;
  assign \A[10][110] [4] = 1'b1;
  assign \A[10][110] [3] = 1'b1;
  assign \A[10][110] [2] = 1'b1;
  assign \A[10][110] [0] = 1'b1;
  assign \A[10][112] [4] = 1'b1;
  assign \A[10][112] [3] = 1'b1;
  assign \A[10][112] [2] = 1'b1;
  assign \A[10][112] [1] = 1'b1;
  assign \A[10][114] [0] = 1'b1;
  assign \A[10][115] [4] = 1'b1;
  assign \A[10][115] [3] = 1'b1;
  assign \A[10][115] [2] = 1'b1;
  assign \A[10][115] [0] = 1'b1;
  assign \A[10][116] [0] = 1'b1;
  assign \A[10][117] [4] = 1'b1;
  assign \A[10][117] [3] = 1'b1;
  assign \A[10][117] [2] = 1'b1;
  assign \A[10][117] [1] = 1'b1;
  assign \A[10][117] [0] = 1'b1;
  assign \A[10][118] [4] = 1'b1;
  assign \A[10][118] [3] = 1'b1;
  assign \A[10][118] [2] = 1'b1;
  assign \A[10][118] [1] = 1'b1;
  assign \A[10][118] [0] = 1'b1;
  assign \A[10][119] [4] = 1'b1;
  assign \A[10][119] [3] = 1'b1;
  assign \A[10][119] [2] = 1'b1;
  assign \A[10][119] [1] = 1'b1;
  assign \A[10][119] [0] = 1'b1;
  assign \A[10][120] [0] = 1'b1;
  assign \A[10][121] [4] = 1'b1;
  assign \A[10][121] [3] = 1'b1;
  assign \A[10][121] [2] = 1'b1;
  assign \A[10][121] [1] = 1'b1;
  assign \A[10][121] [0] = 1'b1;
  assign \A[10][122] [4] = 1'b1;
  assign \A[10][122] [3] = 1'b1;
  assign \A[10][122] [2] = 1'b1;
  assign \A[10][122] [0] = 1'b1;
  assign \A[10][123] [4] = 1'b1;
  assign \A[10][123] [3] = 1'b1;
  assign \A[10][123] [2] = 1'b1;
  assign \A[10][123] [1] = 1'b1;
  assign \A[10][123] [0] = 1'b1;
  assign \A[10][124] [1] = 1'b1;
  assign \A[10][125] [0] = 1'b1;
  assign \A[10][126] [0] = 1'b1;
  assign \A[10][127] [0] = 1'b1;
  assign \A[10][128] [0] = 1'b1;
  assign \A[10][131] [0] = 1'b1;
  assign \A[10][133] [0] = 1'b1;
  assign \A[10][134] [0] = 1'b1;
  assign \A[10][135] [4] = 1'b1;
  assign \A[10][135] [3] = 1'b1;
  assign \A[10][135] [2] = 1'b1;
  assign \A[10][135] [1] = 1'b1;
  assign \A[10][135] [0] = 1'b1;
  assign \A[10][136] [4] = 1'b1;
  assign \A[10][136] [3] = 1'b1;
  assign \A[10][136] [2] = 1'b1;
  assign \A[10][136] [1] = 1'b1;
  assign \A[10][139] [1] = 1'b1;
  assign \A[10][140] [4] = 1'b1;
  assign \A[10][140] [3] = 1'b1;
  assign \A[10][140] [2] = 1'b1;
  assign \A[10][140] [1] = 1'b1;
  assign \A[10][142] [0] = 1'b1;
  assign \A[10][144] [4] = 1'b1;
  assign \A[10][144] [3] = 1'b1;
  assign \A[10][144] [2] = 1'b1;
  assign \A[10][144] [1] = 1'b1;
  assign \A[10][144] [0] = 1'b1;
  assign \A[10][145] [4] = 1'b1;
  assign \A[10][145] [3] = 1'b1;
  assign \A[10][145] [2] = 1'b1;
  assign \A[10][145] [0] = 1'b1;
  assign \A[10][146] [4] = 1'b1;
  assign \A[10][146] [3] = 1'b1;
  assign \A[10][146] [2] = 1'b1;
  assign \A[10][146] [1] = 1'b1;
  assign \A[10][146] [0] = 1'b1;
  assign \A[10][147] [4] = 1'b1;
  assign \A[10][147] [3] = 1'b1;
  assign \A[10][147] [2] = 1'b1;
  assign \A[10][147] [1] = 1'b1;
  assign \A[10][147] [0] = 1'b1;
  assign \A[10][149] [4] = 1'b1;
  assign \A[10][149] [3] = 1'b1;
  assign \A[10][149] [2] = 1'b1;
  assign \A[10][149] [1] = 1'b1;
  assign \A[10][149] [0] = 1'b1;
  assign \A[10][150] [4] = 1'b1;
  assign \A[10][150] [3] = 1'b1;
  assign \A[10][150] [2] = 1'b1;
  assign \A[10][150] [1] = 1'b1;
  assign \A[10][150] [0] = 1'b1;
  assign \A[10][151] [0] = 1'b1;
  assign \A[10][152] [1] = 1'b1;
  assign \A[10][155] [0] = 1'b1;
  assign \A[10][157] [1] = 1'b1;
  assign \A[10][159] [1] = 1'b1;
  assign \A[10][162] [1] = 1'b1;
  assign \A[10][163] [1] = 1'b1;
  assign \A[10][163] [0] = 1'b1;
  assign \A[10][165] [4] = 1'b1;
  assign \A[10][165] [3] = 1'b1;
  assign \A[10][165] [2] = 1'b1;
  assign \A[10][165] [1] = 1'b1;
  assign \A[10][165] [0] = 1'b1;
  assign \A[10][166] [1] = 1'b1;
  assign \A[10][167] [0] = 1'b1;
  assign \A[10][168] [4] = 1'b1;
  assign \A[10][168] [3] = 1'b1;
  assign \A[10][168] [2] = 1'b1;
  assign \A[10][168] [0] = 1'b1;
  assign \A[10][170] [4] = 1'b1;
  assign \A[10][170] [3] = 1'b1;
  assign \A[10][170] [2] = 1'b1;
  assign \A[10][170] [1] = 1'b1;
  assign \A[10][170] [0] = 1'b1;
  assign \A[10][171] [0] = 1'b1;
  assign \A[10][172] [4] = 1'b1;
  assign \A[10][172] [3] = 1'b1;
  assign \A[10][172] [2] = 1'b1;
  assign \A[10][172] [1] = 1'b1;
  assign \A[10][175] [4] = 1'b1;
  assign \A[10][175] [3] = 1'b1;
  assign \A[10][175] [2] = 1'b1;
  assign \A[10][175] [1] = 1'b1;
  assign \A[10][175] [0] = 1'b1;
  assign \A[10][177] [0] = 1'b1;
  assign \A[10][178] [4] = 1'b1;
  assign \A[10][178] [3] = 1'b1;
  assign \A[10][178] [2] = 1'b1;
  assign \A[10][178] [1] = 1'b1;
  assign \A[10][178] [0] = 1'b1;
  assign \A[10][179] [1] = 1'b1;
  assign \A[10][180] [4] = 1'b1;
  assign \A[10][180] [3] = 1'b1;
  assign \A[10][180] [2] = 1'b1;
  assign \A[10][180] [1] = 1'b1;
  assign \A[10][180] [0] = 1'b1;
  assign \A[10][181] [4] = 1'b1;
  assign \A[10][181] [3] = 1'b1;
  assign \A[10][181] [2] = 1'b1;
  assign \A[10][181] [1] = 1'b1;
  assign \A[10][182] [4] = 1'b1;
  assign \A[10][182] [3] = 1'b1;
  assign \A[10][182] [2] = 1'b1;
  assign \A[10][182] [1] = 1'b1;
  assign \A[10][182] [0] = 1'b1;
  assign \A[10][183] [4] = 1'b1;
  assign \A[10][183] [3] = 1'b1;
  assign \A[10][183] [2] = 1'b1;
  assign \A[10][183] [1] = 1'b1;
  assign \A[10][183] [0] = 1'b1;
  assign \A[10][186] [4] = 1'b1;
  assign \A[10][186] [3] = 1'b1;
  assign \A[10][186] [2] = 1'b1;
  assign \A[10][186] [0] = 1'b1;
  assign \A[10][187] [4] = 1'b1;
  assign \A[10][187] [3] = 1'b1;
  assign \A[10][187] [2] = 1'b1;
  assign \A[10][187] [1] = 1'b1;
  assign \A[10][188] [0] = 1'b1;
  assign \A[10][189] [0] = 1'b1;
  assign \A[10][190] [0] = 1'b1;
  assign \A[10][193] [0] = 1'b1;
  assign \A[10][194] [4] = 1'b1;
  assign \A[10][194] [3] = 1'b1;
  assign \A[10][194] [2] = 1'b1;
  assign \A[10][194] [1] = 1'b1;
  assign \A[10][194] [0] = 1'b1;
  assign \A[10][195] [0] = 1'b1;
  assign \A[10][196] [4] = 1'b1;
  assign \A[10][196] [3] = 1'b1;
  assign \A[10][196] [2] = 1'b1;
  assign \A[10][196] [1] = 1'b1;
  assign \A[10][197] [4] = 1'b1;
  assign \A[10][197] [3] = 1'b1;
  assign \A[10][197] [2] = 1'b1;
  assign \A[10][197] [1] = 1'b1;
  assign \A[10][198] [0] = 1'b1;
  assign \A[10][200] [4] = 1'b1;
  assign \A[10][200] [3] = 1'b1;
  assign \A[10][200] [2] = 1'b1;
  assign \A[10][200] [1] = 1'b1;
  assign \A[10][200] [0] = 1'b1;
  assign \A[10][202] [4] = 1'b1;
  assign \A[10][202] [3] = 1'b1;
  assign \A[10][202] [2] = 1'b1;
  assign \A[10][202] [1] = 1'b1;
  assign \A[10][202] [0] = 1'b1;
  assign \A[10][203] [0] = 1'b1;
  assign \A[10][204] [0] = 1'b1;
  assign \A[10][206] [0] = 1'b1;
  assign \A[10][207] [0] = 1'b1;
  assign \A[10][208] [0] = 1'b1;
  assign \A[10][209] [4] = 1'b1;
  assign \A[10][209] [3] = 1'b1;
  assign \A[10][209] [2] = 1'b1;
  assign \A[10][209] [1] = 1'b1;
  assign \A[10][210] [4] = 1'b1;
  assign \A[10][210] [3] = 1'b1;
  assign \A[10][210] [2] = 1'b1;
  assign \A[10][210] [1] = 1'b1;
  assign \A[10][210] [0] = 1'b1;
  assign \A[10][211] [4] = 1'b1;
  assign \A[10][211] [3] = 1'b1;
  assign \A[10][211] [2] = 1'b1;
  assign \A[10][211] [1] = 1'b1;
  assign \A[10][211] [0] = 1'b1;
  assign \A[10][212] [1] = 1'b1;
  assign \A[10][213] [4] = 1'b1;
  assign \A[10][213] [3] = 1'b1;
  assign \A[10][213] [2] = 1'b1;
  assign \A[10][213] [1] = 1'b1;
  assign \A[10][213] [0] = 1'b1;
  assign \A[10][215] [1] = 1'b1;
  assign \A[10][216] [4] = 1'b1;
  assign \A[10][216] [3] = 1'b1;
  assign \A[10][216] [2] = 1'b1;
  assign \A[10][216] [1] = 1'b1;
  assign \A[10][219] [1] = 1'b1;
  assign \A[10][220] [1] = 1'b1;
  assign \A[10][220] [0] = 1'b1;
  assign \A[10][221] [4] = 1'b1;
  assign \A[10][221] [3] = 1'b1;
  assign \A[10][221] [2] = 1'b1;
  assign \A[10][221] [1] = 1'b1;
  assign \A[10][221] [0] = 1'b1;
  assign \A[10][223] [1] = 1'b1;
  assign \A[10][224] [0] = 1'b1;
  assign \A[10][226] [1] = 1'b1;
  assign \A[10][227] [4] = 1'b1;
  assign \A[10][227] [3] = 1'b1;
  assign \A[10][227] [2] = 1'b1;
  assign \A[10][227] [1] = 1'b1;
  assign \A[10][227] [0] = 1'b1;
  assign \A[10][228] [1] = 1'b1;
  assign \A[10][229] [4] = 1'b1;
  assign \A[10][229] [3] = 1'b1;
  assign \A[10][229] [2] = 1'b1;
  assign \A[10][229] [1] = 1'b1;
  assign \A[10][229] [0] = 1'b1;
  assign \A[10][230] [0] = 1'b1;
  assign \A[10][231] [4] = 1'b1;
  assign \A[10][231] [3] = 1'b1;
  assign \A[10][231] [2] = 1'b1;
  assign \A[10][231] [1] = 1'b1;
  assign \A[10][231] [0] = 1'b1;
  assign \A[10][232] [4] = 1'b1;
  assign \A[10][232] [3] = 1'b1;
  assign \A[10][232] [2] = 1'b1;
  assign \A[10][232] [1] = 1'b1;
  assign \A[10][233] [4] = 1'b1;
  assign \A[10][233] [3] = 1'b1;
  assign \A[10][233] [2] = 1'b1;
  assign \A[10][233] [1] = 1'b1;
  assign \A[10][236] [4] = 1'b1;
  assign \A[10][236] [3] = 1'b1;
  assign \A[10][236] [2] = 1'b1;
  assign \A[10][236] [0] = 1'b1;
  assign \A[10][239] [4] = 1'b1;
  assign \A[10][239] [3] = 1'b1;
  assign \A[10][239] [2] = 1'b1;
  assign \A[10][239] [1] = 1'b1;
  assign \A[10][239] [0] = 1'b1;
  assign \A[10][240] [4] = 1'b1;
  assign \A[10][240] [3] = 1'b1;
  assign \A[10][240] [2] = 1'b1;
  assign \A[10][240] [1] = 1'b1;
  assign \A[10][240] [0] = 1'b1;
  assign \A[10][241] [0] = 1'b1;
  assign \A[10][242] [0] = 1'b1;
  assign \A[10][243] [0] = 1'b1;
  assign \A[10][244] [4] = 1'b1;
  assign \A[10][244] [3] = 1'b1;
  assign \A[10][244] [2] = 1'b1;
  assign \A[10][244] [1] = 1'b1;
  assign \A[10][244] [0] = 1'b1;
  assign \A[10][246] [4] = 1'b1;
  assign \A[10][246] [3] = 1'b1;
  assign \A[10][246] [2] = 1'b1;
  assign \A[10][246] [1] = 1'b1;
  assign \A[10][246] [0] = 1'b1;
  assign \A[10][247] [0] = 1'b1;
  assign \A[10][248] [4] = 1'b1;
  assign \A[10][248] [3] = 1'b1;
  assign \A[10][248] [2] = 1'b1;
  assign \A[10][248] [1] = 1'b1;
  assign \A[10][250] [4] = 1'b1;
  assign \A[10][250] [3] = 1'b1;
  assign \A[10][250] [2] = 1'b1;
  assign \A[10][250] [1] = 1'b1;
  assign \A[10][250] [0] = 1'b1;
  assign \A[10][251] [4] = 1'b1;
  assign \A[10][251] [3] = 1'b1;
  assign \A[10][251] [2] = 1'b1;
  assign \A[10][251] [1] = 1'b1;
  assign \A[10][251] [0] = 1'b1;
  assign \A[10][252] [0] = 1'b1;
  assign \A[10][253] [4] = 1'b1;
  assign \A[10][253] [3] = 1'b1;
  assign \A[10][253] [2] = 1'b1;
  assign \A[10][253] [1] = 1'b1;
  assign \A[10][253] [0] = 1'b1;
  assign \A[11][0] [2] = 1'b1;
  assign \A[11][1] [4] = 1'b1;
  assign \A[11][1] [3] = 1'b1;
  assign \A[11][1] [2] = 1'b1;
  assign \A[11][1] [1] = 1'b1;
  assign \A[11][2] [4] = 1'b1;
  assign \A[11][2] [3] = 1'b1;
  assign \A[11][2] [2] = 1'b1;
  assign \A[11][2] [1] = 1'b1;
  assign \A[11][2] [0] = 1'b1;
  assign \A[11][4] [4] = 1'b1;
  assign \A[11][4] [3] = 1'b1;
  assign \A[11][4] [2] = 1'b1;
  assign \A[11][4] [1] = 1'b1;
  assign \A[11][4] [0] = 1'b1;
  assign \A[11][5] [4] = 1'b1;
  assign \A[11][5] [3] = 1'b1;
  assign \A[11][5] [2] = 1'b1;
  assign \A[11][5] [0] = 1'b1;
  assign \A[11][7] [0] = 1'b1;
  assign \A[11][8] [4] = 1'b1;
  assign \A[11][8] [3] = 1'b1;
  assign \A[11][8] [1] = 1'b1;
  assign \A[11][8] [0] = 1'b1;
  assign \A[11][9] [4] = 1'b1;
  assign \A[11][9] [3] = 1'b1;
  assign \A[11][9] [2] = 1'b1;
  assign \A[11][9] [1] = 1'b1;
  assign \A[11][11] [4] = 1'b1;
  assign \A[11][11] [3] = 1'b1;
  assign \A[11][11] [2] = 1'b1;
  assign \A[11][11] [0] = 1'b1;
  assign \A[11][12] [4] = 1'b1;
  assign \A[11][12] [3] = 1'b1;
  assign \A[11][12] [2] = 1'b1;
  assign \A[11][12] [1] = 1'b1;
  assign \A[11][13] [0] = 1'b1;
  assign \A[11][14] [4] = 1'b1;
  assign \A[11][14] [3] = 1'b1;
  assign \A[11][14] [2] = 1'b1;
  assign \A[11][14] [1] = 1'b1;
  assign \A[11][15] [0] = 1'b1;
  assign \A[11][16] [4] = 1'b1;
  assign \A[11][16] [3] = 1'b1;
  assign \A[11][16] [2] = 1'b1;
  assign \A[11][16] [0] = 1'b1;
  assign \A[11][18] [4] = 1'b1;
  assign \A[11][18] [3] = 1'b1;
  assign \A[11][18] [2] = 1'b1;
  assign \A[11][18] [1] = 1'b1;
  assign \A[11][18] [0] = 1'b1;
  assign \A[11][20] [4] = 1'b1;
  assign \A[11][20] [3] = 1'b1;
  assign \A[11][20] [2] = 1'b1;
  assign \A[11][20] [1] = 1'b1;
  assign \A[11][20] [0] = 1'b1;
  assign \A[11][21] [4] = 1'b1;
  assign \A[11][21] [3] = 1'b1;
  assign \A[11][21] [2] = 1'b1;
  assign \A[11][21] [1] = 1'b1;
  assign \A[11][21] [0] = 1'b1;
  assign \A[11][22] [4] = 1'b1;
  assign \A[11][22] [3] = 1'b1;
  assign \A[11][22] [1] = 1'b1;
  assign \A[11][22] [0] = 1'b1;
  assign \A[11][23] [4] = 1'b1;
  assign \A[11][23] [3] = 1'b1;
  assign \A[11][23] [2] = 1'b1;
  assign \A[11][23] [1] = 1'b1;
  assign \A[11][23] [0] = 1'b1;
  assign \A[11][24] [4] = 1'b1;
  assign \A[11][24] [3] = 1'b1;
  assign \A[11][24] [2] = 1'b1;
  assign \A[11][24] [0] = 1'b1;
  assign \A[11][25] [4] = 1'b1;
  assign \A[11][25] [3] = 1'b1;
  assign \A[11][25] [2] = 1'b1;
  assign \A[11][25] [1] = 1'b1;
  assign \A[11][25] [0] = 1'b1;
  assign \A[11][27] [1] = 1'b1;
  assign \A[11][29] [4] = 1'b1;
  assign \A[11][29] [3] = 1'b1;
  assign \A[11][29] [2] = 1'b1;
  assign \A[11][29] [1] = 1'b1;
  assign \A[11][29] [0] = 1'b1;
  assign \A[11][30] [1] = 1'b1;
  assign \A[11][31] [4] = 1'b1;
  assign \A[11][31] [3] = 1'b1;
  assign \A[11][31] [2] = 1'b1;
  assign \A[11][31] [1] = 1'b1;
  assign \A[11][31] [0] = 1'b1;
  assign \A[11][32] [4] = 1'b1;
  assign \A[11][32] [3] = 1'b1;
  assign \A[11][32] [2] = 1'b1;
  assign \A[11][32] [1] = 1'b1;
  assign \A[11][33] [4] = 1'b1;
  assign \A[11][33] [3] = 1'b1;
  assign \A[11][33] [2] = 1'b1;
  assign \A[11][33] [1] = 1'b1;
  assign \A[11][33] [0] = 1'b1;
  assign \A[11][34] [0] = 1'b1;
  assign \A[11][35] [4] = 1'b1;
  assign \A[11][35] [3] = 1'b1;
  assign \A[11][35] [2] = 1'b1;
  assign \A[11][35] [1] = 1'b1;
  assign \A[11][35] [0] = 1'b1;
  assign \A[11][36] [4] = 1'b1;
  assign \A[11][36] [3] = 1'b1;
  assign \A[11][36] [2] = 1'b1;
  assign \A[11][36] [1] = 1'b1;
  assign \A[11][36] [0] = 1'b1;
  assign \A[11][37] [1] = 1'b1;
  assign \A[11][40] [4] = 1'b1;
  assign \A[11][40] [3] = 1'b1;
  assign \A[11][40] [2] = 1'b1;
  assign \A[11][40] [1] = 1'b1;
  assign \A[11][41] [4] = 1'b1;
  assign \A[11][41] [3] = 1'b1;
  assign \A[11][41] [2] = 1'b1;
  assign \A[11][41] [1] = 1'b1;
  assign \A[11][44] [1] = 1'b1;
  assign \A[11][45] [0] = 1'b1;
  assign \A[11][46] [4] = 1'b1;
  assign \A[11][46] [3] = 1'b1;
  assign \A[11][46] [2] = 1'b1;
  assign \A[11][46] [0] = 1'b1;
  assign \A[11][49] [4] = 1'b1;
  assign \A[11][49] [3] = 1'b1;
  assign \A[11][49] [2] = 1'b1;
  assign \A[11][49] [1] = 1'b1;
  assign \A[11][49] [0] = 1'b1;
  assign \A[11][50] [4] = 1'b1;
  assign \A[11][50] [3] = 1'b1;
  assign \A[11][50] [2] = 1'b1;
  assign \A[11][50] [0] = 1'b1;
  assign \A[11][52] [0] = 1'b1;
  assign \A[11][55] [4] = 1'b1;
  assign \A[11][55] [3] = 1'b1;
  assign \A[11][55] [2] = 1'b1;
  assign \A[11][55] [1] = 1'b1;
  assign \A[11][56] [1] = 1'b1;
  assign \A[11][57] [0] = 1'b1;
  assign \A[11][58] [0] = 1'b1;
  assign \A[11][59] [4] = 1'b1;
  assign \A[11][59] [3] = 1'b1;
  assign \A[11][59] [2] = 1'b1;
  assign \A[11][59] [1] = 1'b1;
  assign \A[11][59] [0] = 1'b1;
  assign \A[11][60] [4] = 1'b1;
  assign \A[11][60] [3] = 1'b1;
  assign \A[11][60] [1] = 1'b1;
  assign \A[11][60] [0] = 1'b1;
  assign \A[11][61] [4] = 1'b1;
  assign \A[11][61] [3] = 1'b1;
  assign \A[11][61] [2] = 1'b1;
  assign \A[11][61] [1] = 1'b1;
  assign \A[11][61] [0] = 1'b1;
  assign \A[11][62] [4] = 1'b1;
  assign \A[11][62] [3] = 1'b1;
  assign \A[11][62] [2] = 1'b1;
  assign \A[11][62] [1] = 1'b1;
  assign \A[11][63] [4] = 1'b1;
  assign \A[11][63] [3] = 1'b1;
  assign \A[11][63] [1] = 1'b1;
  assign \A[11][63] [0] = 1'b1;
  assign \A[11][65] [4] = 1'b1;
  assign \A[11][65] [3] = 1'b1;
  assign \A[11][65] [2] = 1'b1;
  assign \A[11][65] [1] = 1'b1;
  assign \A[11][66] [4] = 1'b1;
  assign \A[11][66] [3] = 1'b1;
  assign \A[11][66] [2] = 1'b1;
  assign \A[11][66] [1] = 1'b1;
  assign \A[11][66] [0] = 1'b1;
  assign \A[11][68] [1] = 1'b1;
  assign \A[11][69] [1] = 1'b1;
  assign \A[11][70] [0] = 1'b1;
  assign \A[11][71] [4] = 1'b1;
  assign \A[11][71] [3] = 1'b1;
  assign \A[11][71] [2] = 1'b1;
  assign \A[11][71] [0] = 1'b1;
  assign \A[11][73] [2] = 1'b1;
  assign \A[11][74] [4] = 1'b1;
  assign \A[11][74] [3] = 1'b1;
  assign \A[11][74] [2] = 1'b1;
  assign \A[11][74] [1] = 1'b1;
  assign \A[11][75] [4] = 1'b1;
  assign \A[11][75] [3] = 1'b1;
  assign \A[11][75] [2] = 1'b1;
  assign \A[11][75] [1] = 1'b1;
  assign \A[11][76] [4] = 1'b1;
  assign \A[11][76] [3] = 1'b1;
  assign \A[11][76] [2] = 1'b1;
  assign \A[11][76] [0] = 1'b1;
  assign \A[11][77] [4] = 1'b1;
  assign \A[11][77] [3] = 1'b1;
  assign \A[11][77] [2] = 1'b1;
  assign \A[11][77] [1] = 1'b1;
  assign \A[11][78] [4] = 1'b1;
  assign \A[11][78] [3] = 1'b1;
  assign \A[11][78] [2] = 1'b1;
  assign \A[11][78] [1] = 1'b1;
  assign \A[11][78] [0] = 1'b1;
  assign \A[11][79] [4] = 1'b1;
  assign \A[11][79] [3] = 1'b1;
  assign \A[11][79] [2] = 1'b1;
  assign \A[11][79] [1] = 1'b1;
  assign \A[11][80] [0] = 1'b1;
  assign \A[11][81] [1] = 1'b1;
  assign \A[11][83] [4] = 1'b1;
  assign \A[11][83] [3] = 1'b1;
  assign \A[11][83] [2] = 1'b1;
  assign \A[11][83] [1] = 1'b1;
  assign \A[11][83] [0] = 1'b1;
  assign \A[11][84] [0] = 1'b1;
  assign \A[11][85] [4] = 1'b1;
  assign \A[11][85] [3] = 1'b1;
  assign \A[11][85] [2] = 1'b1;
  assign \A[11][85] [1] = 1'b1;
  assign \A[11][86] [4] = 1'b1;
  assign \A[11][86] [3] = 1'b1;
  assign \A[11][86] [2] = 1'b1;
  assign \A[11][86] [1] = 1'b1;
  assign \A[11][86] [0] = 1'b1;
  assign \A[11][88] [4] = 1'b1;
  assign \A[11][88] [3] = 1'b1;
  assign \A[11][88] [2] = 1'b1;
  assign \A[11][88] [1] = 1'b1;
  assign \A[11][88] [0] = 1'b1;
  assign \A[11][89] [4] = 1'b1;
  assign \A[11][89] [3] = 1'b1;
  assign \A[11][89] [2] = 1'b1;
  assign \A[11][90] [4] = 1'b1;
  assign \A[11][90] [3] = 1'b1;
  assign \A[11][90] [2] = 1'b1;
  assign \A[11][90] [1] = 1'b1;
  assign \A[11][90] [0] = 1'b1;
  assign \A[11][91] [4] = 1'b1;
  assign \A[11][91] [3] = 1'b1;
  assign \A[11][91] [2] = 1'b1;
  assign \A[11][91] [0] = 1'b1;
  assign \A[11][92] [4] = 1'b1;
  assign \A[11][92] [3] = 1'b1;
  assign \A[11][92] [2] = 1'b1;
  assign \A[11][94] [4] = 1'b1;
  assign \A[11][94] [3] = 1'b1;
  assign \A[11][94] [2] = 1'b1;
  assign \A[11][94] [0] = 1'b1;
  assign \A[11][96] [1] = 1'b1;
  assign \A[11][97] [1] = 1'b1;
  assign \A[11][98] [4] = 1'b1;
  assign \A[11][98] [3] = 1'b1;
  assign \A[11][98] [2] = 1'b1;
  assign \A[11][98] [1] = 1'b1;
  assign \A[11][99] [4] = 1'b1;
  assign \A[11][99] [3] = 1'b1;
  assign \A[11][99] [2] = 1'b1;
  assign \A[11][99] [1] = 1'b1;
  assign \A[11][99] [0] = 1'b1;
  assign \A[11][100] [1] = 1'b1;
  assign \A[11][100] [0] = 1'b1;
  assign \A[11][101] [4] = 1'b1;
  assign \A[11][101] [3] = 1'b1;
  assign \A[11][101] [2] = 1'b1;
  assign \A[11][101] [0] = 1'b1;
  assign \A[11][102] [4] = 1'b1;
  assign \A[11][102] [3] = 1'b1;
  assign \A[11][102] [2] = 1'b1;
  assign \A[11][102] [1] = 1'b1;
  assign \A[11][103] [4] = 1'b1;
  assign \A[11][103] [3] = 1'b1;
  assign \A[11][103] [2] = 1'b1;
  assign \A[11][103] [1] = 1'b1;
  assign \A[11][103] [0] = 1'b1;
  assign \A[11][104] [4] = 1'b1;
  assign \A[11][104] [3] = 1'b1;
  assign \A[11][104] [2] = 1'b1;
  assign \A[11][104] [1] = 1'b1;
  assign \A[11][104] [0] = 1'b1;
  assign \A[11][105] [4] = 1'b1;
  assign \A[11][105] [3] = 1'b1;
  assign \A[11][105] [2] = 1'b1;
  assign \A[11][105] [1] = 1'b1;
  assign \A[11][105] [0] = 1'b1;
  assign \A[11][107] [4] = 1'b1;
  assign \A[11][107] [3] = 1'b1;
  assign \A[11][107] [2] = 1'b1;
  assign \A[11][107] [0] = 1'b1;
  assign \A[11][108] [1] = 1'b1;
  assign \A[11][110] [4] = 1'b1;
  assign \A[11][110] [3] = 1'b1;
  assign \A[11][110] [2] = 1'b1;
  assign \A[11][110] [1] = 1'b1;
  assign \A[11][112] [0] = 1'b1;
  assign \A[11][114] [0] = 1'b1;
  assign \A[11][115] [1] = 1'b1;
  assign \A[11][116] [0] = 1'b1;
  assign \A[11][117] [0] = 1'b1;
  assign \A[11][118] [4] = 1'b1;
  assign \A[11][118] [3] = 1'b1;
  assign \A[11][118] [2] = 1'b1;
  assign \A[11][118] [1] = 1'b1;
  assign \A[11][118] [0] = 1'b1;
  assign \A[11][120] [0] = 1'b1;
  assign \A[11][121] [4] = 1'b1;
  assign \A[11][121] [3] = 1'b1;
  assign \A[11][121] [2] = 1'b1;
  assign \A[11][121] [1] = 1'b1;
  assign \A[11][121] [0] = 1'b1;
  assign \A[11][122] [0] = 1'b1;
  assign \A[11][123] [4] = 1'b1;
  assign \A[11][123] [3] = 1'b1;
  assign \A[11][123] [2] = 1'b1;
  assign \A[11][123] [1] = 1'b1;
  assign \A[11][123] [0] = 1'b1;
  assign \A[11][124] [2] = 1'b1;
  assign \A[11][126] [4] = 1'b1;
  assign \A[11][126] [3] = 1'b1;
  assign \A[11][126] [2] = 1'b1;
  assign \A[11][126] [0] = 1'b1;
  assign \A[11][127] [4] = 1'b1;
  assign \A[11][127] [3] = 1'b1;
  assign \A[11][127] [2] = 1'b1;
  assign \A[11][127] [1] = 1'b1;
  assign \A[11][128] [1] = 1'b1;
  assign \A[11][128] [0] = 1'b1;
  assign \A[11][129] [2] = 1'b1;
  assign \A[11][131] [4] = 1'b1;
  assign \A[11][131] [3] = 1'b1;
  assign \A[11][131] [2] = 1'b1;
  assign \A[11][131] [1] = 1'b1;
  assign \A[11][131] [0] = 1'b1;
  assign \A[11][132] [0] = 1'b1;
  assign \A[11][133] [4] = 1'b1;
  assign \A[11][133] [3] = 1'b1;
  assign \A[11][133] [2] = 1'b1;
  assign \A[11][133] [1] = 1'b1;
  assign \A[11][133] [0] = 1'b1;
  assign \A[11][134] [0] = 1'b1;
  assign \A[11][136] [1] = 1'b1;
  assign \A[11][137] [1] = 1'b1;
  assign \A[11][138] [4] = 1'b1;
  assign \A[11][138] [3] = 1'b1;
  assign \A[11][138] [2] = 1'b1;
  assign \A[11][138] [1] = 1'b1;
  assign \A[11][138] [0] = 1'b1;
  assign \A[11][139] [0] = 1'b1;
  assign \A[11][140] [4] = 1'b1;
  assign \A[11][140] [3] = 1'b1;
  assign \A[11][140] [2] = 1'b1;
  assign \A[11][140] [1] = 1'b1;
  assign \A[11][141] [1] = 1'b1;
  assign \A[11][141] [0] = 1'b1;
  assign \A[11][142] [1] = 1'b1;
  assign \A[11][143] [1] = 1'b1;
  assign \A[11][145] [1] = 1'b1;
  assign \A[11][145] [0] = 1'b1;
  assign \A[11][146] [2] = 1'b1;
  assign \A[11][146] [0] = 1'b1;
  assign \A[11][147] [1] = 1'b1;
  assign \A[11][148] [0] = 1'b1;
  assign \A[11][149] [4] = 1'b1;
  assign \A[11][149] [3] = 1'b1;
  assign \A[11][149] [2] = 1'b1;
  assign \A[11][149] [1] = 1'b1;
  assign \A[11][149] [0] = 1'b1;
  assign \A[11][150] [4] = 1'b1;
  assign \A[11][150] [3] = 1'b1;
  assign \A[11][150] [2] = 1'b1;
  assign \A[11][150] [1] = 1'b1;
  assign \A[11][151] [1] = 1'b1;
  assign \A[11][152] [0] = 1'b1;
  assign \A[11][153] [4] = 1'b1;
  assign \A[11][153] [3] = 1'b1;
  assign \A[11][153] [2] = 1'b1;
  assign \A[11][153] [1] = 1'b1;
  assign \A[11][155] [1] = 1'b1;
  assign \A[11][156] [4] = 1'b1;
  assign \A[11][156] [3] = 1'b1;
  assign \A[11][156] [2] = 1'b1;
  assign \A[11][156] [1] = 1'b1;
  assign \A[11][156] [0] = 1'b1;
  assign \A[11][157] [1] = 1'b1;
  assign \A[11][158] [4] = 1'b1;
  assign \A[11][158] [3] = 1'b1;
  assign \A[11][158] [2] = 1'b1;
  assign \A[11][158] [1] = 1'b1;
  assign \A[11][158] [0] = 1'b1;
  assign \A[11][159] [0] = 1'b1;
  assign \A[11][160] [4] = 1'b1;
  assign \A[11][160] [3] = 1'b1;
  assign \A[11][160] [2] = 1'b1;
  assign \A[11][160] [1] = 1'b1;
  assign \A[11][160] [0] = 1'b1;
  assign \A[11][161] [2] = 1'b1;
  assign \A[11][161] [1] = 1'b1;
  assign \A[11][161] [0] = 1'b1;
  assign \A[11][162] [0] = 1'b1;
  assign \A[11][163] [1] = 1'b1;
  assign \A[11][164] [4] = 1'b1;
  assign \A[11][164] [3] = 1'b1;
  assign \A[11][164] [2] = 1'b1;
  assign \A[11][164] [1] = 1'b1;
  assign \A[11][165] [4] = 1'b1;
  assign \A[11][165] [3] = 1'b1;
  assign \A[11][165] [2] = 1'b1;
  assign \A[11][165] [1] = 1'b1;
  assign \A[11][165] [0] = 1'b1;
  assign \A[11][166] [4] = 1'b1;
  assign \A[11][166] [3] = 1'b1;
  assign \A[11][166] [2] = 1'b1;
  assign \A[11][166] [1] = 1'b1;
  assign \A[11][166] [0] = 1'b1;
  assign \A[11][167] [1] = 1'b1;
  assign \A[11][167] [0] = 1'b1;
  assign \A[11][168] [1] = 1'b1;
  assign \A[11][168] [0] = 1'b1;
  assign \A[11][169] [0] = 1'b1;
  assign \A[11][170] [2] = 1'b1;
  assign \A[11][171] [0] = 1'b1;
  assign \A[11][172] [0] = 1'b1;
  assign \A[11][173] [1] = 1'b1;
  assign \A[11][174] [1] = 1'b1;
  assign \A[11][175] [1] = 1'b1;
  assign \A[11][176] [1] = 1'b1;
  assign \A[11][177] [1] = 1'b1;
  assign \A[11][179] [0] = 1'b1;
  assign \A[11][180] [1] = 1'b1;
  assign \A[11][181] [0] = 1'b1;
  assign \A[11][182] [4] = 1'b1;
  assign \A[11][182] [3] = 1'b1;
  assign \A[11][182] [2] = 1'b1;
  assign \A[11][182] [1] = 1'b1;
  assign \A[11][182] [0] = 1'b1;
  assign \A[11][183] [0] = 1'b1;
  assign \A[11][185] [1] = 1'b1;
  assign \A[11][187] [1] = 1'b1;
  assign \A[11][188] [4] = 1'b1;
  assign \A[11][188] [3] = 1'b1;
  assign \A[11][188] [2] = 1'b1;
  assign \A[11][188] [1] = 1'b1;
  assign \A[11][188] [0] = 1'b1;
  assign \A[11][189] [1] = 1'b1;
  assign \A[11][190] [0] = 1'b1;
  assign \A[11][193] [0] = 1'b1;
  assign \A[11][194] [1] = 1'b1;
  assign \A[11][194] [0] = 1'b1;
  assign \A[11][195] [0] = 1'b1;
  assign \A[11][196] [0] = 1'b1;
  assign \A[11][197] [1] = 1'b1;
  assign \A[11][198] [4] = 1'b1;
  assign \A[11][198] [3] = 1'b1;
  assign \A[11][198] [2] = 1'b1;
  assign \A[11][198] [1] = 1'b1;
  assign \A[11][199] [1] = 1'b1;
  assign \A[11][199] [0] = 1'b1;
  assign \A[11][200] [4] = 1'b1;
  assign \A[11][200] [3] = 1'b1;
  assign \A[11][200] [2] = 1'b1;
  assign \A[11][200] [1] = 1'b1;
  assign \A[11][202] [1] = 1'b1;
  assign \A[11][205] [4] = 1'b1;
  assign \A[11][205] [3] = 1'b1;
  assign \A[11][205] [2] = 1'b1;
  assign \A[11][205] [1] = 1'b1;
  assign \A[11][205] [0] = 1'b1;
  assign \A[11][207] [0] = 1'b1;
  assign \A[11][208] [0] = 1'b1;
  assign \A[11][209] [4] = 1'b1;
  assign \A[11][209] [3] = 1'b1;
  assign \A[11][209] [2] = 1'b1;
  assign \A[11][209] [1] = 1'b1;
  assign \A[11][209] [0] = 1'b1;
  assign \A[11][210] [4] = 1'b1;
  assign \A[11][210] [3] = 1'b1;
  assign \A[11][210] [2] = 1'b1;
  assign \A[11][210] [1] = 1'b1;
  assign \A[11][210] [0] = 1'b1;
  assign \A[11][211] [0] = 1'b1;
  assign \A[11][212] [4] = 1'b1;
  assign \A[11][212] [3] = 1'b1;
  assign \A[11][212] [2] = 1'b1;
  assign \A[11][213] [4] = 1'b1;
  assign \A[11][213] [3] = 1'b1;
  assign \A[11][213] [2] = 1'b1;
  assign \A[11][213] [1] = 1'b1;
  assign \A[11][213] [0] = 1'b1;
  assign \A[11][215] [0] = 1'b1;
  assign \A[11][216] [4] = 1'b1;
  assign \A[11][216] [3] = 1'b1;
  assign \A[11][216] [2] = 1'b1;
  assign \A[11][216] [1] = 1'b1;
  assign \A[11][216] [0] = 1'b1;
  assign \A[11][217] [0] = 1'b1;
  assign \A[11][218] [4] = 1'b1;
  assign \A[11][218] [3] = 1'b1;
  assign \A[11][218] [2] = 1'b1;
  assign \A[11][218] [1] = 1'b1;
  assign \A[11][220] [4] = 1'b1;
  assign \A[11][220] [3] = 1'b1;
  assign \A[11][220] [2] = 1'b1;
  assign \A[11][220] [1] = 1'b1;
  assign \A[11][220] [0] = 1'b1;
  assign \A[11][221] [0] = 1'b1;
  assign \A[11][222] [4] = 1'b1;
  assign \A[11][222] [3] = 1'b1;
  assign \A[11][222] [2] = 1'b1;
  assign \A[11][222] [0] = 1'b1;
  assign \A[11][223] [4] = 1'b1;
  assign \A[11][223] [3] = 1'b1;
  assign \A[11][223] [2] = 1'b1;
  assign \A[11][223] [1] = 1'b1;
  assign \A[11][223] [0] = 1'b1;
  assign \A[11][224] [0] = 1'b1;
  assign \A[11][225] [0] = 1'b1;
  assign \A[11][226] [4] = 1'b1;
  assign \A[11][226] [3] = 1'b1;
  assign \A[11][226] [2] = 1'b1;
  assign \A[11][226] [1] = 1'b1;
  assign \A[11][227] [4] = 1'b1;
  assign \A[11][227] [3] = 1'b1;
  assign \A[11][227] [2] = 1'b1;
  assign \A[11][227] [1] = 1'b1;
  assign \A[11][227] [0] = 1'b1;
  assign \A[11][229] [1] = 1'b1;
  assign \A[11][229] [0] = 1'b1;
  assign \A[11][230] [4] = 1'b1;
  assign \A[11][230] [3] = 1'b1;
  assign \A[11][230] [2] = 1'b1;
  assign \A[11][230] [1] = 1'b1;
  assign \A[11][233] [4] = 1'b1;
  assign \A[11][233] [3] = 1'b1;
  assign \A[11][233] [2] = 1'b1;
  assign \A[11][233] [1] = 1'b1;
  assign \A[11][233] [0] = 1'b1;
  assign \A[11][235] [0] = 1'b1;
  assign \A[11][238] [4] = 1'b1;
  assign \A[11][238] [3] = 1'b1;
  assign \A[11][238] [2] = 1'b1;
  assign \A[11][238] [1] = 1'b1;
  assign \A[11][238] [0] = 1'b1;
  assign \A[11][239] [4] = 1'b1;
  assign \A[11][239] [3] = 1'b1;
  assign \A[11][239] [2] = 1'b1;
  assign \A[11][239] [1] = 1'b1;
  assign \A[11][240] [4] = 1'b1;
  assign \A[11][240] [3] = 1'b1;
  assign \A[11][240] [2] = 1'b1;
  assign \A[11][240] [1] = 1'b1;
  assign \A[11][240] [0] = 1'b1;
  assign \A[11][241] [4] = 1'b1;
  assign \A[11][241] [3] = 1'b1;
  assign \A[11][241] [2] = 1'b1;
  assign \A[11][241] [1] = 1'b1;
  assign \A[11][241] [0] = 1'b1;
  assign \A[11][242] [0] = 1'b1;
  assign \A[11][243] [4] = 1'b1;
  assign \A[11][243] [3] = 1'b1;
  assign \A[11][243] [2] = 1'b1;
  assign \A[11][243] [1] = 1'b1;
  assign \A[11][243] [0] = 1'b1;
  assign \A[11][244] [4] = 1'b1;
  assign \A[11][244] [3] = 1'b1;
  assign \A[11][244] [2] = 1'b1;
  assign \A[11][244] [0] = 1'b1;
  assign \A[11][245] [4] = 1'b1;
  assign \A[11][245] [3] = 1'b1;
  assign \A[11][245] [2] = 1'b1;
  assign \A[11][245] [1] = 1'b1;
  assign \A[11][245] [0] = 1'b1;
  assign \A[11][246] [4] = 1'b1;
  assign \A[11][246] [3] = 1'b1;
  assign \A[11][246] [2] = 1'b1;
  assign \A[11][246] [1] = 1'b1;
  assign \A[11][246] [0] = 1'b1;
  assign \A[11][247] [0] = 1'b1;
  assign \A[11][251] [4] = 1'b1;
  assign \A[11][251] [3] = 1'b1;
  assign \A[11][251] [2] = 1'b1;
  assign \A[11][251] [1] = 1'b1;
  assign \A[11][252] [4] = 1'b1;
  assign \A[11][252] [3] = 1'b1;
  assign \A[11][252] [2] = 1'b1;
  assign \A[11][252] [1] = 1'b1;
  assign \A[11][252] [0] = 1'b1;
  assign \A[11][254] [4] = 1'b1;
  assign \A[11][254] [3] = 1'b1;
  assign \A[11][254] [2] = 1'b1;
  assign \A[11][254] [1] = 1'b1;
  assign \A[11][255] [4] = 1'b1;
  assign \A[11][255] [3] = 1'b1;
  assign \A[11][255] [2] = 1'b1;
  assign \A[11][255] [1] = 1'b1;
  assign \A[11][255] [0] = 1'b1;
  assign \A[12][0] [0] = 1'b1;
  assign \A[12][1] [4] = 1'b1;
  assign \A[12][1] [3] = 1'b1;
  assign \A[12][1] [2] = 1'b1;
  assign \A[12][1] [1] = 1'b1;
  assign \A[12][2] [4] = 1'b1;
  assign \A[12][2] [3] = 1'b1;
  assign \A[12][2] [2] = 1'b1;
  assign \A[12][2] [1] = 1'b1;
  assign \A[12][4] [0] = 1'b1;
  assign \A[12][5] [1] = 1'b1;
  assign \A[12][6] [4] = 1'b1;
  assign \A[12][6] [3] = 1'b1;
  assign \A[12][6] [2] = 1'b1;
  assign \A[12][6] [1] = 1'b1;
  assign \A[12][8] [4] = 1'b1;
  assign \A[12][8] [3] = 1'b1;
  assign \A[12][8] [2] = 1'b1;
  assign \A[12][8] [0] = 1'b1;
  assign \A[12][9] [4] = 1'b1;
  assign \A[12][9] [3] = 1'b1;
  assign \A[12][9] [2] = 1'b1;
  assign \A[12][9] [1] = 1'b1;
  assign \A[12][9] [0] = 1'b1;
  assign \A[12][10] [4] = 1'b1;
  assign \A[12][10] [3] = 1'b1;
  assign \A[12][10] [2] = 1'b1;
  assign \A[12][10] [1] = 1'b1;
  assign \A[12][11] [4] = 1'b1;
  assign \A[12][11] [3] = 1'b1;
  assign \A[12][11] [2] = 1'b1;
  assign \A[12][11] [1] = 1'b1;
  assign \A[12][11] [0] = 1'b1;
  assign \A[12][13] [1] = 1'b1;
  assign \A[12][14] [0] = 1'b1;
  assign \A[12][15] [4] = 1'b1;
  assign \A[12][15] [3] = 1'b1;
  assign \A[12][15] [2] = 1'b1;
  assign \A[12][15] [1] = 1'b1;
  assign \A[12][15] [0] = 1'b1;
  assign \A[12][16] [4] = 1'b1;
  assign \A[12][16] [3] = 1'b1;
  assign \A[12][16] [2] = 1'b1;
  assign \A[12][16] [1] = 1'b1;
  assign \A[12][16] [0] = 1'b1;
  assign \A[12][17] [4] = 1'b1;
  assign \A[12][17] [3] = 1'b1;
  assign \A[12][17] [2] = 1'b1;
  assign \A[12][17] [1] = 1'b1;
  assign \A[12][17] [0] = 1'b1;
  assign \A[12][18] [4] = 1'b1;
  assign \A[12][18] [3] = 1'b1;
  assign \A[12][18] [2] = 1'b1;
  assign \A[12][18] [1] = 1'b1;
  assign \A[12][18] [0] = 1'b1;
  assign \A[12][21] [0] = 1'b1;
  assign \A[12][22] [4] = 1'b1;
  assign \A[12][22] [3] = 1'b1;
  assign \A[12][22] [2] = 1'b1;
  assign \A[12][22] [1] = 1'b1;
  assign \A[12][22] [0] = 1'b1;
  assign \A[12][23] [0] = 1'b1;
  assign \A[12][25] [4] = 1'b1;
  assign \A[12][25] [3] = 1'b1;
  assign \A[12][25] [2] = 1'b1;
  assign \A[12][25] [1] = 1'b1;
  assign \A[12][25] [0] = 1'b1;
  assign \A[12][26] [4] = 1'b1;
  assign \A[12][26] [3] = 1'b1;
  assign \A[12][26] [2] = 1'b1;
  assign \A[12][26] [1] = 1'b1;
  assign \A[12][26] [0] = 1'b1;
  assign \A[12][27] [0] = 1'b1;
  assign \A[12][29] [0] = 1'b1;
  assign \A[12][30] [4] = 1'b1;
  assign \A[12][30] [3] = 1'b1;
  assign \A[12][30] [2] = 1'b1;
  assign \A[12][30] [1] = 1'b1;
  assign \A[12][31] [4] = 1'b1;
  assign \A[12][31] [3] = 1'b1;
  assign \A[12][31] [2] = 1'b1;
  assign \A[12][31] [1] = 1'b1;
  assign \A[12][32] [0] = 1'b1;
  assign \A[12][33] [0] = 1'b1;
  assign \A[12][37] [0] = 1'b1;
  assign \A[12][39] [4] = 1'b1;
  assign \A[12][39] [3] = 1'b1;
  assign \A[12][39] [2] = 1'b1;
  assign \A[12][39] [1] = 1'b1;
  assign \A[12][39] [0] = 1'b1;
  assign \A[12][40] [4] = 1'b1;
  assign \A[12][40] [3] = 1'b1;
  assign \A[12][40] [2] = 1'b1;
  assign \A[12][40] [1] = 1'b1;
  assign \A[12][40] [0] = 1'b1;
  assign \A[12][41] [0] = 1'b1;
  assign \A[12][42] [0] = 1'b1;
  assign \A[12][43] [0] = 1'b1;
  assign \A[12][44] [4] = 1'b1;
  assign \A[12][44] [3] = 1'b1;
  assign \A[12][44] [2] = 1'b1;
  assign \A[12][44] [1] = 1'b1;
  assign \A[12][44] [0] = 1'b1;
  assign \A[12][46] [1] = 1'b1;
  assign \A[12][47] [4] = 1'b1;
  assign \A[12][47] [3] = 1'b1;
  assign \A[12][47] [2] = 1'b1;
  assign \A[12][47] [1] = 1'b1;
  assign \A[12][47] [0] = 1'b1;
  assign \A[12][48] [4] = 1'b1;
  assign \A[12][48] [3] = 1'b1;
  assign \A[12][48] [2] = 1'b1;
  assign \A[12][48] [1] = 1'b1;
  assign \A[12][48] [0] = 1'b1;
  assign \A[12][49] [0] = 1'b1;
  assign \A[12][50] [4] = 1'b1;
  assign \A[12][50] [3] = 1'b1;
  assign \A[12][50] [2] = 1'b1;
  assign \A[12][50] [0] = 1'b1;
  assign \A[12][51] [4] = 1'b1;
  assign \A[12][51] [3] = 1'b1;
  assign \A[12][51] [2] = 1'b1;
  assign \A[12][51] [1] = 1'b1;
  assign \A[12][52] [0] = 1'b1;
  assign \A[12][53] [1] = 1'b1;
  assign \A[12][53] [0] = 1'b1;
  assign \A[12][54] [4] = 1'b1;
  assign \A[12][54] [3] = 1'b1;
  assign \A[12][54] [2] = 1'b1;
  assign \A[12][54] [1] = 1'b1;
  assign \A[12][55] [0] = 1'b1;
  assign \A[12][56] [1] = 1'b1;
  assign \A[12][58] [0] = 1'b1;
  assign \A[12][59] [4] = 1'b1;
  assign \A[12][59] [3] = 1'b1;
  assign \A[12][59] [2] = 1'b1;
  assign \A[12][59] [1] = 1'b1;
  assign \A[12][59] [0] = 1'b1;
  assign \A[12][60] [4] = 1'b1;
  assign \A[12][60] [3] = 1'b1;
  assign \A[12][60] [2] = 1'b1;
  assign \A[12][60] [1] = 1'b1;
  assign \A[12][60] [0] = 1'b1;
  assign \A[12][62] [1] = 1'b1;
  assign \A[12][63] [0] = 1'b1;
  assign \A[12][64] [1] = 1'b1;
  assign \A[12][64] [0] = 1'b1;
  assign \A[12][66] [0] = 1'b1;
  assign \A[12][68] [0] = 1'b1;
  assign \A[12][69] [1] = 1'b1;
  assign \A[12][69] [0] = 1'b1;
  assign \A[12][70] [4] = 1'b1;
  assign \A[12][70] [3] = 1'b1;
  assign \A[12][70] [2] = 1'b1;
  assign \A[12][70] [1] = 1'b1;
  assign \A[12][71] [4] = 1'b1;
  assign \A[12][71] [3] = 1'b1;
  assign \A[12][71] [2] = 1'b1;
  assign \A[12][71] [0] = 1'b1;
  assign \A[12][72] [0] = 1'b1;
  assign \A[12][74] [4] = 1'b1;
  assign \A[12][74] [3] = 1'b1;
  assign \A[12][74] [2] = 1'b1;
  assign \A[12][74] [0] = 1'b1;
  assign \A[12][75] [4] = 1'b1;
  assign \A[12][75] [3] = 1'b1;
  assign \A[12][75] [2] = 1'b1;
  assign \A[12][75] [1] = 1'b1;
  assign \A[12][75] [0] = 1'b1;
  assign \A[12][76] [4] = 1'b1;
  assign \A[12][76] [3] = 1'b1;
  assign \A[12][76] [2] = 1'b1;
  assign \A[12][76] [1] = 1'b1;
  assign \A[12][76] [0] = 1'b1;
  assign \A[12][77] [0] = 1'b1;
  assign \A[12][78] [4] = 1'b1;
  assign \A[12][78] [3] = 1'b1;
  assign \A[12][78] [2] = 1'b1;
  assign \A[12][78] [1] = 1'b1;
  assign \A[12][79] [4] = 1'b1;
  assign \A[12][79] [3] = 1'b1;
  assign \A[12][79] [2] = 1'b1;
  assign \A[12][79] [1] = 1'b1;
  assign \A[12][79] [0] = 1'b1;
  assign \A[12][80] [0] = 1'b1;
  assign \A[12][81] [4] = 1'b1;
  assign \A[12][81] [3] = 1'b1;
  assign \A[12][81] [2] = 1'b1;
  assign \A[12][81] [1] = 1'b1;
  assign \A[12][82] [4] = 1'b1;
  assign \A[12][82] [3] = 1'b1;
  assign \A[12][82] [2] = 1'b1;
  assign \A[12][82] [1] = 1'b1;
  assign \A[12][82] [0] = 1'b1;
  assign \A[12][83] [4] = 1'b1;
  assign \A[12][83] [3] = 1'b1;
  assign \A[12][83] [2] = 1'b1;
  assign \A[12][83] [1] = 1'b1;
  assign \A[12][84] [1] = 1'b1;
  assign \A[12][84] [0] = 1'b1;
  assign \A[12][85] [1] = 1'b1;
  assign \A[12][86] [0] = 1'b1;
  assign \A[12][87] [4] = 1'b1;
  assign \A[12][87] [3] = 1'b1;
  assign \A[12][87] [2] = 1'b1;
  assign \A[12][87] [1] = 1'b1;
  assign \A[12][87] [0] = 1'b1;
  assign \A[12][88] [0] = 1'b1;
  assign \A[12][90] [0] = 1'b1;
  assign \A[12][91] [4] = 1'b1;
  assign \A[12][91] [3] = 1'b1;
  assign \A[12][91] [2] = 1'b1;
  assign \A[12][91] [1] = 1'b1;
  assign \A[12][91] [0] = 1'b1;
  assign \A[12][92] [4] = 1'b1;
  assign \A[12][92] [3] = 1'b1;
  assign \A[12][92] [2] = 1'b1;
  assign \A[12][92] [1] = 1'b1;
  assign \A[12][93] [4] = 1'b1;
  assign \A[12][93] [3] = 1'b1;
  assign \A[12][93] [2] = 1'b1;
  assign \A[12][93] [1] = 1'b1;
  assign \A[12][93] [0] = 1'b1;
  assign \A[12][94] [0] = 1'b1;
  assign \A[12][95] [4] = 1'b1;
  assign \A[12][95] [3] = 1'b1;
  assign \A[12][95] [2] = 1'b1;
  assign \A[12][95] [1] = 1'b1;
  assign \A[12][95] [0] = 1'b1;
  assign \A[12][96] [4] = 1'b1;
  assign \A[12][96] [3] = 1'b1;
  assign \A[12][96] [2] = 1'b1;
  assign \A[12][96] [1] = 1'b1;
  assign \A[12][96] [0] = 1'b1;
  assign \A[12][98] [4] = 1'b1;
  assign \A[12][98] [3] = 1'b1;
  assign \A[12][98] [2] = 1'b1;
  assign \A[12][98] [1] = 1'b1;
  assign \A[12][98] [0] = 1'b1;
  assign \A[12][100] [4] = 1'b1;
  assign \A[12][100] [3] = 1'b1;
  assign \A[12][100] [2] = 1'b1;
  assign \A[12][100] [1] = 1'b1;
  assign \A[12][101] [4] = 1'b1;
  assign \A[12][101] [3] = 1'b1;
  assign \A[12][101] [2] = 1'b1;
  assign \A[12][101] [1] = 1'b1;
  assign \A[12][101] [0] = 1'b1;
  assign \A[12][102] [0] = 1'b1;
  assign \A[12][104] [0] = 1'b1;
  assign \A[12][105] [1] = 1'b1;
  assign \A[12][106] [4] = 1'b1;
  assign \A[12][106] [3] = 1'b1;
  assign \A[12][106] [2] = 1'b1;
  assign \A[12][106] [1] = 1'b1;
  assign \A[12][108] [0] = 1'b1;
  assign \A[12][110] [0] = 1'b1;
  assign \A[12][111] [1] = 1'b1;
  assign \A[12][112] [0] = 1'b1;
  assign \A[12][113] [1] = 1'b1;
  assign \A[12][114] [1] = 1'b1;
  assign \A[12][115] [4] = 1'b1;
  assign \A[12][115] [3] = 1'b1;
  assign \A[12][115] [2] = 1'b1;
  assign \A[12][115] [1] = 1'b1;
  assign \A[12][116] [4] = 1'b1;
  assign \A[12][116] [3] = 1'b1;
  assign \A[12][116] [2] = 1'b1;
  assign \A[12][116] [0] = 1'b1;
  assign \A[12][117] [0] = 1'b1;
  assign \A[12][118] [4] = 1'b1;
  assign \A[12][118] [3] = 1'b1;
  assign \A[12][118] [2] = 1'b1;
  assign \A[12][118] [1] = 1'b1;
  assign \A[12][118] [0] = 1'b1;
  assign \A[12][120] [1] = 1'b1;
  assign \A[12][121] [0] = 1'b1;
  assign \A[12][122] [4] = 1'b1;
  assign \A[12][122] [3] = 1'b1;
  assign \A[12][122] [2] = 1'b1;
  assign \A[12][122] [0] = 1'b1;
  assign \A[12][123] [4] = 1'b1;
  assign \A[12][123] [3] = 1'b1;
  assign \A[12][123] [2] = 1'b1;
  assign \A[12][123] [1] = 1'b1;
  assign \A[12][123] [0] = 1'b1;
  assign \A[12][124] [4] = 1'b1;
  assign \A[12][124] [3] = 1'b1;
  assign \A[12][124] [2] = 1'b1;
  assign \A[12][124] [1] = 1'b1;
  assign \A[12][125] [4] = 1'b1;
  assign \A[12][125] [3] = 1'b1;
  assign \A[12][125] [2] = 1'b1;
  assign \A[12][125] [1] = 1'b1;
  assign \A[12][126] [1] = 1'b1;
  assign \A[12][127] [4] = 1'b1;
  assign \A[12][127] [3] = 1'b1;
  assign \A[12][127] [2] = 1'b1;
  assign \A[12][127] [1] = 1'b1;
  assign \A[12][128] [4] = 1'b1;
  assign \A[12][128] [3] = 1'b1;
  assign \A[12][128] [2] = 1'b1;
  assign \A[12][128] [0] = 1'b1;
  assign \A[12][129] [4] = 1'b1;
  assign \A[12][129] [3] = 1'b1;
  assign \A[12][129] [2] = 1'b1;
  assign \A[12][129] [1] = 1'b1;
  assign \A[12][130] [4] = 1'b1;
  assign \A[12][130] [3] = 1'b1;
  assign \A[12][130] [2] = 1'b1;
  assign \A[12][130] [1] = 1'b1;
  assign \A[12][130] [0] = 1'b1;
  assign \A[12][131] [4] = 1'b1;
  assign \A[12][131] [3] = 1'b1;
  assign \A[12][131] [2] = 1'b1;
  assign \A[12][131] [1] = 1'b1;
  assign \A[12][131] [0] = 1'b1;
  assign \A[12][132] [4] = 1'b1;
  assign \A[12][132] [3] = 1'b1;
  assign \A[12][132] [2] = 1'b1;
  assign \A[12][132] [1] = 1'b1;
  assign \A[12][134] [1] = 1'b1;
  assign \A[12][134] [0] = 1'b1;
  assign \A[12][135] [1] = 1'b1;
  assign \A[12][140] [1] = 1'b1;
  assign \A[12][140] [0] = 1'b1;
  assign \A[12][141] [1] = 1'b1;
  assign \A[12][141] [0] = 1'b1;
  assign \A[12][142] [0] = 1'b1;
  assign \A[12][143] [1] = 1'b1;
  assign \A[12][144] [0] = 1'b1;
  assign \A[12][146] [0] = 1'b1;
  assign \A[12][147] [0] = 1'b1;
  assign \A[12][148] [4] = 1'b1;
  assign \A[12][148] [3] = 1'b1;
  assign \A[12][148] [2] = 1'b1;
  assign \A[12][148] [1] = 1'b1;
  assign \A[12][148] [0] = 1'b1;
  assign \A[12][150] [2] = 1'b1;
  assign \A[12][151] [1] = 1'b1;
  assign \A[12][151] [0] = 1'b1;
  assign \A[12][152] [4] = 1'b1;
  assign \A[12][152] [3] = 1'b1;
  assign \A[12][152] [2] = 1'b1;
  assign \A[12][152] [1] = 1'b1;
  assign \A[12][152] [0] = 1'b1;
  assign \A[12][153] [1] = 1'b1;
  assign \A[12][154] [1] = 1'b1;
  assign \A[12][155] [4] = 1'b1;
  assign \A[12][155] [3] = 1'b1;
  assign \A[12][155] [2] = 1'b1;
  assign \A[12][155] [0] = 1'b1;
  assign \A[12][156] [0] = 1'b1;
  assign \A[12][158] [4] = 1'b1;
  assign \A[12][158] [3] = 1'b1;
  assign \A[12][158] [2] = 1'b1;
  assign \A[12][158] [1] = 1'b1;
  assign \A[12][160] [0] = 1'b1;
  assign \A[12][163] [4] = 1'b1;
  assign \A[12][163] [3] = 1'b1;
  assign \A[12][163] [2] = 1'b1;
  assign \A[12][163] [1] = 1'b1;
  assign \A[12][164] [1] = 1'b1;
  assign \A[12][165] [1] = 1'b1;
  assign \A[12][167] [1] = 1'b1;
  assign \A[12][168] [0] = 1'b1;
  assign \A[12][170] [1] = 1'b1;
  assign \A[12][172] [4] = 1'b1;
  assign \A[12][172] [3] = 1'b1;
  assign \A[12][172] [2] = 1'b1;
  assign \A[12][172] [1] = 1'b1;
  assign \A[12][172] [0] = 1'b1;
  assign \A[12][173] [4] = 1'b1;
  assign \A[12][173] [3] = 1'b1;
  assign \A[12][173] [2] = 1'b1;
  assign \A[12][173] [1] = 1'b1;
  assign \A[12][173] [0] = 1'b1;
  assign \A[12][176] [4] = 1'b1;
  assign \A[12][176] [3] = 1'b1;
  assign \A[12][176] [2] = 1'b1;
  assign \A[12][176] [1] = 1'b1;
  assign \A[12][177] [4] = 1'b1;
  assign \A[12][177] [3] = 1'b1;
  assign \A[12][177] [2] = 1'b1;
  assign \A[12][177] [1] = 1'b1;
  assign \A[12][177] [0] = 1'b1;
  assign \A[12][178] [0] = 1'b1;
  assign \A[12][179] [4] = 1'b1;
  assign \A[12][179] [3] = 1'b1;
  assign \A[12][179] [2] = 1'b1;
  assign \A[12][179] [1] = 1'b1;
  assign \A[12][180] [4] = 1'b1;
  assign \A[12][180] [3] = 1'b1;
  assign \A[12][180] [2] = 1'b1;
  assign \A[12][180] [1] = 1'b1;
  assign \A[12][180] [0] = 1'b1;
  assign \A[12][181] [4] = 1'b1;
  assign \A[12][181] [3] = 1'b1;
  assign \A[12][181] [2] = 1'b1;
  assign \A[12][181] [1] = 1'b1;
  assign \A[12][181] [0] = 1'b1;
  assign \A[12][185] [1] = 1'b1;
  assign \A[12][187] [4] = 1'b1;
  assign \A[12][187] [3] = 1'b1;
  assign \A[12][187] [2] = 1'b1;
  assign \A[12][187] [1] = 1'b1;
  assign \A[12][188] [1] = 1'b1;
  assign \A[12][189] [4] = 1'b1;
  assign \A[12][189] [3] = 1'b1;
  assign \A[12][189] [2] = 1'b1;
  assign \A[12][189] [1] = 1'b1;
  assign \A[12][189] [0] = 1'b1;
  assign \A[12][190] [4] = 1'b1;
  assign \A[12][190] [3] = 1'b1;
  assign \A[12][190] [2] = 1'b1;
  assign \A[12][190] [0] = 1'b1;
  assign \A[12][191] [4] = 1'b1;
  assign \A[12][191] [3] = 1'b1;
  assign \A[12][191] [2] = 1'b1;
  assign \A[12][191] [1] = 1'b1;
  assign \A[12][191] [0] = 1'b1;
  assign \A[12][192] [1] = 1'b1;
  assign \A[12][194] [0] = 1'b1;
  assign \A[12][195] [0] = 1'b1;
  assign \A[12][196] [4] = 1'b1;
  assign \A[12][196] [3] = 1'b1;
  assign \A[12][196] [2] = 1'b1;
  assign \A[12][196] [0] = 1'b1;
  assign \A[12][198] [1] = 1'b1;
  assign \A[12][199] [4] = 1'b1;
  assign \A[12][199] [3] = 1'b1;
  assign \A[12][199] [2] = 1'b1;
  assign \A[12][199] [1] = 1'b1;
  assign \A[12][199] [0] = 1'b1;
  assign \A[12][200] [0] = 1'b1;
  assign \A[12][202] [0] = 1'b1;
  assign \A[12][203] [4] = 1'b1;
  assign \A[12][203] [3] = 1'b1;
  assign \A[12][203] [2] = 1'b1;
  assign \A[12][203] [1] = 1'b1;
  assign \A[12][203] [0] = 1'b1;
  assign \A[12][205] [4] = 1'b1;
  assign \A[12][205] [3] = 1'b1;
  assign \A[12][205] [2] = 1'b1;
  assign \A[12][205] [1] = 1'b1;
  assign \A[12][206] [4] = 1'b1;
  assign \A[12][206] [3] = 1'b1;
  assign \A[12][206] [2] = 1'b1;
  assign \A[12][206] [1] = 1'b1;
  assign \A[12][206] [0] = 1'b1;
  assign \A[12][207] [1] = 1'b1;
  assign \A[12][207] [0] = 1'b1;
  assign \A[12][210] [4] = 1'b1;
  assign \A[12][210] [3] = 1'b1;
  assign \A[12][210] [2] = 1'b1;
  assign \A[12][210] [0] = 1'b1;
  assign \A[12][213] [4] = 1'b1;
  assign \A[12][213] [3] = 1'b1;
  assign \A[12][213] [2] = 1'b1;
  assign \A[12][213] [1] = 1'b1;
  assign \A[12][214] [0] = 1'b1;
  assign \A[12][215] [4] = 1'b1;
  assign \A[12][215] [3] = 1'b1;
  assign \A[12][215] [2] = 1'b1;
  assign \A[12][215] [1] = 1'b1;
  assign \A[12][215] [0] = 1'b1;
  assign \A[12][217] [0] = 1'b1;
  assign \A[12][218] [4] = 1'b1;
  assign \A[12][218] [3] = 1'b1;
  assign \A[12][218] [2] = 1'b1;
  assign \A[12][218] [1] = 1'b1;
  assign \A[12][219] [4] = 1'b1;
  assign \A[12][219] [3] = 1'b1;
  assign \A[12][219] [2] = 1'b1;
  assign \A[12][219] [1] = 1'b1;
  assign \A[12][219] [0] = 1'b1;
  assign \A[12][220] [1] = 1'b1;
  assign \A[12][221] [1] = 1'b1;
  assign \A[12][221] [0] = 1'b1;
  assign \A[12][223] [4] = 1'b1;
  assign \A[12][223] [3] = 1'b1;
  assign \A[12][223] [2] = 1'b1;
  assign \A[12][223] [1] = 1'b1;
  assign \A[12][223] [0] = 1'b1;
  assign \A[12][224] [0] = 1'b1;
  assign \A[12][225] [4] = 1'b1;
  assign \A[12][225] [3] = 1'b1;
  assign \A[12][225] [2] = 1'b1;
  assign \A[12][225] [1] = 1'b1;
  assign \A[12][225] [0] = 1'b1;
  assign \A[12][226] [4] = 1'b1;
  assign \A[12][226] [3] = 1'b1;
  assign \A[12][226] [2] = 1'b1;
  assign \A[12][226] [1] = 1'b1;
  assign \A[12][226] [0] = 1'b1;
  assign \A[12][227] [0] = 1'b1;
  assign \A[12][229] [4] = 1'b1;
  assign \A[12][229] [3] = 1'b1;
  assign \A[12][229] [2] = 1'b1;
  assign \A[12][229] [1] = 1'b1;
  assign \A[12][229] [0] = 1'b1;
  assign \A[12][231] [4] = 1'b1;
  assign \A[12][231] [3] = 1'b1;
  assign \A[12][231] [2] = 1'b1;
  assign \A[12][231] [1] = 1'b1;
  assign \A[12][231] [0] = 1'b1;
  assign \A[12][232] [4] = 1'b1;
  assign \A[12][232] [3] = 1'b1;
  assign \A[12][232] [2] = 1'b1;
  assign \A[12][232] [0] = 1'b1;
  assign \A[12][233] [0] = 1'b1;
  assign \A[12][234] [4] = 1'b1;
  assign \A[12][234] [3] = 1'b1;
  assign \A[12][234] [2] = 1'b1;
  assign \A[12][234] [1] = 1'b1;
  assign \A[12][235] [0] = 1'b1;
  assign \A[12][236] [4] = 1'b1;
  assign \A[12][236] [3] = 1'b1;
  assign \A[12][236] [2] = 1'b1;
  assign \A[12][236] [1] = 1'b1;
  assign \A[12][236] [0] = 1'b1;
  assign \A[12][237] [4] = 1'b1;
  assign \A[12][237] [3] = 1'b1;
  assign \A[12][237] [2] = 1'b1;
  assign \A[12][237] [1] = 1'b1;
  assign \A[12][239] [4] = 1'b1;
  assign \A[12][239] [3] = 1'b1;
  assign \A[12][239] [2] = 1'b1;
  assign \A[12][239] [1] = 1'b1;
  assign \A[12][240] [4] = 1'b1;
  assign \A[12][240] [3] = 1'b1;
  assign \A[12][240] [2] = 1'b1;
  assign \A[12][240] [1] = 1'b1;
  assign \A[12][240] [0] = 1'b1;
  assign \A[12][242] [1] = 1'b1;
  assign \A[12][243] [0] = 1'b1;
  assign \A[12][244] [0] = 1'b1;
  assign \A[12][249] [4] = 1'b1;
  assign \A[12][249] [3] = 1'b1;
  assign \A[12][249] [2] = 1'b1;
  assign \A[12][249] [1] = 1'b1;
  assign \A[12][250] [1] = 1'b1;
  assign \A[12][251] [2] = 1'b1;
  assign \A[12][252] [4] = 1'b1;
  assign \A[12][252] [3] = 1'b1;
  assign \A[12][252] [2] = 1'b1;
  assign \A[12][252] [1] = 1'b1;
  assign \A[12][252] [0] = 1'b1;
  assign \A[12][253] [4] = 1'b1;
  assign \A[12][253] [3] = 1'b1;
  assign \A[12][253] [2] = 1'b1;
  assign \A[12][253] [1] = 1'b1;
  assign \A[13][1] [4] = 1'b1;
  assign \A[13][1] [3] = 1'b1;
  assign \A[13][1] [2] = 1'b1;
  assign \A[13][1] [1] = 1'b1;
  assign \A[13][1] [0] = 1'b1;
  assign \A[13][2] [4] = 1'b1;
  assign \A[13][2] [3] = 1'b1;
  assign \A[13][2] [2] = 1'b1;
  assign \A[13][2] [1] = 1'b1;
  assign \A[13][2] [0] = 1'b1;
  assign \A[13][3] [0] = 1'b1;
  assign \A[13][4] [2] = 1'b1;
  assign \A[13][5] [4] = 1'b1;
  assign \A[13][5] [3] = 1'b1;
  assign \A[13][5] [2] = 1'b1;
  assign \A[13][5] [1] = 1'b1;
  assign \A[13][6] [0] = 1'b1;
  assign \A[13][7] [4] = 1'b1;
  assign \A[13][7] [3] = 1'b1;
  assign \A[13][7] [2] = 1'b1;
  assign \A[13][7] [1] = 1'b1;
  assign \A[13][7] [0] = 1'b1;
  assign \A[13][8] [0] = 1'b1;
  assign \A[13][9] [0] = 1'b1;
  assign \A[13][11] [4] = 1'b1;
  assign \A[13][11] [3] = 1'b1;
  assign \A[13][11] [2] = 1'b1;
  assign \A[13][11] [1] = 1'b1;
  assign \A[13][11] [0] = 1'b1;
  assign \A[13][12] [0] = 1'b1;
  assign \A[13][13] [4] = 1'b1;
  assign \A[13][13] [3] = 1'b1;
  assign \A[13][13] [2] = 1'b1;
  assign \A[13][13] [1] = 1'b1;
  assign \A[13][13] [0] = 1'b1;
  assign \A[13][14] [0] = 1'b1;
  assign \A[13][15] [0] = 1'b1;
  assign \A[13][16] [4] = 1'b1;
  assign \A[13][16] [3] = 1'b1;
  assign \A[13][16] [2] = 1'b1;
  assign \A[13][16] [1] = 1'b1;
  assign \A[13][17] [4] = 1'b1;
  assign \A[13][17] [3] = 1'b1;
  assign \A[13][17] [2] = 1'b1;
  assign \A[13][17] [1] = 1'b1;
  assign \A[13][19] [4] = 1'b1;
  assign \A[13][19] [3] = 1'b1;
  assign \A[13][19] [2] = 1'b1;
  assign \A[13][19] [1] = 1'b1;
  assign \A[13][19] [0] = 1'b1;
  assign \A[13][20] [4] = 1'b1;
  assign \A[13][20] [3] = 1'b1;
  assign \A[13][20] [2] = 1'b1;
  assign \A[13][20] [1] = 1'b1;
  assign \A[13][21] [0] = 1'b1;
  assign \A[13][22] [0] = 1'b1;
  assign \A[13][26] [4] = 1'b1;
  assign \A[13][26] [3] = 1'b1;
  assign \A[13][26] [2] = 1'b1;
  assign \A[13][26] [1] = 1'b1;
  assign \A[13][27] [4] = 1'b1;
  assign \A[13][27] [3] = 1'b1;
  assign \A[13][27] [2] = 1'b1;
  assign \A[13][27] [1] = 1'b1;
  assign \A[13][27] [0] = 1'b1;
  assign \A[13][28] [1] = 1'b1;
  assign \A[13][30] [0] = 1'b1;
  assign \A[13][31] [0] = 1'b1;
  assign \A[13][32] [1] = 1'b1;
  assign \A[13][32] [0] = 1'b1;
  assign \A[13][33] [0] = 1'b1;
  assign \A[13][36] [4] = 1'b1;
  assign \A[13][36] [3] = 1'b1;
  assign \A[13][36] [2] = 1'b1;
  assign \A[13][37] [4] = 1'b1;
  assign \A[13][37] [3] = 1'b1;
  assign \A[13][37] [2] = 1'b1;
  assign \A[13][37] [1] = 1'b1;
  assign \A[13][37] [0] = 1'b1;
  assign \A[13][41] [0] = 1'b1;
  assign \A[13][42] [0] = 1'b1;
  assign \A[13][43] [0] = 1'b1;
  assign \A[13][44] [0] = 1'b1;
  assign \A[13][46] [4] = 1'b1;
  assign \A[13][46] [3] = 1'b1;
  assign \A[13][46] [2] = 1'b1;
  assign \A[13][46] [1] = 1'b1;
  assign \A[13][46] [0] = 1'b1;
  assign \A[13][48] [1] = 1'b1;
  assign \A[13][50] [0] = 1'b1;
  assign \A[13][51] [1] = 1'b1;
  assign \A[13][51] [0] = 1'b1;
  assign \A[13][52] [1] = 1'b1;
  assign \A[13][54] [4] = 1'b1;
  assign \A[13][54] [3] = 1'b1;
  assign \A[13][54] [2] = 1'b1;
  assign \A[13][54] [1] = 1'b1;
  assign \A[13][56] [4] = 1'b1;
  assign \A[13][56] [3] = 1'b1;
  assign \A[13][56] [2] = 1'b1;
  assign \A[13][56] [1] = 1'b1;
  assign \A[13][56] [0] = 1'b1;
  assign \A[13][57] [4] = 1'b1;
  assign \A[13][57] [3] = 1'b1;
  assign \A[13][57] [2] = 1'b1;
  assign \A[13][57] [1] = 1'b1;
  assign \A[13][57] [0] = 1'b1;
  assign \A[13][59] [4] = 1'b1;
  assign \A[13][59] [3] = 1'b1;
  assign \A[13][59] [2] = 1'b1;
  assign \A[13][59] [1] = 1'b1;
  assign \A[13][60] [4] = 1'b1;
  assign \A[13][60] [3] = 1'b1;
  assign \A[13][60] [2] = 1'b1;
  assign \A[13][60] [0] = 1'b1;
  assign \A[13][61] [0] = 1'b1;
  assign \A[13][62] [0] = 1'b1;
  assign \A[13][63] [1] = 1'b1;
  assign \A[13][63] [0] = 1'b1;
  assign \A[13][64] [0] = 1'b1;
  assign \A[13][65] [0] = 1'b1;
  assign \A[13][67] [4] = 1'b1;
  assign \A[13][67] [3] = 1'b1;
  assign \A[13][67] [2] = 1'b1;
  assign \A[13][67] [1] = 1'b1;
  assign \A[13][68] [0] = 1'b1;
  assign \A[13][69] [0] = 1'b1;
  assign \A[13][70] [4] = 1'b1;
  assign \A[13][70] [3] = 1'b1;
  assign \A[13][70] [2] = 1'b1;
  assign \A[13][70] [0] = 1'b1;
  assign \A[13][72] [1] = 1'b1;
  assign \A[13][72] [0] = 1'b1;
  assign \A[13][73] [4] = 1'b1;
  assign \A[13][73] [3] = 1'b1;
  assign \A[13][73] [2] = 1'b1;
  assign \A[13][73] [1] = 1'b1;
  assign \A[13][73] [0] = 1'b1;
  assign \A[13][75] [0] = 1'b1;
  assign \A[13][77] [0] = 1'b1;
  assign \A[13][79] [4] = 1'b1;
  assign \A[13][79] [3] = 1'b1;
  assign \A[13][79] [2] = 1'b1;
  assign \A[13][79] [1] = 1'b1;
  assign \A[13][81] [4] = 1'b1;
  assign \A[13][81] [3] = 1'b1;
  assign \A[13][81] [2] = 1'b1;
  assign \A[13][81] [1] = 1'b1;
  assign \A[13][81] [0] = 1'b1;
  assign \A[13][82] [1] = 1'b1;
  assign \A[13][82] [0] = 1'b1;
  assign \A[13][83] [0] = 1'b1;
  assign \A[13][84] [4] = 1'b1;
  assign \A[13][84] [3] = 1'b1;
  assign \A[13][84] [2] = 1'b1;
  assign \A[13][84] [1] = 1'b1;
  assign \A[13][85] [4] = 1'b1;
  assign \A[13][85] [3] = 1'b1;
  assign \A[13][85] [2] = 1'b1;
  assign \A[13][85] [1] = 1'b1;
  assign \A[13][87] [4] = 1'b1;
  assign \A[13][87] [3] = 1'b1;
  assign \A[13][87] [2] = 1'b1;
  assign \A[13][87] [1] = 1'b1;
  assign \A[13][88] [0] = 1'b1;
  assign \A[13][89] [0] = 1'b1;
  assign \A[13][90] [4] = 1'b1;
  assign \A[13][90] [3] = 1'b1;
  assign \A[13][90] [2] = 1'b1;
  assign \A[13][90] [1] = 1'b1;
  assign \A[13][91] [4] = 1'b1;
  assign \A[13][91] [3] = 1'b1;
  assign \A[13][91] [2] = 1'b1;
  assign \A[13][91] [1] = 1'b1;
  assign \A[13][91] [0] = 1'b1;
  assign \A[13][92] [1] = 1'b1;
  assign \A[13][93] [1] = 1'b1;
  assign \A[13][94] [0] = 1'b1;
  assign \A[13][95] [0] = 1'b1;
  assign \A[13][97] [4] = 1'b1;
  assign \A[13][97] [3] = 1'b1;
  assign \A[13][97] [2] = 1'b1;
  assign \A[13][97] [0] = 1'b1;
  assign \A[13][98] [0] = 1'b1;
  assign \A[13][99] [1] = 1'b1;
  assign \A[13][101] [0] = 1'b1;
  assign \A[13][102] [0] = 1'b1;
  assign \A[13][103] [4] = 1'b1;
  assign \A[13][103] [3] = 1'b1;
  assign \A[13][103] [2] = 1'b1;
  assign \A[13][103] [1] = 1'b1;
  assign \A[13][104] [4] = 1'b1;
  assign \A[13][104] [3] = 1'b1;
  assign \A[13][104] [2] = 1'b1;
  assign \A[13][104] [1] = 1'b1;
  assign \A[13][104] [0] = 1'b1;
  assign \A[13][106] [4] = 1'b1;
  assign \A[13][106] [3] = 1'b1;
  assign \A[13][106] [2] = 1'b1;
  assign \A[13][106] [1] = 1'b1;
  assign \A[13][106] [0] = 1'b1;
  assign \A[13][107] [0] = 1'b1;
  assign \A[13][108] [0] = 1'b1;
  assign \A[13][109] [4] = 1'b1;
  assign \A[13][109] [3] = 1'b1;
  assign \A[13][109] [2] = 1'b1;
  assign \A[13][109] [1] = 1'b1;
  assign \A[13][109] [0] = 1'b1;
  assign \A[13][112] [0] = 1'b1;
  assign \A[13][113] [4] = 1'b1;
  assign \A[13][113] [3] = 1'b1;
  assign \A[13][113] [2] = 1'b1;
  assign \A[13][113] [1] = 1'b1;
  assign \A[13][113] [0] = 1'b1;
  assign \A[13][114] [4] = 1'b1;
  assign \A[13][114] [3] = 1'b1;
  assign \A[13][114] [2] = 1'b1;
  assign \A[13][114] [1] = 1'b1;
  assign \A[13][114] [0] = 1'b1;
  assign \A[13][117] [4] = 1'b1;
  assign \A[13][117] [3] = 1'b1;
  assign \A[13][117] [2] = 1'b1;
  assign \A[13][117] [1] = 1'b1;
  assign \A[13][117] [0] = 1'b1;
  assign \A[13][118] [4] = 1'b1;
  assign \A[13][118] [3] = 1'b1;
  assign \A[13][118] [2] = 1'b1;
  assign \A[13][118] [1] = 1'b1;
  assign \A[13][118] [0] = 1'b1;
  assign \A[13][119] [0] = 1'b1;
  assign \A[13][120] [4] = 1'b1;
  assign \A[13][120] [3] = 1'b1;
  assign \A[13][120] [2] = 1'b1;
  assign \A[13][120] [1] = 1'b1;
  assign \A[13][120] [0] = 1'b1;
  assign \A[13][121] [0] = 1'b1;
  assign \A[13][123] [0] = 1'b1;
  assign \A[13][125] [0] = 1'b1;
  assign \A[13][126] [4] = 1'b1;
  assign \A[13][126] [3] = 1'b1;
  assign \A[13][126] [2] = 1'b1;
  assign \A[13][126] [1] = 1'b1;
  assign \A[13][126] [0] = 1'b1;
  assign \A[13][127] [0] = 1'b1;
  assign \A[13][128] [1] = 1'b1;
  assign \A[13][130] [4] = 1'b1;
  assign \A[13][130] [3] = 1'b1;
  assign \A[13][130] [2] = 1'b1;
  assign \A[13][130] [1] = 1'b1;
  assign \A[13][131] [1] = 1'b1;
  assign \A[13][133] [0] = 1'b1;
  assign \A[13][134] [4] = 1'b1;
  assign \A[13][134] [3] = 1'b1;
  assign \A[13][134] [2] = 1'b1;
  assign \A[13][134] [1] = 1'b1;
  assign \A[13][135] [4] = 1'b1;
  assign \A[13][135] [3] = 1'b1;
  assign \A[13][135] [2] = 1'b1;
  assign \A[13][135] [1] = 1'b1;
  assign \A[13][135] [0] = 1'b1;
  assign \A[13][137] [4] = 1'b1;
  assign \A[13][137] [3] = 1'b1;
  assign \A[13][137] [2] = 1'b1;
  assign \A[13][137] [1] = 1'b1;
  assign \A[13][137] [0] = 1'b1;
  assign \A[13][139] [4] = 1'b1;
  assign \A[13][139] [3] = 1'b1;
  assign \A[13][139] [2] = 1'b1;
  assign \A[13][139] [1] = 1'b1;
  assign \A[13][140] [4] = 1'b1;
  assign \A[13][140] [3] = 1'b1;
  assign \A[13][140] [2] = 1'b1;
  assign \A[13][140] [1] = 1'b1;
  assign \A[13][140] [0] = 1'b1;
  assign \A[13][141] [4] = 1'b1;
  assign \A[13][141] [3] = 1'b1;
  assign \A[13][141] [2] = 1'b1;
  assign \A[13][141] [1] = 1'b1;
  assign \A[13][143] [4] = 1'b1;
  assign \A[13][143] [3] = 1'b1;
  assign \A[13][143] [1] = 1'b1;
  assign \A[13][143] [0] = 1'b1;
  assign \A[13][144] [0] = 1'b1;
  assign \A[13][146] [4] = 1'b1;
  assign \A[13][146] [3] = 1'b1;
  assign \A[13][146] [2] = 1'b1;
  assign \A[13][146] [1] = 1'b1;
  assign \A[13][146] [0] = 1'b1;
  assign \A[13][148] [4] = 1'b1;
  assign \A[13][148] [3] = 1'b1;
  assign \A[13][148] [2] = 1'b1;
  assign \A[13][148] [1] = 1'b1;
  assign \A[13][150] [1] = 1'b1;
  assign \A[13][152] [1] = 1'b1;
  assign \A[13][153] [1] = 1'b1;
  assign \A[13][156] [0] = 1'b1;
  assign \A[13][157] [1] = 1'b1;
  assign \A[13][158] [0] = 1'b1;
  assign \A[13][159] [4] = 1'b1;
  assign \A[13][159] [3] = 1'b1;
  assign \A[13][159] [2] = 1'b1;
  assign \A[13][159] [1] = 1'b1;
  assign \A[13][160] [0] = 1'b1;
  assign \A[13][161] [1] = 1'b1;
  assign \A[13][162] [4] = 1'b1;
  assign \A[13][162] [3] = 1'b1;
  assign \A[13][162] [2] = 1'b1;
  assign \A[13][162] [1] = 1'b1;
  assign \A[13][162] [0] = 1'b1;
  assign \A[13][165] [0] = 1'b1;
  assign \A[13][166] [4] = 1'b1;
  assign \A[13][166] [3] = 1'b1;
  assign \A[13][166] [2] = 1'b1;
  assign \A[13][166] [1] = 1'b1;
  assign \A[13][166] [0] = 1'b1;
  assign \A[13][167] [1] = 1'b1;
  assign \A[13][167] [0] = 1'b1;
  assign \A[13][168] [4] = 1'b1;
  assign \A[13][168] [3] = 1'b1;
  assign \A[13][168] [2] = 1'b1;
  assign \A[13][168] [1] = 1'b1;
  assign \A[13][168] [0] = 1'b1;
  assign \A[13][169] [4] = 1'b1;
  assign \A[13][169] [3] = 1'b1;
  assign \A[13][169] [2] = 1'b1;
  assign \A[13][169] [1] = 1'b1;
  assign \A[13][169] [0] = 1'b1;
  assign \A[13][171] [4] = 1'b1;
  assign \A[13][171] [3] = 1'b1;
  assign \A[13][171] [2] = 1'b1;
  assign \A[13][171] [1] = 1'b1;
  assign \A[13][171] [0] = 1'b1;
  assign \A[13][172] [4] = 1'b1;
  assign \A[13][172] [3] = 1'b1;
  assign \A[13][172] [2] = 1'b1;
  assign \A[13][172] [1] = 1'b1;
  assign \A[13][173] [0] = 1'b1;
  assign \A[13][174] [4] = 1'b1;
  assign \A[13][174] [3] = 1'b1;
  assign \A[13][174] [2] = 1'b1;
  assign \A[13][174] [1] = 1'b1;
  assign \A[13][174] [0] = 1'b1;
  assign \A[13][175] [1] = 1'b1;
  assign \A[13][176] [1] = 1'b1;
  assign \A[13][179] [0] = 1'b1;
  assign \A[13][180] [0] = 1'b1;
  assign \A[13][181] [1] = 1'b1;
  assign \A[13][182] [0] = 1'b1;
  assign \A[13][184] [1] = 1'b1;
  assign \A[13][186] [4] = 1'b1;
  assign \A[13][186] [3] = 1'b1;
  assign \A[13][186] [2] = 1'b1;
  assign \A[13][186] [1] = 1'b1;
  assign \A[13][186] [0] = 1'b1;
  assign \A[13][187] [4] = 1'b1;
  assign \A[13][187] [3] = 1'b1;
  assign \A[13][187] [2] = 1'b1;
  assign \A[13][187] [1] = 1'b1;
  assign \A[13][189] [4] = 1'b1;
  assign \A[13][189] [3] = 1'b1;
  assign \A[13][189] [2] = 1'b1;
  assign \A[13][189] [1] = 1'b1;
  assign \A[13][189] [0] = 1'b1;
  assign \A[13][191] [1] = 1'b1;
  assign \A[13][192] [1] = 1'b1;
  assign \A[13][192] [0] = 1'b1;
  assign \A[13][193] [4] = 1'b1;
  assign \A[13][193] [3] = 1'b1;
  assign \A[13][193] [2] = 1'b1;
  assign \A[13][193] [1] = 1'b1;
  assign \A[13][194] [0] = 1'b1;
  assign \A[13][195] [1] = 1'b1;
  assign \A[13][198] [0] = 1'b1;
  assign \A[13][199] [0] = 1'b1;
  assign \A[13][201] [0] = 1'b1;
  assign \A[13][202] [0] = 1'b1;
  assign \A[13][203] [4] = 1'b1;
  assign \A[13][203] [3] = 1'b1;
  assign \A[13][203] [2] = 1'b1;
  assign \A[13][203] [1] = 1'b1;
  assign \A[13][203] [0] = 1'b1;
  assign \A[13][204] [0] = 1'b1;
  assign \A[13][205] [1] = 1'b1;
  assign \A[13][205] [0] = 1'b1;
  assign \A[13][207] [4] = 1'b1;
  assign \A[13][207] [3] = 1'b1;
  assign \A[13][207] [2] = 1'b1;
  assign \A[13][207] [1] = 1'b1;
  assign \A[13][207] [0] = 1'b1;
  assign \A[13][208] [1] = 1'b1;
  assign \A[13][210] [1] = 1'b1;
  assign \A[13][211] [4] = 1'b1;
  assign \A[13][211] [3] = 1'b1;
  assign \A[13][211] [2] = 1'b1;
  assign \A[13][211] [1] = 1'b1;
  assign \A[13][211] [0] = 1'b1;
  assign \A[13][213] [1] = 1'b1;
  assign \A[13][215] [4] = 1'b1;
  assign \A[13][215] [3] = 1'b1;
  assign \A[13][215] [2] = 1'b1;
  assign \A[13][215] [1] = 1'b1;
  assign \A[13][215] [0] = 1'b1;
  assign \A[13][216] [4] = 1'b1;
  assign \A[13][216] [3] = 1'b1;
  assign \A[13][216] [2] = 1'b1;
  assign \A[13][216] [1] = 1'b1;
  assign \A[13][216] [0] = 1'b1;
  assign \A[13][217] [1] = 1'b1;
  assign \A[13][217] [0] = 1'b1;
  assign \A[13][220] [1] = 1'b1;
  assign \A[13][220] [0] = 1'b1;
  assign \A[13][222] [4] = 1'b1;
  assign \A[13][222] [3] = 1'b1;
  assign \A[13][222] [2] = 1'b1;
  assign \A[13][222] [1] = 1'b1;
  assign \A[13][222] [0] = 1'b1;
  assign \A[13][223] [4] = 1'b1;
  assign \A[13][223] [3] = 1'b1;
  assign \A[13][223] [2] = 1'b1;
  assign \A[13][223] [1] = 1'b1;
  assign \A[13][223] [0] = 1'b1;
  assign \A[13][224] [1] = 1'b1;
  assign \A[13][225] [4] = 1'b1;
  assign \A[13][225] [3] = 1'b1;
  assign \A[13][225] [2] = 1'b1;
  assign \A[13][225] [1] = 1'b1;
  assign \A[13][225] [0] = 1'b1;
  assign \A[13][226] [4] = 1'b1;
  assign \A[13][226] [3] = 1'b1;
  assign \A[13][226] [2] = 1'b1;
  assign \A[13][226] [1] = 1'b1;
  assign \A[13][228] [4] = 1'b1;
  assign \A[13][228] [3] = 1'b1;
  assign \A[13][228] [2] = 1'b1;
  assign \A[13][228] [1] = 1'b1;
  assign \A[13][228] [0] = 1'b1;
  assign \A[13][229] [1] = 1'b1;
  assign \A[13][230] [1] = 1'b1;
  assign \A[13][231] [1] = 1'b1;
  assign \A[13][231] [0] = 1'b1;
  assign \A[13][233] [1] = 1'b1;
  assign \A[13][233] [0] = 1'b1;
  assign \A[13][235] [0] = 1'b1;
  assign \A[13][236] [4] = 1'b1;
  assign \A[13][236] [3] = 1'b1;
  assign \A[13][236] [2] = 1'b1;
  assign \A[13][236] [1] = 1'b1;
  assign \A[13][236] [0] = 1'b1;
  assign \A[13][237] [4] = 1'b1;
  assign \A[13][237] [3] = 1'b1;
  assign \A[13][237] [2] = 1'b1;
  assign \A[13][237] [1] = 1'b1;
  assign \A[13][237] [0] = 1'b1;
  assign \A[13][239] [4] = 1'b1;
  assign \A[13][239] [3] = 1'b1;
  assign \A[13][239] [2] = 1'b1;
  assign \A[13][239] [1] = 1'b1;
  assign \A[13][241] [4] = 1'b1;
  assign \A[13][241] [3] = 1'b1;
  assign \A[13][241] [2] = 1'b1;
  assign \A[13][241] [1] = 1'b1;
  assign \A[13][241] [0] = 1'b1;
  assign \A[13][242] [4] = 1'b1;
  assign \A[13][242] [3] = 1'b1;
  assign \A[13][242] [2] = 1'b1;
  assign \A[13][242] [1] = 1'b1;
  assign \A[13][244] [1] = 1'b1;
  assign \A[13][245] [0] = 1'b1;
  assign \A[13][246] [1] = 1'b1;
  assign \A[13][247] [4] = 1'b1;
  assign \A[13][247] [3] = 1'b1;
  assign \A[13][247] [2] = 1'b1;
  assign \A[13][247] [1] = 1'b1;
  assign \A[13][248] [0] = 1'b1;
  assign \A[13][249] [4] = 1'b1;
  assign \A[13][249] [3] = 1'b1;
  assign \A[13][249] [2] = 1'b1;
  assign \A[13][249] [1] = 1'b1;
  assign \A[13][249] [0] = 1'b1;
  assign \A[13][250] [0] = 1'b1;
  assign \A[13][251] [0] = 1'b1;
  assign \A[13][252] [4] = 1'b1;
  assign \A[13][252] [3] = 1'b1;
  assign \A[13][252] [2] = 1'b1;
  assign \A[13][252] [1] = 1'b1;
  assign \A[13][253] [4] = 1'b1;
  assign \A[13][253] [3] = 1'b1;
  assign \A[13][253] [2] = 1'b1;
  assign \A[13][253] [1] = 1'b1;
  assign \A[13][253] [0] = 1'b1;
  assign \A[13][254] [0] = 1'b1;
  assign \A[14][0] [0] = 1'b1;
  assign \A[14][1] [4] = 1'b1;
  assign \A[14][1] [3] = 1'b1;
  assign \A[14][1] [2] = 1'b1;
  assign \A[14][3] [4] = 1'b1;
  assign \A[14][3] [3] = 1'b1;
  assign \A[14][3] [2] = 1'b1;
  assign \A[14][3] [1] = 1'b1;
  assign \A[14][3] [0] = 1'b1;
  assign \A[14][4] [4] = 1'b1;
  assign \A[14][4] [3] = 1'b1;
  assign \A[14][4] [2] = 1'b1;
  assign \A[14][4] [1] = 1'b1;
  assign \A[14][4] [0] = 1'b1;
  assign \A[14][5] [1] = 1'b1;
  assign \A[14][6] [0] = 1'b1;
  assign \A[14][7] [1] = 1'b1;
  assign \A[14][8] [0] = 1'b1;
  assign \A[14][10] [4] = 1'b1;
  assign \A[14][10] [3] = 1'b1;
  assign \A[14][10] [2] = 1'b1;
  assign \A[14][10] [1] = 1'b1;
  assign \A[14][10] [0] = 1'b1;
  assign \A[14][11] [4] = 1'b1;
  assign \A[14][11] [3] = 1'b1;
  assign \A[14][11] [2] = 1'b1;
  assign \A[14][11] [1] = 1'b1;
  assign \A[14][11] [0] = 1'b1;
  assign \A[14][12] [4] = 1'b1;
  assign \A[14][12] [3] = 1'b1;
  assign \A[14][12] [2] = 1'b1;
  assign \A[14][12] [1] = 1'b1;
  assign \A[14][12] [0] = 1'b1;
  assign \A[14][15] [4] = 1'b1;
  assign \A[14][15] [3] = 1'b1;
  assign \A[14][15] [2] = 1'b1;
  assign \A[14][15] [0] = 1'b1;
  assign \A[14][17] [1] = 1'b1;
  assign \A[14][17] [0] = 1'b1;
  assign \A[14][18] [0] = 1'b1;
  assign \A[14][19] [4] = 1'b1;
  assign \A[14][19] [3] = 1'b1;
  assign \A[14][19] [2] = 1'b1;
  assign \A[14][19] [1] = 1'b1;
  assign \A[14][19] [0] = 1'b1;
  assign \A[14][21] [4] = 1'b1;
  assign \A[14][21] [3] = 1'b1;
  assign \A[14][21] [2] = 1'b1;
  assign \A[14][21] [0] = 1'b1;
  assign \A[14][23] [0] = 1'b1;
  assign \A[14][24] [1] = 1'b1;
  assign \A[14][24] [0] = 1'b1;
  assign \A[14][27] [1] = 1'b1;
  assign \A[14][30] [4] = 1'b1;
  assign \A[14][30] [3] = 1'b1;
  assign \A[14][30] [2] = 1'b1;
  assign \A[14][30] [1] = 1'b1;
  assign \A[14][32] [4] = 1'b1;
  assign \A[14][32] [3] = 1'b1;
  assign \A[14][32] [2] = 1'b1;
  assign \A[14][32] [1] = 1'b1;
  assign \A[14][32] [0] = 1'b1;
  assign \A[14][33] [2] = 1'b1;
  assign \A[14][34] [4] = 1'b1;
  assign \A[14][34] [3] = 1'b1;
  assign \A[14][34] [2] = 1'b1;
  assign \A[14][34] [1] = 1'b1;
  assign \A[14][34] [0] = 1'b1;
  assign \A[14][35] [4] = 1'b1;
  assign \A[14][35] [3] = 1'b1;
  assign \A[14][35] [2] = 1'b1;
  assign \A[14][35] [1] = 1'b1;
  assign \A[14][36] [4] = 1'b1;
  assign \A[14][36] [3] = 1'b1;
  assign \A[14][36] [2] = 1'b1;
  assign \A[14][36] [1] = 1'b1;
  assign \A[14][36] [0] = 1'b1;
  assign \A[14][37] [1] = 1'b1;
  assign \A[14][38] [4] = 1'b1;
  assign \A[14][38] [3] = 1'b1;
  assign \A[14][38] [2] = 1'b1;
  assign \A[14][38] [1] = 1'b1;
  assign \A[14][38] [0] = 1'b1;
  assign \A[14][39] [1] = 1'b1;
  assign \A[14][40] [4] = 1'b1;
  assign \A[14][40] [3] = 1'b1;
  assign \A[14][40] [2] = 1'b1;
  assign \A[14][40] [1] = 1'b1;
  assign \A[14][40] [0] = 1'b1;
  assign \A[14][42] [4] = 1'b1;
  assign \A[14][42] [3] = 1'b1;
  assign \A[14][42] [2] = 1'b1;
  assign \A[14][42] [1] = 1'b1;
  assign \A[14][44] [4] = 1'b1;
  assign \A[14][44] [3] = 1'b1;
  assign \A[14][44] [2] = 1'b1;
  assign \A[14][44] [1] = 1'b1;
  assign \A[14][45] [4] = 1'b1;
  assign \A[14][45] [3] = 1'b1;
  assign \A[14][45] [2] = 1'b1;
  assign \A[14][45] [0] = 1'b1;
  assign \A[14][46] [4] = 1'b1;
  assign \A[14][46] [3] = 1'b1;
  assign \A[14][46] [2] = 1'b1;
  assign \A[14][46] [1] = 1'b1;
  assign \A[14][47] [0] = 1'b1;
  assign \A[14][48] [0] = 1'b1;
  assign \A[14][49] [1] = 1'b1;
  assign \A[14][49] [0] = 1'b1;
  assign \A[14][50] [1] = 1'b1;
  assign \A[14][50] [0] = 1'b1;
  assign \A[14][51] [4] = 1'b1;
  assign \A[14][51] [3] = 1'b1;
  assign \A[14][51] [2] = 1'b1;
  assign \A[14][51] [1] = 1'b1;
  assign \A[14][52] [0] = 1'b1;
  assign \A[14][54] [0] = 1'b1;
  assign \A[14][55] [4] = 1'b1;
  assign \A[14][55] [3] = 1'b1;
  assign \A[14][55] [2] = 1'b1;
  assign \A[14][55] [0] = 1'b1;
  assign \A[14][56] [0] = 1'b1;
  assign \A[14][57] [4] = 1'b1;
  assign \A[14][57] [3] = 1'b1;
  assign \A[14][57] [2] = 1'b1;
  assign \A[14][57] [1] = 1'b1;
  assign \A[14][59] [4] = 1'b1;
  assign \A[14][59] [3] = 1'b1;
  assign \A[14][59] [2] = 1'b1;
  assign \A[14][59] [1] = 1'b1;
  assign \A[14][59] [0] = 1'b1;
  assign \A[14][60] [4] = 1'b1;
  assign \A[14][60] [3] = 1'b1;
  assign \A[14][60] [2] = 1'b1;
  assign \A[14][60] [1] = 1'b1;
  assign \A[14][60] [0] = 1'b1;
  assign \A[14][61] [4] = 1'b1;
  assign \A[14][61] [3] = 1'b1;
  assign \A[14][61] [2] = 1'b1;
  assign \A[14][61] [1] = 1'b1;
  assign \A[14][61] [0] = 1'b1;
  assign \A[14][62] [0] = 1'b1;
  assign \A[14][63] [1] = 1'b1;
  assign \A[14][64] [0] = 1'b1;
  assign \A[14][65] [1] = 1'b1;
  assign \A[14][66] [0] = 1'b1;
  assign \A[14][68] [0] = 1'b1;
  assign \A[14][69] [0] = 1'b1;
  assign \A[14][72] [4] = 1'b1;
  assign \A[14][72] [3] = 1'b1;
  assign \A[14][72] [2] = 1'b1;
  assign \A[14][72] [1] = 1'b1;
  assign \A[14][72] [0] = 1'b1;
  assign \A[14][73] [0] = 1'b1;
  assign \A[14][74] [4] = 1'b1;
  assign \A[14][74] [3] = 1'b1;
  assign \A[14][74] [2] = 1'b1;
  assign \A[14][74] [1] = 1'b1;
  assign \A[14][75] [1] = 1'b1;
  assign \A[14][76] [4] = 1'b1;
  assign \A[14][76] [3] = 1'b1;
  assign \A[14][76] [2] = 1'b1;
  assign \A[14][76] [1] = 1'b1;
  assign \A[14][76] [0] = 1'b1;
  assign \A[14][77] [4] = 1'b1;
  assign \A[14][77] [3] = 1'b1;
  assign \A[14][77] [2] = 1'b1;
  assign \A[14][77] [1] = 1'b1;
  assign \A[14][79] [4] = 1'b1;
  assign \A[14][79] [3] = 1'b1;
  assign \A[14][79] [2] = 1'b1;
  assign \A[14][79] [1] = 1'b1;
  assign \A[14][79] [0] = 1'b1;
  assign \A[14][80] [4] = 1'b1;
  assign \A[14][80] [3] = 1'b1;
  assign \A[14][80] [2] = 1'b1;
  assign \A[14][80] [1] = 1'b1;
  assign \A[14][82] [2] = 1'b1;
  assign \A[14][86] [2] = 1'b1;
  assign \A[14][87] [4] = 1'b1;
  assign \A[14][87] [3] = 1'b1;
  assign \A[14][87] [2] = 1'b1;
  assign \A[14][87] [0] = 1'b1;
  assign \A[14][88] [0] = 1'b1;
  assign \A[14][94] [0] = 1'b1;
  assign \A[14][95] [4] = 1'b1;
  assign \A[14][95] [3] = 1'b1;
  assign \A[14][95] [2] = 1'b1;
  assign \A[14][95] [1] = 1'b1;
  assign \A[14][95] [0] = 1'b1;
  assign \A[14][96] [4] = 1'b1;
  assign \A[14][96] [3] = 1'b1;
  assign \A[14][96] [2] = 1'b1;
  assign \A[14][96] [1] = 1'b1;
  assign \A[14][96] [0] = 1'b1;
  assign \A[14][98] [0] = 1'b1;
  assign \A[14][99] [4] = 1'b1;
  assign \A[14][99] [3] = 1'b1;
  assign \A[14][99] [2] = 1'b1;
  assign \A[14][99] [0] = 1'b1;
  assign \A[14][101] [4] = 1'b1;
  assign \A[14][101] [3] = 1'b1;
  assign \A[14][101] [2] = 1'b1;
  assign \A[14][101] [1] = 1'b1;
  assign \A[14][101] [0] = 1'b1;
  assign \A[14][102] [1] = 1'b1;
  assign \A[14][103] [4] = 1'b1;
  assign \A[14][103] [3] = 1'b1;
  assign \A[14][103] [2] = 1'b1;
  assign \A[14][103] [0] = 1'b1;
  assign \A[14][105] [4] = 1'b1;
  assign \A[14][105] [3] = 1'b1;
  assign \A[14][105] [2] = 1'b1;
  assign \A[14][105] [1] = 1'b1;
  assign \A[14][105] [0] = 1'b1;
  assign \A[14][106] [4] = 1'b1;
  assign \A[14][106] [3] = 1'b1;
  assign \A[14][106] [2] = 1'b1;
  assign \A[14][106] [1] = 1'b1;
  assign \A[14][106] [0] = 1'b1;
  assign \A[14][107] [0] = 1'b1;
  assign \A[14][109] [0] = 1'b1;
  assign \A[14][110] [0] = 1'b1;
  assign \A[14][111] [4] = 1'b1;
  assign \A[14][111] [3] = 1'b1;
  assign \A[14][111] [2] = 1'b1;
  assign \A[14][111] [1] = 1'b1;
  assign \A[14][112] [4] = 1'b1;
  assign \A[14][112] [3] = 1'b1;
  assign \A[14][112] [2] = 1'b1;
  assign \A[14][112] [1] = 1'b1;
  assign \A[14][113] [0] = 1'b1;
  assign \A[14][114] [4] = 1'b1;
  assign \A[14][114] [3] = 1'b1;
  assign \A[14][114] [2] = 1'b1;
  assign \A[14][114] [0] = 1'b1;
  assign \A[14][115] [0] = 1'b1;
  assign \A[14][116] [4] = 1'b1;
  assign \A[14][116] [3] = 1'b1;
  assign \A[14][116] [2] = 1'b1;
  assign \A[14][116] [1] = 1'b1;
  assign \A[14][116] [0] = 1'b1;
  assign \A[14][117] [0] = 1'b1;
  assign \A[14][118] [4] = 1'b1;
  assign \A[14][118] [3] = 1'b1;
  assign \A[14][118] [2] = 1'b1;
  assign \A[14][118] [1] = 1'b1;
  assign \A[14][118] [0] = 1'b1;
  assign \A[14][123] [0] = 1'b1;
  assign \A[14][124] [0] = 1'b1;
  assign \A[14][125] [4] = 1'b1;
  assign \A[14][125] [3] = 1'b1;
  assign \A[14][125] [2] = 1'b1;
  assign \A[14][125] [1] = 1'b1;
  assign \A[14][126] [1] = 1'b1;
  assign \A[14][128] [0] = 1'b1;
  assign \A[14][129] [4] = 1'b1;
  assign \A[14][129] [3] = 1'b1;
  assign \A[14][129] [2] = 1'b1;
  assign \A[14][129] [1] = 1'b1;
  assign \A[14][129] [0] = 1'b1;
  assign \A[14][131] [4] = 1'b1;
  assign \A[14][131] [3] = 1'b1;
  assign \A[14][131] [2] = 1'b1;
  assign \A[14][131] [0] = 1'b1;
  assign \A[14][132] [0] = 1'b1;
  assign \A[14][133] [4] = 1'b1;
  assign \A[14][133] [3] = 1'b1;
  assign \A[14][133] [2] = 1'b1;
  assign \A[14][133] [1] = 1'b1;
  assign \A[14][133] [0] = 1'b1;
  assign \A[14][134] [4] = 1'b1;
  assign \A[14][134] [3] = 1'b1;
  assign \A[14][134] [2] = 1'b1;
  assign \A[14][134] [1] = 1'b1;
  assign \A[14][134] [0] = 1'b1;
  assign \A[14][135] [4] = 1'b1;
  assign \A[14][135] [3] = 1'b1;
  assign \A[14][135] [2] = 1'b1;
  assign \A[14][135] [1] = 1'b1;
  assign \A[14][135] [0] = 1'b1;
  assign \A[14][137] [4] = 1'b1;
  assign \A[14][137] [3] = 1'b1;
  assign \A[14][137] [2] = 1'b1;
  assign \A[14][137] [1] = 1'b1;
  assign \A[14][138] [2] = 1'b1;
  assign \A[14][139] [0] = 1'b1;
  assign \A[14][141] [4] = 1'b1;
  assign \A[14][141] [3] = 1'b1;
  assign \A[14][141] [2] = 1'b1;
  assign \A[14][141] [1] = 1'b1;
  assign \A[14][141] [0] = 1'b1;
  assign \A[14][142] [4] = 1'b1;
  assign \A[14][142] [3] = 1'b1;
  assign \A[14][142] [2] = 1'b1;
  assign \A[14][142] [1] = 1'b1;
  assign \A[14][142] [0] = 1'b1;
  assign \A[14][145] [4] = 1'b1;
  assign \A[14][145] [3] = 1'b1;
  assign \A[14][145] [2] = 1'b1;
  assign \A[14][145] [1] = 1'b1;
  assign \A[14][145] [0] = 1'b1;
  assign \A[14][146] [4] = 1'b1;
  assign \A[14][146] [3] = 1'b1;
  assign \A[14][146] [2] = 1'b1;
  assign \A[14][146] [1] = 1'b1;
  assign \A[14][146] [0] = 1'b1;
  assign \A[14][147] [4] = 1'b1;
  assign \A[14][147] [3] = 1'b1;
  assign \A[14][147] [2] = 1'b1;
  assign \A[14][147] [1] = 1'b1;
  assign \A[14][147] [0] = 1'b1;
  assign \A[14][149] [4] = 1'b1;
  assign \A[14][149] [3] = 1'b1;
  assign \A[14][149] [2] = 1'b1;
  assign \A[14][149] [1] = 1'b1;
  assign \A[14][149] [0] = 1'b1;
  assign \A[14][150] [4] = 1'b1;
  assign \A[14][150] [3] = 1'b1;
  assign \A[14][150] [2] = 1'b1;
  assign \A[14][150] [1] = 1'b1;
  assign \A[14][150] [0] = 1'b1;
  assign \A[14][151] [4] = 1'b1;
  assign \A[14][151] [3] = 1'b1;
  assign \A[14][151] [2] = 1'b1;
  assign \A[14][151] [1] = 1'b1;
  assign \A[14][151] [0] = 1'b1;
  assign \A[14][153] [0] = 1'b1;
  assign \A[14][154] [4] = 1'b1;
  assign \A[14][154] [3] = 1'b1;
  assign \A[14][154] [2] = 1'b1;
  assign \A[14][154] [1] = 1'b1;
  assign \A[14][154] [0] = 1'b1;
  assign \A[14][155] [1] = 1'b1;
  assign \A[14][156] [0] = 1'b1;
  assign \A[14][157] [4] = 1'b1;
  assign \A[14][157] [3] = 1'b1;
  assign \A[14][157] [2] = 1'b1;
  assign \A[14][157] [1] = 1'b1;
  assign \A[14][159] [4] = 1'b1;
  assign \A[14][159] [3] = 1'b1;
  assign \A[14][159] [2] = 1'b1;
  assign \A[14][159] [1] = 1'b1;
  assign \A[14][159] [0] = 1'b1;
  assign \A[14][160] [0] = 1'b1;
  assign \A[14][161] [1] = 1'b1;
  assign \A[14][164] [4] = 1'b1;
  assign \A[14][164] [3] = 1'b1;
  assign \A[14][164] [2] = 1'b1;
  assign \A[14][164] [1] = 1'b1;
  assign \A[14][165] [0] = 1'b1;
  assign \A[14][169] [0] = 1'b1;
  assign \A[14][171] [4] = 1'b1;
  assign \A[14][171] [3] = 1'b1;
  assign \A[14][171] [2] = 1'b1;
  assign \A[14][171] [1] = 1'b1;
  assign \A[14][171] [0] = 1'b1;
  assign \A[14][173] [1] = 1'b1;
  assign \A[14][173] [0] = 1'b1;
  assign \A[14][174] [0] = 1'b1;
  assign \A[14][175] [0] = 1'b1;
  assign \A[14][177] [0] = 1'b1;
  assign \A[14][178] [4] = 1'b1;
  assign \A[14][178] [3] = 1'b1;
  assign \A[14][178] [2] = 1'b1;
  assign \A[14][178] [1] = 1'b1;
  assign \A[14][178] [0] = 1'b1;
  assign \A[14][180] [1] = 1'b1;
  assign \A[14][181] [0] = 1'b1;
  assign \A[14][182] [4] = 1'b1;
  assign \A[14][182] [3] = 1'b1;
  assign \A[14][182] [2] = 1'b1;
  assign \A[14][182] [1] = 1'b1;
  assign \A[14][182] [0] = 1'b1;
  assign \A[14][183] [4] = 1'b1;
  assign \A[14][183] [3] = 1'b1;
  assign \A[14][183] [2] = 1'b1;
  assign \A[14][185] [4] = 1'b1;
  assign \A[14][185] [3] = 1'b1;
  assign \A[14][185] [2] = 1'b1;
  assign \A[14][185] [1] = 1'b1;
  assign \A[14][185] [0] = 1'b1;
  assign \A[14][187] [1] = 1'b1;
  assign \A[14][189] [4] = 1'b1;
  assign \A[14][189] [3] = 1'b1;
  assign \A[14][189] [2] = 1'b1;
  assign \A[14][189] [1] = 1'b1;
  assign \A[14][189] [0] = 1'b1;
  assign \A[14][190] [1] = 1'b1;
  assign \A[14][191] [0] = 1'b1;
  assign \A[14][193] [4] = 1'b1;
  assign \A[14][193] [3] = 1'b1;
  assign \A[14][193] [2] = 1'b1;
  assign \A[14][193] [1] = 1'b1;
  assign \A[14][194] [4] = 1'b1;
  assign \A[14][194] [3] = 1'b1;
  assign \A[14][194] [2] = 1'b1;
  assign \A[14][194] [1] = 1'b1;
  assign \A[14][194] [0] = 1'b1;
  assign \A[14][195] [1] = 1'b1;
  assign \A[14][195] [0] = 1'b1;
  assign \A[14][196] [0] = 1'b1;
  assign \A[14][198] [1] = 1'b1;
  assign \A[14][198] [0] = 1'b1;
  assign \A[14][200] [4] = 1'b1;
  assign \A[14][200] [3] = 1'b1;
  assign \A[14][200] [2] = 1'b1;
  assign \A[14][200] [1] = 1'b1;
  assign \A[14][201] [4] = 1'b1;
  assign \A[14][201] [3] = 1'b1;
  assign \A[14][201] [2] = 1'b1;
  assign \A[14][201] [1] = 1'b1;
  assign \A[14][201] [0] = 1'b1;
  assign \A[14][202] [0] = 1'b1;
  assign \A[14][203] [1] = 1'b1;
  assign \A[14][203] [0] = 1'b1;
  assign \A[14][204] [0] = 1'b1;
  assign \A[14][205] [0] = 1'b1;
  assign \A[14][206] [4] = 1'b1;
  assign \A[14][206] [3] = 1'b1;
  assign \A[14][206] [2] = 1'b1;
  assign \A[14][206] [1] = 1'b1;
  assign \A[14][206] [0] = 1'b1;
  assign \A[14][207] [4] = 1'b1;
  assign \A[14][207] [3] = 1'b1;
  assign \A[14][207] [2] = 1'b1;
  assign \A[14][207] [1] = 1'b1;
  assign \A[14][207] [0] = 1'b1;
  assign \A[14][208] [1] = 1'b1;
  assign \A[14][208] [0] = 1'b1;
  assign \A[14][209] [4] = 1'b1;
  assign \A[14][209] [3] = 1'b1;
  assign \A[14][209] [2] = 1'b1;
  assign \A[14][209] [1] = 1'b1;
  assign \A[14][209] [0] = 1'b1;
  assign \A[14][210] [4] = 1'b1;
  assign \A[14][210] [3] = 1'b1;
  assign \A[14][210] [2] = 1'b1;
  assign \A[14][210] [0] = 1'b1;
  assign \A[14][213] [4] = 1'b1;
  assign \A[14][213] [3] = 1'b1;
  assign \A[14][213] [2] = 1'b1;
  assign \A[14][213] [0] = 1'b1;
  assign \A[14][214] [4] = 1'b1;
  assign \A[14][214] [3] = 1'b1;
  assign \A[14][214] [2] = 1'b1;
  assign \A[14][214] [1] = 1'b1;
  assign \A[14][214] [0] = 1'b1;
  assign \A[14][216] [0] = 1'b1;
  assign \A[14][218] [1] = 1'b1;
  assign \A[14][219] [0] = 1'b1;
  assign \A[14][220] [4] = 1'b1;
  assign \A[14][220] [3] = 1'b1;
  assign \A[14][220] [2] = 1'b1;
  assign \A[14][220] [1] = 1'b1;
  assign \A[14][220] [0] = 1'b1;
  assign \A[14][221] [4] = 1'b1;
  assign \A[14][221] [3] = 1'b1;
  assign \A[14][221] [2] = 1'b1;
  assign \A[14][221] [1] = 1'b1;
  assign \A[14][221] [0] = 1'b1;
  assign \A[14][223] [0] = 1'b1;
  assign \A[14][224] [4] = 1'b1;
  assign \A[14][224] [3] = 1'b1;
  assign \A[14][224] [2] = 1'b1;
  assign \A[14][224] [0] = 1'b1;
  assign \A[14][225] [4] = 1'b1;
  assign \A[14][225] [3] = 1'b1;
  assign \A[14][225] [2] = 1'b1;
  assign \A[14][225] [1] = 1'b1;
  assign \A[14][225] [0] = 1'b1;
  assign \A[14][227] [4] = 1'b1;
  assign \A[14][227] [3] = 1'b1;
  assign \A[14][227] [2] = 1'b1;
  assign \A[14][227] [1] = 1'b1;
  assign \A[14][227] [0] = 1'b1;
  assign \A[14][228] [0] = 1'b1;
  assign \A[14][229] [0] = 1'b1;
  assign \A[14][230] [4] = 1'b1;
  assign \A[14][230] [3] = 1'b1;
  assign \A[14][230] [2] = 1'b1;
  assign \A[14][230] [1] = 1'b1;
  assign \A[14][230] [0] = 1'b1;
  assign \A[14][231] [4] = 1'b1;
  assign \A[14][231] [3] = 1'b1;
  assign \A[14][231] [2] = 1'b1;
  assign \A[14][231] [1] = 1'b1;
  assign \A[14][231] [0] = 1'b1;
  assign \A[14][232] [4] = 1'b1;
  assign \A[14][232] [3] = 1'b1;
  assign \A[14][232] [2] = 1'b1;
  assign \A[14][232] [1] = 1'b1;
  assign \A[14][232] [0] = 1'b1;
  assign \A[14][233] [0] = 1'b1;
  assign \A[14][234] [0] = 1'b1;
  assign \A[14][235] [4] = 1'b1;
  assign \A[14][235] [3] = 1'b1;
  assign \A[14][235] [2] = 1'b1;
  assign \A[14][235] [1] = 1'b1;
  assign \A[14][235] [0] = 1'b1;
  assign \A[14][236] [4] = 1'b1;
  assign \A[14][236] [3] = 1'b1;
  assign \A[14][236] [2] = 1'b1;
  assign \A[14][236] [1] = 1'b1;
  assign \A[14][236] [0] = 1'b1;
  assign \A[14][238] [4] = 1'b1;
  assign \A[14][238] [3] = 1'b1;
  assign \A[14][238] [2] = 1'b1;
  assign \A[14][238] [1] = 1'b1;
  assign \A[14][238] [0] = 1'b1;
  assign \A[14][239] [4] = 1'b1;
  assign \A[14][239] [3] = 1'b1;
  assign \A[14][239] [2] = 1'b1;
  assign \A[14][239] [1] = 1'b1;
  assign \A[14][239] [0] = 1'b1;
  assign \A[14][240] [0] = 1'b1;
  assign \A[14][241] [4] = 1'b1;
  assign \A[14][241] [3] = 1'b1;
  assign \A[14][241] [2] = 1'b1;
  assign \A[14][241] [1] = 1'b1;
  assign \A[14][243] [1] = 1'b1;
  assign \A[14][246] [4] = 1'b1;
  assign \A[14][246] [3] = 1'b1;
  assign \A[14][246] [2] = 1'b1;
  assign \A[14][246] [1] = 1'b1;
  assign \A[14][246] [0] = 1'b1;
  assign \A[14][248] [4] = 1'b1;
  assign \A[14][248] [3] = 1'b1;
  assign \A[14][248] [2] = 1'b1;
  assign \A[14][248] [1] = 1'b1;
  assign \A[14][249] [4] = 1'b1;
  assign \A[14][249] [3] = 1'b1;
  assign \A[14][249] [1] = 1'b1;
  assign \A[14][249] [0] = 1'b1;
  assign \A[14][250] [0] = 1'b1;
  assign \A[14][251] [4] = 1'b1;
  assign \A[14][251] [3] = 1'b1;
  assign \A[14][251] [2] = 1'b1;
  assign \A[14][251] [1] = 1'b1;
  assign \A[14][251] [0] = 1'b1;
  assign \A[14][252] [4] = 1'b1;
  assign \A[14][252] [3] = 1'b1;
  assign \A[14][252] [2] = 1'b1;
  assign \A[14][252] [1] = 1'b1;
  assign \A[14][252] [0] = 1'b1;
  assign \A[14][253] [1] = 1'b1;
  assign \A[14][254] [1] = 1'b1;
  assign \A[14][254] [0] = 1'b1;
  assign \A[14][255] [1] = 1'b1;
  assign \A[14][255] [0] = 1'b1;
  assign \A[15][1] [1] = 1'b1;
  assign \A[15][2] [1] = 1'b1;
  assign \A[15][3] [4] = 1'b1;
  assign \A[15][3] [3] = 1'b1;
  assign \A[15][3] [2] = 1'b1;
  assign \A[15][3] [1] = 1'b1;
  assign \A[15][7] [4] = 1'b1;
  assign \A[15][7] [3] = 1'b1;
  assign \A[15][7] [2] = 1'b1;
  assign \A[15][7] [1] = 1'b1;
  assign \A[15][7] [0] = 1'b1;
  assign \A[15][9] [0] = 1'b1;
  assign \A[15][10] [4] = 1'b1;
  assign \A[15][10] [3] = 1'b1;
  assign \A[15][10] [2] = 1'b1;
  assign \A[15][10] [1] = 1'b1;
  assign \A[15][11] [4] = 1'b1;
  assign \A[15][11] [3] = 1'b1;
  assign \A[15][11] [2] = 1'b1;
  assign \A[15][11] [1] = 1'b1;
  assign \A[15][11] [0] = 1'b1;
  assign \A[15][12] [4] = 1'b1;
  assign \A[15][12] [3] = 1'b1;
  assign \A[15][12] [2] = 1'b1;
  assign \A[15][12] [1] = 1'b1;
  assign \A[15][12] [0] = 1'b1;
  assign \A[15][13] [4] = 1'b1;
  assign \A[15][13] [3] = 1'b1;
  assign \A[15][13] [2] = 1'b1;
  assign \A[15][13] [1] = 1'b1;
  assign \A[15][15] [4] = 1'b1;
  assign \A[15][15] [3] = 1'b1;
  assign \A[15][15] [2] = 1'b1;
  assign \A[15][15] [1] = 1'b1;
  assign \A[15][15] [0] = 1'b1;
  assign \A[15][16] [4] = 1'b1;
  assign \A[15][16] [3] = 1'b1;
  assign \A[15][16] [2] = 1'b1;
  assign \A[15][16] [1] = 1'b1;
  assign \A[15][16] [0] = 1'b1;
  assign \A[15][17] [4] = 1'b1;
  assign \A[15][17] [3] = 1'b1;
  assign \A[15][17] [2] = 1'b1;
  assign \A[15][17] [1] = 1'b1;
  assign \A[15][17] [0] = 1'b1;
  assign \A[15][18] [4] = 1'b1;
  assign \A[15][18] [3] = 1'b1;
  assign \A[15][18] [2] = 1'b1;
  assign \A[15][18] [1] = 1'b1;
  assign \A[15][18] [0] = 1'b1;
  assign \A[15][19] [4] = 1'b1;
  assign \A[15][19] [3] = 1'b1;
  assign \A[15][19] [2] = 1'b1;
  assign \A[15][19] [1] = 1'b1;
  assign \A[15][19] [0] = 1'b1;
  assign \A[15][20] [0] = 1'b1;
  assign \A[15][21] [4] = 1'b1;
  assign \A[15][21] [3] = 1'b1;
  assign \A[15][21] [2] = 1'b1;
  assign \A[15][21] [1] = 1'b1;
  assign \A[15][22] [4] = 1'b1;
  assign \A[15][22] [3] = 1'b1;
  assign \A[15][22] [2] = 1'b1;
  assign \A[15][22] [1] = 1'b1;
  assign \A[15][24] [4] = 1'b1;
  assign \A[15][24] [3] = 1'b1;
  assign \A[15][24] [2] = 1'b1;
  assign \A[15][24] [1] = 1'b1;
  assign \A[15][24] [0] = 1'b1;
  assign \A[15][26] [4] = 1'b1;
  assign \A[15][26] [3] = 1'b1;
  assign \A[15][26] [2] = 1'b1;
  assign \A[15][26] [1] = 1'b1;
  assign \A[15][27] [4] = 1'b1;
  assign \A[15][27] [3] = 1'b1;
  assign \A[15][27] [2] = 1'b1;
  assign \A[15][27] [1] = 1'b1;
  assign \A[15][27] [0] = 1'b1;
  assign \A[15][28] [4] = 1'b1;
  assign \A[15][28] [3] = 1'b1;
  assign \A[15][28] [2] = 1'b1;
  assign \A[15][28] [1] = 1'b1;
  assign \A[15][29] [0] = 1'b1;
  assign \A[15][31] [4] = 1'b1;
  assign \A[15][31] [3] = 1'b1;
  assign \A[15][31] [2] = 1'b1;
  assign \A[15][31] [1] = 1'b1;
  assign \A[15][31] [0] = 1'b1;
  assign \A[15][32] [4] = 1'b1;
  assign \A[15][32] [3] = 1'b1;
  assign \A[15][32] [2] = 1'b1;
  assign \A[15][32] [1] = 1'b1;
  assign \A[15][33] [0] = 1'b1;
  assign \A[15][34] [4] = 1'b1;
  assign \A[15][34] [3] = 1'b1;
  assign \A[15][34] [2] = 1'b1;
  assign \A[15][34] [1] = 1'b1;
  assign \A[15][35] [0] = 1'b1;
  assign \A[15][36] [4] = 1'b1;
  assign \A[15][36] [3] = 1'b1;
  assign \A[15][36] [2] = 1'b1;
  assign \A[15][36] [1] = 1'b1;
  assign \A[15][37] [4] = 1'b1;
  assign \A[15][37] [3] = 1'b1;
  assign \A[15][37] [2] = 1'b1;
  assign \A[15][37] [1] = 1'b1;
  assign \A[15][37] [0] = 1'b1;
  assign \A[15][38] [4] = 1'b1;
  assign \A[15][38] [3] = 1'b1;
  assign \A[15][38] [2] = 1'b1;
  assign \A[15][38] [1] = 1'b1;
  assign \A[15][40] [0] = 1'b1;
  assign \A[15][41] [0] = 1'b1;
  assign \A[15][42] [4] = 1'b1;
  assign \A[15][42] [3] = 1'b1;
  assign \A[15][42] [2] = 1'b1;
  assign \A[15][42] [0] = 1'b1;
  assign \A[15][43] [4] = 1'b1;
  assign \A[15][43] [3] = 1'b1;
  assign \A[15][43] [2] = 1'b1;
  assign \A[15][43] [1] = 1'b1;
  assign \A[15][44] [4] = 1'b1;
  assign \A[15][44] [3] = 1'b1;
  assign \A[15][44] [2] = 1'b1;
  assign \A[15][44] [1] = 1'b1;
  assign \A[15][44] [0] = 1'b1;
  assign \A[15][45] [4] = 1'b1;
  assign \A[15][45] [3] = 1'b1;
  assign \A[15][45] [2] = 1'b1;
  assign \A[15][45] [1] = 1'b1;
  assign \A[15][45] [0] = 1'b1;
  assign \A[15][47] [1] = 1'b1;
  assign \A[15][49] [1] = 1'b1;
  assign \A[15][50] [1] = 1'b1;
  assign \A[15][52] [4] = 1'b1;
  assign \A[15][52] [3] = 1'b1;
  assign \A[15][52] [2] = 1'b1;
  assign \A[15][52] [1] = 1'b1;
  assign \A[15][52] [0] = 1'b1;
  assign \A[15][53] [4] = 1'b1;
  assign \A[15][53] [3] = 1'b1;
  assign \A[15][53] [2] = 1'b1;
  assign \A[15][53] [1] = 1'b1;
  assign \A[15][53] [0] = 1'b1;
  assign \A[15][54] [1] = 1'b1;
  assign \A[15][55] [4] = 1'b1;
  assign \A[15][55] [3] = 1'b1;
  assign \A[15][55] [2] = 1'b1;
  assign \A[15][55] [1] = 1'b1;
  assign \A[15][55] [0] = 1'b1;
  assign \A[15][56] [0] = 1'b1;
  assign \A[15][57] [0] = 1'b1;
  assign \A[15][58] [2] = 1'b1;
  assign \A[15][59] [4] = 1'b1;
  assign \A[15][59] [3] = 1'b1;
  assign \A[15][59] [2] = 1'b1;
  assign \A[15][59] [1] = 1'b1;
  assign \A[15][59] [0] = 1'b1;
  assign \A[15][60] [0] = 1'b1;
  assign \A[15][61] [4] = 1'b1;
  assign \A[15][61] [3] = 1'b1;
  assign \A[15][61] [2] = 1'b1;
  assign \A[15][61] [1] = 1'b1;
  assign \A[15][64] [4] = 1'b1;
  assign \A[15][64] [3] = 1'b1;
  assign \A[15][64] [2] = 1'b1;
  assign \A[15][64] [1] = 1'b1;
  assign \A[15][64] [0] = 1'b1;
  assign \A[15][65] [0] = 1'b1;
  assign \A[15][67] [0] = 1'b1;
  assign \A[15][69] [4] = 1'b1;
  assign \A[15][69] [3] = 1'b1;
  assign \A[15][69] [2] = 1'b1;
  assign \A[15][69] [1] = 1'b1;
  assign \A[15][69] [0] = 1'b1;
  assign \A[15][70] [1] = 1'b1;
  assign \A[15][71] [1] = 1'b1;
  assign \A[15][72] [4] = 1'b1;
  assign \A[15][72] [3] = 1'b1;
  assign \A[15][72] [2] = 1'b1;
  assign \A[15][72] [1] = 1'b1;
  assign \A[15][72] [0] = 1'b1;
  assign \A[15][73] [4] = 1'b1;
  assign \A[15][73] [3] = 1'b1;
  assign \A[15][73] [2] = 1'b1;
  assign \A[15][73] [1] = 1'b1;
  assign \A[15][74] [4] = 1'b1;
  assign \A[15][74] [3] = 1'b1;
  assign \A[15][74] [2] = 1'b1;
  assign \A[15][74] [0] = 1'b1;
  assign \A[15][75] [0] = 1'b1;
  assign \A[15][76] [4] = 1'b1;
  assign \A[15][76] [3] = 1'b1;
  assign \A[15][76] [2] = 1'b1;
  assign \A[15][76] [1] = 1'b1;
  assign \A[15][76] [0] = 1'b1;
  assign \A[15][78] [0] = 1'b1;
  assign \A[15][80] [0] = 1'b1;
  assign \A[15][81] [4] = 1'b1;
  assign \A[15][81] [3] = 1'b1;
  assign \A[15][81] [2] = 1'b1;
  assign \A[15][81] [0] = 1'b1;
  assign \A[15][83] [4] = 1'b1;
  assign \A[15][83] [3] = 1'b1;
  assign \A[15][83] [2] = 1'b1;
  assign \A[15][83] [1] = 1'b1;
  assign \A[15][85] [1] = 1'b1;
  assign \A[15][86] [4] = 1'b1;
  assign \A[15][86] [3] = 1'b1;
  assign \A[15][86] [2] = 1'b1;
  assign \A[15][86] [1] = 1'b1;
  assign \A[15][91] [0] = 1'b1;
  assign \A[15][92] [0] = 1'b1;
  assign \A[15][93] [4] = 1'b1;
  assign \A[15][93] [3] = 1'b1;
  assign \A[15][93] [2] = 1'b1;
  assign \A[15][93] [1] = 1'b1;
  assign \A[15][94] [0] = 1'b1;
  assign \A[15][96] [0] = 1'b1;
  assign \A[15][97] [4] = 1'b1;
  assign \A[15][97] [3] = 1'b1;
  assign \A[15][97] [2] = 1'b1;
  assign \A[15][97] [1] = 1'b1;
  assign \A[15][97] [0] = 1'b1;
  assign \A[15][98] [0] = 1'b1;
  assign \A[15][99] [1] = 1'b1;
  assign \A[15][99] [0] = 1'b1;
  assign \A[15][100] [4] = 1'b1;
  assign \A[15][100] [3] = 1'b1;
  assign \A[15][100] [2] = 1'b1;
  assign \A[15][100] [0] = 1'b1;
  assign \A[15][101] [1] = 1'b1;
  assign \A[15][101] [0] = 1'b1;
  assign \A[15][102] [0] = 1'b1;
  assign \A[15][103] [4] = 1'b1;
  assign \A[15][103] [3] = 1'b1;
  assign \A[15][103] [2] = 1'b1;
  assign \A[15][103] [1] = 1'b1;
  assign \A[15][103] [0] = 1'b1;
  assign \A[15][104] [0] = 1'b1;
  assign \A[15][105] [4] = 1'b1;
  assign \A[15][105] [3] = 1'b1;
  assign \A[15][105] [2] = 1'b1;
  assign \A[15][105] [1] = 1'b1;
  assign \A[15][106] [0] = 1'b1;
  assign \A[15][107] [4] = 1'b1;
  assign \A[15][107] [3] = 1'b1;
  assign \A[15][107] [2] = 1'b1;
  assign \A[15][107] [1] = 1'b1;
  assign \A[15][107] [0] = 1'b1;
  assign \A[15][108] [4] = 1'b1;
  assign \A[15][108] [3] = 1'b1;
  assign \A[15][108] [2] = 1'b1;
  assign \A[15][108] [1] = 1'b1;
  assign \A[15][108] [0] = 1'b1;
  assign \A[15][109] [0] = 1'b1;
  assign \A[15][111] [4] = 1'b1;
  assign \A[15][111] [3] = 1'b1;
  assign \A[15][111] [2] = 1'b1;
  assign \A[15][111] [1] = 1'b1;
  assign \A[15][113] [4] = 1'b1;
  assign \A[15][113] [3] = 1'b1;
  assign \A[15][113] [2] = 1'b1;
  assign \A[15][113] [1] = 1'b1;
  assign \A[15][113] [0] = 1'b1;
  assign \A[15][114] [4] = 1'b1;
  assign \A[15][114] [3] = 1'b1;
  assign \A[15][114] [2] = 1'b1;
  assign \A[15][114] [1] = 1'b1;
  assign \A[15][114] [0] = 1'b1;
  assign \A[15][115] [1] = 1'b1;
  assign \A[15][117] [4] = 1'b1;
  assign \A[15][117] [3] = 1'b1;
  assign \A[15][117] [2] = 1'b1;
  assign \A[15][117] [1] = 1'b1;
  assign \A[15][117] [0] = 1'b1;
  assign \A[15][118] [0] = 1'b1;
  assign \A[15][119] [4] = 1'b1;
  assign \A[15][119] [3] = 1'b1;
  assign \A[15][119] [2] = 1'b1;
  assign \A[15][119] [1] = 1'b1;
  assign \A[15][119] [0] = 1'b1;
  assign \A[15][125] [4] = 1'b1;
  assign \A[15][125] [3] = 1'b1;
  assign \A[15][125] [2] = 1'b1;
  assign \A[15][125] [0] = 1'b1;
  assign \A[15][126] [1] = 1'b1;
  assign \A[15][127] [0] = 1'b1;
  assign \A[15][128] [4] = 1'b1;
  assign \A[15][128] [3] = 1'b1;
  assign \A[15][128] [2] = 1'b1;
  assign \A[15][128] [1] = 1'b1;
  assign \A[15][128] [0] = 1'b1;
  assign \A[15][130] [4] = 1'b1;
  assign \A[15][130] [3] = 1'b1;
  assign \A[15][130] [2] = 1'b1;
  assign \A[15][130] [1] = 1'b1;
  assign \A[15][130] [0] = 1'b1;
  assign \A[15][131] [4] = 1'b1;
  assign \A[15][131] [3] = 1'b1;
  assign \A[15][131] [2] = 1'b1;
  assign \A[15][131] [1] = 1'b1;
  assign \A[15][131] [0] = 1'b1;
  assign \A[15][132] [4] = 1'b1;
  assign \A[15][132] [3] = 1'b1;
  assign \A[15][132] [2] = 1'b1;
  assign \A[15][132] [1] = 1'b1;
  assign \A[15][133] [4] = 1'b1;
  assign \A[15][133] [3] = 1'b1;
  assign \A[15][133] [2] = 1'b1;
  assign \A[15][133] [1] = 1'b1;
  assign \A[15][133] [0] = 1'b1;
  assign \A[15][134] [4] = 1'b1;
  assign \A[15][134] [3] = 1'b1;
  assign \A[15][134] [2] = 1'b1;
  assign \A[15][134] [1] = 1'b1;
  assign \A[15][135] [4] = 1'b1;
  assign \A[15][135] [3] = 1'b1;
  assign \A[15][135] [2] = 1'b1;
  assign \A[15][135] [1] = 1'b1;
  assign \A[15][137] [0] = 1'b1;
  assign \A[15][139] [4] = 1'b1;
  assign \A[15][139] [3] = 1'b1;
  assign \A[15][139] [2] = 1'b1;
  assign \A[15][139] [1] = 1'b1;
  assign \A[15][140] [1] = 1'b1;
  assign \A[15][140] [0] = 1'b1;
  assign \A[15][141] [0] = 1'b1;
  assign \A[15][143] [4] = 1'b1;
  assign \A[15][143] [3] = 1'b1;
  assign \A[15][143] [2] = 1'b1;
  assign \A[15][143] [1] = 1'b1;
  assign \A[15][144] [4] = 1'b1;
  assign \A[15][144] [3] = 1'b1;
  assign \A[15][144] [2] = 1'b1;
  assign \A[15][144] [1] = 1'b1;
  assign \A[15][144] [0] = 1'b1;
  assign \A[15][145] [4] = 1'b1;
  assign \A[15][145] [3] = 1'b1;
  assign \A[15][145] [2] = 1'b1;
  assign \A[15][145] [1] = 1'b1;
  assign \A[15][146] [0] = 1'b1;
  assign \A[15][148] [4] = 1'b1;
  assign \A[15][148] [3] = 1'b1;
  assign \A[15][148] [2] = 1'b1;
  assign \A[15][148] [1] = 1'b1;
  assign \A[15][148] [0] = 1'b1;
  assign \A[15][151] [4] = 1'b1;
  assign \A[15][151] [3] = 1'b1;
  assign \A[15][151] [2] = 1'b1;
  assign \A[15][151] [1] = 1'b1;
  assign \A[15][151] [0] = 1'b1;
  assign \A[15][152] [4] = 1'b1;
  assign \A[15][152] [3] = 1'b1;
  assign \A[15][152] [2] = 1'b1;
  assign \A[15][152] [1] = 1'b1;
  assign \A[15][153] [4] = 1'b1;
  assign \A[15][153] [3] = 1'b1;
  assign \A[15][153] [2] = 1'b1;
  assign \A[15][153] [1] = 1'b1;
  assign \A[15][153] [0] = 1'b1;
  assign \A[15][154] [4] = 1'b1;
  assign \A[15][154] [3] = 1'b1;
  assign \A[15][154] [2] = 1'b1;
  assign \A[15][154] [0] = 1'b1;
  assign \A[15][156] [2] = 1'b1;
  assign \A[15][158] [4] = 1'b1;
  assign \A[15][158] [3] = 1'b1;
  assign \A[15][158] [2] = 1'b1;
  assign \A[15][158] [1] = 1'b1;
  assign \A[15][158] [0] = 1'b1;
  assign \A[15][159] [0] = 1'b1;
  assign \A[15][160] [0] = 1'b1;
  assign \A[15][162] [4] = 1'b1;
  assign \A[15][162] [3] = 1'b1;
  assign \A[15][162] [2] = 1'b1;
  assign \A[15][162] [1] = 1'b1;
  assign \A[15][162] [0] = 1'b1;
  assign \A[15][163] [4] = 1'b1;
  assign \A[15][163] [3] = 1'b1;
  assign \A[15][163] [2] = 1'b1;
  assign \A[15][163] [1] = 1'b1;
  assign \A[15][163] [0] = 1'b1;
  assign \A[15][165] [0] = 1'b1;
  assign \A[15][166] [0] = 1'b1;
  assign \A[15][169] [4] = 1'b1;
  assign \A[15][169] [3] = 1'b1;
  assign \A[15][169] [2] = 1'b1;
  assign \A[15][169] [0] = 1'b1;
  assign \A[15][170] [1] = 1'b1;
  assign \A[15][172] [4] = 1'b1;
  assign \A[15][172] [3] = 1'b1;
  assign \A[15][172] [2] = 1'b1;
  assign \A[15][172] [1] = 1'b1;
  assign \A[15][173] [4] = 1'b1;
  assign \A[15][173] [3] = 1'b1;
  assign \A[15][173] [2] = 1'b1;
  assign \A[15][173] [0] = 1'b1;
  assign \A[15][174] [4] = 1'b1;
  assign \A[15][174] [3] = 1'b1;
  assign \A[15][174] [2] = 1'b1;
  assign \A[15][174] [1] = 1'b1;
  assign \A[15][174] [0] = 1'b1;
  assign \A[15][175] [0] = 1'b1;
  assign \A[15][176] [4] = 1'b1;
  assign \A[15][176] [3] = 1'b1;
  assign \A[15][176] [2] = 1'b1;
  assign \A[15][176] [1] = 1'b1;
  assign \A[15][176] [0] = 1'b1;
  assign \A[15][177] [4] = 1'b1;
  assign \A[15][177] [3] = 1'b1;
  assign \A[15][177] [2] = 1'b1;
  assign \A[15][177] [1] = 1'b1;
  assign \A[15][178] [4] = 1'b1;
  assign \A[15][178] [3] = 1'b1;
  assign \A[15][178] [2] = 1'b1;
  assign \A[15][178] [1] = 1'b1;
  assign \A[15][179] [4] = 1'b1;
  assign \A[15][179] [3] = 1'b1;
  assign \A[15][179] [2] = 1'b1;
  assign \A[15][179] [1] = 1'b1;
  assign \A[15][179] [0] = 1'b1;
  assign \A[15][180] [0] = 1'b1;
  assign \A[15][181] [4] = 1'b1;
  assign \A[15][181] [3] = 1'b1;
  assign \A[15][181] [2] = 1'b1;
  assign \A[15][181] [1] = 1'b1;
  assign \A[15][182] [4] = 1'b1;
  assign \A[15][182] [3] = 1'b1;
  assign \A[15][182] [2] = 1'b1;
  assign \A[15][182] [1] = 1'b1;
  assign \A[15][182] [0] = 1'b1;
  assign \A[15][184] [0] = 1'b1;
  assign \A[15][185] [0] = 1'b1;
  assign \A[15][186] [4] = 1'b1;
  assign \A[15][186] [3] = 1'b1;
  assign \A[15][186] [2] = 1'b1;
  assign \A[15][186] [1] = 1'b1;
  assign \A[15][186] [0] = 1'b1;
  assign \A[15][188] [0] = 1'b1;
  assign \A[15][189] [4] = 1'b1;
  assign \A[15][189] [3] = 1'b1;
  assign \A[15][189] [2] = 1'b1;
  assign \A[15][189] [0] = 1'b1;
  assign \A[15][190] [1] = 1'b1;
  assign \A[15][192] [0] = 1'b1;
  assign \A[15][193] [0] = 1'b1;
  assign \A[15][195] [4] = 1'b1;
  assign \A[15][195] [3] = 1'b1;
  assign \A[15][195] [2] = 1'b1;
  assign \A[15][195] [1] = 1'b1;
  assign \A[15][195] [0] = 1'b1;
  assign \A[15][196] [4] = 1'b1;
  assign \A[15][196] [3] = 1'b1;
  assign \A[15][196] [2] = 1'b1;
  assign \A[15][196] [1] = 1'b1;
  assign \A[15][196] [0] = 1'b1;
  assign \A[15][198] [4] = 1'b1;
  assign \A[15][198] [3] = 1'b1;
  assign \A[15][198] [2] = 1'b1;
  assign \A[15][198] [1] = 1'b1;
  assign \A[15][199] [4] = 1'b1;
  assign \A[15][199] [3] = 1'b1;
  assign \A[15][199] [2] = 1'b1;
  assign \A[15][199] [1] = 1'b1;
  assign \A[15][199] [0] = 1'b1;
  assign \A[15][200] [4] = 1'b1;
  assign \A[15][200] [3] = 1'b1;
  assign \A[15][200] [2] = 1'b1;
  assign \A[15][200] [1] = 1'b1;
  assign \A[15][200] [0] = 1'b1;
  assign \A[15][202] [1] = 1'b1;
  assign \A[15][204] [4] = 1'b1;
  assign \A[15][204] [3] = 1'b1;
  assign \A[15][204] [2] = 1'b1;
  assign \A[15][204] [1] = 1'b1;
  assign \A[15][204] [0] = 1'b1;
  assign \A[15][205] [4] = 1'b1;
  assign \A[15][205] [3] = 1'b1;
  assign \A[15][205] [2] = 1'b1;
  assign \A[15][205] [1] = 1'b1;
  assign \A[15][205] [0] = 1'b1;
  assign \A[15][206] [4] = 1'b1;
  assign \A[15][206] [3] = 1'b1;
  assign \A[15][206] [2] = 1'b1;
  assign \A[15][206] [1] = 1'b1;
  assign \A[15][206] [0] = 1'b1;
  assign \A[15][209] [0] = 1'b1;
  assign \A[15][210] [0] = 1'b1;
  assign \A[15][212] [4] = 1'b1;
  assign \A[15][212] [3] = 1'b1;
  assign \A[15][212] [2] = 1'b1;
  assign \A[15][212] [1] = 1'b1;
  assign \A[15][212] [0] = 1'b1;
  assign \A[15][213] [4] = 1'b1;
  assign \A[15][213] [3] = 1'b1;
  assign \A[15][213] [2] = 1'b1;
  assign \A[15][213] [1] = 1'b1;
  assign \A[15][214] [1] = 1'b1;
  assign \A[15][215] [4] = 1'b1;
  assign \A[15][215] [3] = 1'b1;
  assign \A[15][215] [2] = 1'b1;
  assign \A[15][215] [1] = 1'b1;
  assign \A[15][215] [0] = 1'b1;
  assign \A[15][216] [0] = 1'b1;
  assign \A[15][217] [0] = 1'b1;
  assign \A[15][218] [4] = 1'b1;
  assign \A[15][218] [3] = 1'b1;
  assign \A[15][218] [2] = 1'b1;
  assign \A[15][218] [1] = 1'b1;
  assign \A[15][218] [0] = 1'b1;
  assign \A[15][219] [0] = 1'b1;
  assign \A[15][220] [4] = 1'b1;
  assign \A[15][220] [3] = 1'b1;
  assign \A[15][220] [2] = 1'b1;
  assign \A[15][220] [1] = 1'b1;
  assign \A[15][221] [4] = 1'b1;
  assign \A[15][221] [3] = 1'b1;
  assign \A[15][221] [2] = 1'b1;
  assign \A[15][221] [1] = 1'b1;
  assign \A[15][221] [0] = 1'b1;
  assign \A[15][222] [4] = 1'b1;
  assign \A[15][222] [3] = 1'b1;
  assign \A[15][222] [2] = 1'b1;
  assign \A[15][222] [1] = 1'b1;
  assign \A[15][223] [4] = 1'b1;
  assign \A[15][223] [3] = 1'b1;
  assign \A[15][223] [2] = 1'b1;
  assign \A[15][223] [1] = 1'b1;
  assign \A[15][223] [0] = 1'b1;
  assign \A[15][225] [1] = 1'b1;
  assign \A[15][225] [0] = 1'b1;
  assign \A[15][227] [1] = 1'b1;
  assign \A[15][229] [4] = 1'b1;
  assign \A[15][229] [3] = 1'b1;
  assign \A[15][229] [2] = 1'b1;
  assign \A[15][229] [1] = 1'b1;
  assign \A[15][229] [0] = 1'b1;
  assign \A[15][232] [4] = 1'b1;
  assign \A[15][232] [3] = 1'b1;
  assign \A[15][232] [2] = 1'b1;
  assign \A[15][232] [1] = 1'b1;
  assign \A[15][232] [0] = 1'b1;
  assign \A[15][233] [0] = 1'b1;
  assign \A[15][234] [4] = 1'b1;
  assign \A[15][234] [3] = 1'b1;
  assign \A[15][234] [2] = 1'b1;
  assign \A[15][234] [1] = 1'b1;
  assign \A[15][234] [0] = 1'b1;
  assign \A[15][237] [1] = 1'b1;
  assign \A[15][238] [4] = 1'b1;
  assign \A[15][238] [3] = 1'b1;
  assign \A[15][238] [2] = 1'b1;
  assign \A[15][238] [1] = 1'b1;
  assign \A[15][238] [0] = 1'b1;
  assign \A[15][240] [1] = 1'b1;
  assign \A[15][241] [0] = 1'b1;
  assign \A[15][242] [1] = 1'b1;
  assign \A[15][243] [4] = 1'b1;
  assign \A[15][243] [3] = 1'b1;
  assign \A[15][243] [2] = 1'b1;
  assign \A[15][243] [1] = 1'b1;
  assign \A[15][245] [4] = 1'b1;
  assign \A[15][245] [3] = 1'b1;
  assign \A[15][245] [2] = 1'b1;
  assign \A[15][245] [1] = 1'b1;
  assign \A[15][245] [0] = 1'b1;
  assign \A[15][246] [0] = 1'b1;
  assign \A[15][248] [4] = 1'b1;
  assign \A[15][248] [3] = 1'b1;
  assign \A[15][248] [2] = 1'b1;
  assign \A[15][248] [0] = 1'b1;
  assign \A[15][250] [1] = 1'b1;
  assign \A[15][251] [0] = 1'b1;
  assign \A[15][252] [0] = 1'b1;
  assign \A[15][254] [0] = 1'b1;
  assign \A[15][255] [4] = 1'b1;
  assign \A[15][255] [3] = 1'b1;
  assign \A[15][255] [2] = 1'b1;
  assign \A[15][255] [1] = 1'b1;
  assign \A[15][255] [0] = 1'b1;
  assign \A[16][2] [4] = 1'b1;
  assign \A[16][2] [3] = 1'b1;
  assign \A[16][2] [2] = 1'b1;
  assign \A[16][2] [1] = 1'b1;
  assign \A[16][2] [0] = 1'b1;
  assign \A[16][3] [4] = 1'b1;
  assign \A[16][3] [3] = 1'b1;
  assign \A[16][3] [2] = 1'b1;
  assign \A[16][3] [1] = 1'b1;
  assign \A[16][5] [1] = 1'b1;
  assign \A[16][6] [4] = 1'b1;
  assign \A[16][6] [3] = 1'b1;
  assign \A[16][6] [2] = 1'b1;
  assign \A[16][6] [1] = 1'b1;
  assign \A[16][7] [4] = 1'b1;
  assign \A[16][7] [3] = 1'b1;
  assign \A[16][7] [2] = 1'b1;
  assign \A[16][7] [1] = 1'b1;
  assign \A[16][7] [0] = 1'b1;
  assign \A[16][8] [4] = 1'b1;
  assign \A[16][8] [3] = 1'b1;
  assign \A[16][8] [2] = 1'b1;
  assign \A[16][8] [1] = 1'b1;
  assign \A[16][8] [0] = 1'b1;
  assign \A[16][9] [1] = 1'b1;
  assign \A[16][10] [4] = 1'b1;
  assign \A[16][10] [3] = 1'b1;
  assign \A[16][10] [2] = 1'b1;
  assign \A[16][10] [1] = 1'b1;
  assign \A[16][10] [0] = 1'b1;
  assign \A[16][12] [1] = 1'b1;
  assign \A[16][12] [0] = 1'b1;
  assign \A[16][13] [4] = 1'b1;
  assign \A[16][13] [3] = 1'b1;
  assign \A[16][13] [2] = 1'b1;
  assign \A[16][13] [1] = 1'b1;
  assign \A[16][14] [4] = 1'b1;
  assign \A[16][14] [3] = 1'b1;
  assign \A[16][14] [2] = 1'b1;
  assign \A[16][15] [4] = 1'b1;
  assign \A[16][15] [3] = 1'b1;
  assign \A[16][15] [2] = 1'b1;
  assign \A[16][15] [1] = 1'b1;
  assign \A[16][16] [1] = 1'b1;
  assign \A[16][16] [0] = 1'b1;
  assign \A[16][18] [4] = 1'b1;
  assign \A[16][18] [3] = 1'b1;
  assign \A[16][18] [2] = 1'b1;
  assign \A[16][18] [1] = 1'b1;
  assign \A[16][18] [0] = 1'b1;
  assign \A[16][19] [4] = 1'b1;
  assign \A[16][19] [3] = 1'b1;
  assign \A[16][19] [2] = 1'b1;
  assign \A[16][19] [0] = 1'b1;
  assign \A[16][20] [4] = 1'b1;
  assign \A[16][20] [3] = 1'b1;
  assign \A[16][20] [2] = 1'b1;
  assign \A[16][20] [1] = 1'b1;
  assign \A[16][20] [0] = 1'b1;
  assign \A[16][21] [4] = 1'b1;
  assign \A[16][21] [3] = 1'b1;
  assign \A[16][21] [2] = 1'b1;
  assign \A[16][21] [1] = 1'b1;
  assign \A[16][22] [4] = 1'b1;
  assign \A[16][22] [3] = 1'b1;
  assign \A[16][22] [2] = 1'b1;
  assign \A[16][22] [1] = 1'b1;
  assign \A[16][22] [0] = 1'b1;
  assign \A[16][23] [4] = 1'b1;
  assign \A[16][23] [3] = 1'b1;
  assign \A[16][23] [2] = 1'b1;
  assign \A[16][23] [1] = 1'b1;
  assign \A[16][24] [4] = 1'b1;
  assign \A[16][24] [3] = 1'b1;
  assign \A[16][24] [2] = 1'b1;
  assign \A[16][24] [1] = 1'b1;
  assign \A[16][24] [0] = 1'b1;
  assign \A[16][26] [4] = 1'b1;
  assign \A[16][26] [3] = 1'b1;
  assign \A[16][26] [2] = 1'b1;
  assign \A[16][26] [1] = 1'b1;
  assign \A[16][26] [0] = 1'b1;
  assign \A[16][27] [0] = 1'b1;
  assign \A[16][28] [4] = 1'b1;
  assign \A[16][28] [3] = 1'b1;
  assign \A[16][28] [2] = 1'b1;
  assign \A[16][28] [0] = 1'b1;
  assign \A[16][30] [0] = 1'b1;
  assign \A[16][33] [0] = 1'b1;
  assign \A[16][36] [4] = 1'b1;
  assign \A[16][36] [3] = 1'b1;
  assign \A[16][36] [2] = 1'b1;
  assign \A[16][36] [1] = 1'b1;
  assign \A[16][37] [4] = 1'b1;
  assign \A[16][37] [3] = 1'b1;
  assign \A[16][37] [2] = 1'b1;
  assign \A[16][37] [1] = 1'b1;
  assign \A[16][37] [0] = 1'b1;
  assign \A[16][39] [0] = 1'b1;
  assign \A[16][41] [4] = 1'b1;
  assign \A[16][41] [3] = 1'b1;
  assign \A[16][41] [2] = 1'b1;
  assign \A[16][41] [1] = 1'b1;
  assign \A[16][42] [4] = 1'b1;
  assign \A[16][42] [3] = 1'b1;
  assign \A[16][42] [2] = 1'b1;
  assign \A[16][42] [1] = 1'b1;
  assign \A[16][42] [0] = 1'b1;
  assign \A[16][43] [4] = 1'b1;
  assign \A[16][43] [3] = 1'b1;
  assign \A[16][43] [2] = 1'b1;
  assign \A[16][43] [1] = 1'b1;
  assign \A[16][44] [4] = 1'b1;
  assign \A[16][44] [3] = 1'b1;
  assign \A[16][44] [2] = 1'b1;
  assign \A[16][44] [1] = 1'b1;
  assign \A[16][45] [4] = 1'b1;
  assign \A[16][45] [3] = 1'b1;
  assign \A[16][45] [2] = 1'b1;
  assign \A[16][45] [1] = 1'b1;
  assign \A[16][46] [1] = 1'b1;
  assign \A[16][47] [4] = 1'b1;
  assign \A[16][47] [3] = 1'b1;
  assign \A[16][47] [2] = 1'b1;
  assign \A[16][47] [1] = 1'b1;
  assign \A[16][50] [0] = 1'b1;
  assign \A[16][51] [1] = 1'b1;
  assign \A[16][52] [0] = 1'b1;
  assign \A[16][53] [4] = 1'b1;
  assign \A[16][53] [3] = 1'b1;
  assign \A[16][53] [2] = 1'b1;
  assign \A[16][53] [1] = 1'b1;
  assign \A[16][53] [0] = 1'b1;
  assign \A[16][54] [1] = 1'b1;
  assign \A[16][55] [4] = 1'b1;
  assign \A[16][55] [3] = 1'b1;
  assign \A[16][55] [2] = 1'b1;
  assign \A[16][55] [1] = 1'b1;
  assign \A[16][55] [0] = 1'b1;
  assign \A[16][56] [4] = 1'b1;
  assign \A[16][56] [3] = 1'b1;
  assign \A[16][56] [2] = 1'b1;
  assign \A[16][56] [1] = 1'b1;
  assign \A[16][56] [0] = 1'b1;
  assign \A[16][57] [0] = 1'b1;
  assign \A[16][58] [4] = 1'b1;
  assign \A[16][58] [3] = 1'b1;
  assign \A[16][58] [2] = 1'b1;
  assign \A[16][58] [1] = 1'b1;
  assign \A[16][58] [0] = 1'b1;
  assign \A[16][59] [4] = 1'b1;
  assign \A[16][59] [3] = 1'b1;
  assign \A[16][59] [2] = 1'b1;
  assign \A[16][59] [1] = 1'b1;
  assign \A[16][59] [0] = 1'b1;
  assign \A[16][60] [0] = 1'b1;
  assign \A[16][61] [4] = 1'b1;
  assign \A[16][61] [3] = 1'b1;
  assign \A[16][61] [2] = 1'b1;
  assign \A[16][61] [1] = 1'b1;
  assign \A[16][61] [0] = 1'b1;
  assign \A[16][62] [4] = 1'b1;
  assign \A[16][62] [3] = 1'b1;
  assign \A[16][62] [2] = 1'b1;
  assign \A[16][62] [1] = 1'b1;
  assign \A[16][62] [0] = 1'b1;
  assign \A[16][63] [0] = 1'b1;
  assign \A[16][64] [0] = 1'b1;
  assign \A[16][65] [4] = 1'b1;
  assign \A[16][65] [3] = 1'b1;
  assign \A[16][65] [2] = 1'b1;
  assign \A[16][65] [1] = 1'b1;
  assign \A[16][66] [4] = 1'b1;
  assign \A[16][66] [3] = 1'b1;
  assign \A[16][66] [2] = 1'b1;
  assign \A[16][66] [1] = 1'b1;
  assign \A[16][67] [4] = 1'b1;
  assign \A[16][67] [3] = 1'b1;
  assign \A[16][67] [2] = 1'b1;
  assign \A[16][67] [1] = 1'b1;
  assign \A[16][67] [0] = 1'b1;
  assign \A[16][69] [4] = 1'b1;
  assign \A[16][69] [3] = 1'b1;
  assign \A[16][69] [2] = 1'b1;
  assign \A[16][69] [1] = 1'b1;
  assign \A[16][69] [0] = 1'b1;
  assign \A[16][71] [4] = 1'b1;
  assign \A[16][71] [3] = 1'b1;
  assign \A[16][71] [2] = 1'b1;
  assign \A[16][71] [1] = 1'b1;
  assign \A[16][71] [0] = 1'b1;
  assign \A[16][73] [4] = 1'b1;
  assign \A[16][73] [3] = 1'b1;
  assign \A[16][73] [2] = 1'b1;
  assign \A[16][73] [1] = 1'b1;
  assign \A[16][73] [0] = 1'b1;
  assign \A[16][74] [1] = 1'b1;
  assign \A[16][74] [0] = 1'b1;
  assign \A[16][76] [2] = 1'b1;
  assign \A[16][76] [0] = 1'b1;
  assign \A[16][77] [4] = 1'b1;
  assign \A[16][77] [3] = 1'b1;
  assign \A[16][77] [2] = 1'b1;
  assign \A[16][77] [1] = 1'b1;
  assign \A[16][77] [0] = 1'b1;
  assign \A[16][78] [0] = 1'b1;
  assign \A[16][79] [4] = 1'b1;
  assign \A[16][79] [3] = 1'b1;
  assign \A[16][79] [2] = 1'b1;
  assign \A[16][79] [1] = 1'b1;
  assign \A[16][79] [0] = 1'b1;
  assign \A[16][80] [4] = 1'b1;
  assign \A[16][80] [3] = 1'b1;
  assign \A[16][80] [2] = 1'b1;
  assign \A[16][80] [1] = 1'b1;
  assign \A[16][81] [0] = 1'b1;
  assign \A[16][82] [4] = 1'b1;
  assign \A[16][82] [3] = 1'b1;
  assign \A[16][82] [2] = 1'b1;
  assign \A[16][82] [1] = 1'b1;
  assign \A[16][82] [0] = 1'b1;
  assign \A[16][83] [4] = 1'b1;
  assign \A[16][83] [3] = 1'b1;
  assign \A[16][83] [2] = 1'b1;
  assign \A[16][83] [0] = 1'b1;
  assign \A[16][84] [4] = 1'b1;
  assign \A[16][84] [3] = 1'b1;
  assign \A[16][84] [2] = 1'b1;
  assign \A[16][84] [1] = 1'b1;
  assign \A[16][84] [0] = 1'b1;
  assign \A[16][85] [4] = 1'b1;
  assign \A[16][85] [3] = 1'b1;
  assign \A[16][85] [2] = 1'b1;
  assign \A[16][85] [0] = 1'b1;
  assign \A[16][86] [4] = 1'b1;
  assign \A[16][86] [3] = 1'b1;
  assign \A[16][86] [2] = 1'b1;
  assign \A[16][86] [1] = 1'b1;
  assign \A[16][86] [0] = 1'b1;
  assign \A[16][87] [1] = 1'b1;
  assign \A[16][88] [0] = 1'b1;
  assign \A[16][89] [4] = 1'b1;
  assign \A[16][89] [3] = 1'b1;
  assign \A[16][89] [2] = 1'b1;
  assign \A[16][89] [1] = 1'b1;
  assign \A[16][91] [4] = 1'b1;
  assign \A[16][91] [3] = 1'b1;
  assign \A[16][91] [2] = 1'b1;
  assign \A[16][91] [1] = 1'b1;
  assign \A[16][92] [1] = 1'b1;
  assign \A[16][93] [0] = 1'b1;
  assign \A[16][94] [4] = 1'b1;
  assign \A[16][94] [3] = 1'b1;
  assign \A[16][94] [2] = 1'b1;
  assign \A[16][94] [1] = 1'b1;
  assign \A[16][94] [0] = 1'b1;
  assign \A[16][96] [0] = 1'b1;
  assign \A[16][97] [0] = 1'b1;
  assign \A[16][99] [0] = 1'b1;
  assign \A[16][100] [0] = 1'b1;
  assign \A[16][101] [1] = 1'b1;
  assign \A[16][102] [4] = 1'b1;
  assign \A[16][102] [3] = 1'b1;
  assign \A[16][102] [2] = 1'b1;
  assign \A[16][103] [4] = 1'b1;
  assign \A[16][103] [3] = 1'b1;
  assign \A[16][103] [2] = 1'b1;
  assign \A[16][103] [1] = 1'b1;
  assign \A[16][103] [0] = 1'b1;
  assign \A[16][105] [0] = 1'b1;
  assign \A[16][106] [4] = 1'b1;
  assign \A[16][106] [3] = 1'b1;
  assign \A[16][106] [2] = 1'b1;
  assign \A[16][106] [1] = 1'b1;
  assign \A[16][107] [1] = 1'b1;
  assign \A[16][107] [0] = 1'b1;
  assign \A[16][108] [0] = 1'b1;
  assign \A[16][109] [0] = 1'b1;
  assign \A[16][110] [0] = 1'b1;
  assign \A[16][111] [4] = 1'b1;
  assign \A[16][111] [3] = 1'b1;
  assign \A[16][111] [2] = 1'b1;
  assign \A[16][111] [1] = 1'b1;
  assign \A[16][114] [4] = 1'b1;
  assign \A[16][114] [3] = 1'b1;
  assign \A[16][114] [2] = 1'b1;
  assign \A[16][114] [1] = 1'b1;
  assign \A[16][114] [0] = 1'b1;
  assign \A[16][115] [4] = 1'b1;
  assign \A[16][115] [3] = 1'b1;
  assign \A[16][115] [2] = 1'b1;
  assign \A[16][115] [1] = 1'b1;
  assign \A[16][115] [0] = 1'b1;
  assign \A[16][117] [1] = 1'b1;
  assign \A[16][118] [4] = 1'b1;
  assign \A[16][118] [3] = 1'b1;
  assign \A[16][118] [2] = 1'b1;
  assign \A[16][118] [1] = 1'b1;
  assign \A[16][120] [4] = 1'b1;
  assign \A[16][120] [3] = 1'b1;
  assign \A[16][120] [2] = 1'b1;
  assign \A[16][120] [1] = 1'b1;
  assign \A[16][120] [0] = 1'b1;
  assign \A[16][121] [0] = 1'b1;
  assign \A[16][123] [4] = 1'b1;
  assign \A[16][123] [3] = 1'b1;
  assign \A[16][123] [2] = 1'b1;
  assign \A[16][123] [1] = 1'b1;
  assign \A[16][123] [0] = 1'b1;
  assign \A[16][124] [1] = 1'b1;
  assign \A[16][124] [0] = 1'b1;
  assign \A[16][125] [0] = 1'b1;
  assign \A[16][126] [4] = 1'b1;
  assign \A[16][126] [3] = 1'b1;
  assign \A[16][126] [2] = 1'b1;
  assign \A[16][126] [1] = 1'b1;
  assign \A[16][127] [4] = 1'b1;
  assign \A[16][127] [3] = 1'b1;
  assign \A[16][127] [2] = 1'b1;
  assign \A[16][127] [1] = 1'b1;
  assign \A[16][127] [0] = 1'b1;
  assign \A[16][129] [1] = 1'b1;
  assign \A[16][130] [1] = 1'b1;
  assign \A[16][131] [4] = 1'b1;
  assign \A[16][131] [3] = 1'b1;
  assign \A[16][131] [2] = 1'b1;
  assign \A[16][131] [1] = 1'b1;
  assign \A[16][131] [0] = 1'b1;
  assign \A[16][132] [0] = 1'b1;
  assign \A[16][134] [0] = 1'b1;
  assign \A[16][135] [4] = 1'b1;
  assign \A[16][135] [3] = 1'b1;
  assign \A[16][135] [2] = 1'b1;
  assign \A[16][135] [1] = 1'b1;
  assign \A[16][139] [4] = 1'b1;
  assign \A[16][139] [3] = 1'b1;
  assign \A[16][139] [2] = 1'b1;
  assign \A[16][139] [1] = 1'b1;
  assign \A[16][140] [4] = 1'b1;
  assign \A[16][140] [3] = 1'b1;
  assign \A[16][140] [2] = 1'b1;
  assign \A[16][140] [1] = 1'b1;
  assign \A[16][140] [0] = 1'b1;
  assign \A[16][141] [4] = 1'b1;
  assign \A[16][141] [3] = 1'b1;
  assign \A[16][141] [2] = 1'b1;
  assign \A[16][141] [1] = 1'b1;
  assign \A[16][142] [4] = 1'b1;
  assign \A[16][142] [3] = 1'b1;
  assign \A[16][142] [2] = 1'b1;
  assign \A[16][142] [1] = 1'b1;
  assign \A[16][142] [0] = 1'b1;
  assign \A[16][143] [4] = 1'b1;
  assign \A[16][143] [3] = 1'b1;
  assign \A[16][143] [2] = 1'b1;
  assign \A[16][143] [1] = 1'b1;
  assign \A[16][143] [0] = 1'b1;
  assign \A[16][145] [0] = 1'b1;
  assign \A[16][147] [1] = 1'b1;
  assign \A[16][147] [0] = 1'b1;
  assign \A[16][150] [0] = 1'b1;
  assign \A[16][151] [4] = 1'b1;
  assign \A[16][151] [3] = 1'b1;
  assign \A[16][151] [2] = 1'b1;
  assign \A[16][151] [0] = 1'b1;
  assign \A[16][152] [0] = 1'b1;
  assign \A[16][153] [4] = 1'b1;
  assign \A[16][153] [3] = 1'b1;
  assign \A[16][153] [2] = 1'b1;
  assign \A[16][153] [1] = 1'b1;
  assign \A[16][155] [0] = 1'b1;
  assign \A[16][156] [4] = 1'b1;
  assign \A[16][156] [3] = 1'b1;
  assign \A[16][156] [2] = 1'b1;
  assign \A[16][156] [1] = 1'b1;
  assign \A[16][156] [0] = 1'b1;
  assign \A[16][157] [4] = 1'b1;
  assign \A[16][157] [3] = 1'b1;
  assign \A[16][157] [2] = 1'b1;
  assign \A[16][157] [1] = 1'b1;
  assign \A[16][158] [4] = 1'b1;
  assign \A[16][158] [3] = 1'b1;
  assign \A[16][158] [2] = 1'b1;
  assign \A[16][158] [1] = 1'b1;
  assign \A[16][158] [0] = 1'b1;
  assign \A[16][159] [4] = 1'b1;
  assign \A[16][159] [3] = 1'b1;
  assign \A[16][159] [2] = 1'b1;
  assign \A[16][159] [1] = 1'b1;
  assign \A[16][160] [1] = 1'b1;
  assign \A[16][162] [1] = 1'b1;
  assign \A[16][164] [1] = 1'b1;
  assign \A[16][165] [4] = 1'b1;
  assign \A[16][165] [3] = 1'b1;
  assign \A[16][165] [2] = 1'b1;
  assign \A[16][165] [1] = 1'b1;
  assign \A[16][165] [0] = 1'b1;
  assign \A[16][166] [4] = 1'b1;
  assign \A[16][166] [3] = 1'b1;
  assign \A[16][166] [2] = 1'b1;
  assign \A[16][166] [1] = 1'b1;
  assign \A[16][167] [1] = 1'b1;
  assign \A[16][168] [1] = 1'b1;
  assign \A[16][170] [1] = 1'b1;
  assign \A[16][171] [4] = 1'b1;
  assign \A[16][171] [3] = 1'b1;
  assign \A[16][171] [2] = 1'b1;
  assign \A[16][171] [1] = 1'b1;
  assign \A[16][171] [0] = 1'b1;
  assign \A[16][173] [4] = 1'b1;
  assign \A[16][173] [3] = 1'b1;
  assign \A[16][173] [2] = 1'b1;
  assign \A[16][173] [1] = 1'b1;
  assign \A[16][174] [4] = 1'b1;
  assign \A[16][174] [3] = 1'b1;
  assign \A[16][174] [2] = 1'b1;
  assign \A[16][174] [1] = 1'b1;
  assign \A[16][174] [0] = 1'b1;
  assign \A[16][175] [1] = 1'b1;
  assign \A[16][176] [0] = 1'b1;
  assign \A[16][177] [1] = 1'b1;
  assign \A[16][178] [4] = 1'b1;
  assign \A[16][178] [3] = 1'b1;
  assign \A[16][178] [2] = 1'b1;
  assign \A[16][178] [1] = 1'b1;
  assign \A[16][179] [0] = 1'b1;
  assign \A[16][181] [1] = 1'b1;
  assign \A[16][181] [0] = 1'b1;
  assign \A[16][182] [0] = 1'b1;
  assign \A[16][184] [4] = 1'b1;
  assign \A[16][184] [3] = 1'b1;
  assign \A[16][184] [2] = 1'b1;
  assign \A[16][184] [1] = 1'b1;
  assign \A[16][185] [4] = 1'b1;
  assign \A[16][185] [3] = 1'b1;
  assign \A[16][185] [2] = 1'b1;
  assign \A[16][185] [1] = 1'b1;
  assign \A[16][185] [0] = 1'b1;
  assign \A[16][186] [0] = 1'b1;
  assign \A[16][189] [4] = 1'b1;
  assign \A[16][189] [3] = 1'b1;
  assign \A[16][189] [2] = 1'b1;
  assign \A[16][189] [1] = 1'b1;
  assign \A[16][189] [0] = 1'b1;
  assign \A[16][190] [4] = 1'b1;
  assign \A[16][190] [3] = 1'b1;
  assign \A[16][190] [2] = 1'b1;
  assign \A[16][190] [1] = 1'b1;
  assign \A[16][191] [0] = 1'b1;
  assign \A[16][192] [4] = 1'b1;
  assign \A[16][192] [3] = 1'b1;
  assign \A[16][192] [2] = 1'b1;
  assign \A[16][192] [1] = 1'b1;
  assign \A[16][192] [0] = 1'b1;
  assign \A[16][194] [4] = 1'b1;
  assign \A[16][194] [3] = 1'b1;
  assign \A[16][194] [2] = 1'b1;
  assign \A[16][194] [1] = 1'b1;
  assign \A[16][195] [1] = 1'b1;
  assign \A[16][196] [4] = 1'b1;
  assign \A[16][196] [3] = 1'b1;
  assign \A[16][196] [2] = 1'b1;
  assign \A[16][196] [1] = 1'b1;
  assign \A[16][198] [4] = 1'b1;
  assign \A[16][198] [3] = 1'b1;
  assign \A[16][198] [2] = 1'b1;
  assign \A[16][198] [1] = 1'b1;
  assign \A[16][198] [0] = 1'b1;
  assign \A[16][199] [0] = 1'b1;
  assign \A[16][200] [4] = 1'b1;
  assign \A[16][200] [3] = 1'b1;
  assign \A[16][200] [2] = 1'b1;
  assign \A[16][200] [1] = 1'b1;
  assign \A[16][202] [4] = 1'b1;
  assign \A[16][202] [3] = 1'b1;
  assign \A[16][202] [2] = 1'b1;
  assign \A[16][202] [0] = 1'b1;
  assign \A[16][203] [4] = 1'b1;
  assign \A[16][203] [3] = 1'b1;
  assign \A[16][203] [2] = 1'b1;
  assign \A[16][203] [1] = 1'b1;
  assign \A[16][203] [0] = 1'b1;
  assign \A[16][204] [4] = 1'b1;
  assign \A[16][204] [3] = 1'b1;
  assign \A[16][204] [2] = 1'b1;
  assign \A[16][204] [1] = 1'b1;
  assign \A[16][205] [4] = 1'b1;
  assign \A[16][205] [3] = 1'b1;
  assign \A[16][205] [2] = 1'b1;
  assign \A[16][205] [1] = 1'b1;
  assign \A[16][205] [0] = 1'b1;
  assign \A[16][206] [4] = 1'b1;
  assign \A[16][206] [3] = 1'b1;
  assign \A[16][206] [2] = 1'b1;
  assign \A[16][206] [1] = 1'b1;
  assign \A[16][206] [0] = 1'b1;
  assign \A[16][209] [0] = 1'b1;
  assign \A[16][211] [1] = 1'b1;
  assign \A[16][212] [0] = 1'b1;
  assign \A[16][213] [4] = 1'b1;
  assign \A[16][213] [3] = 1'b1;
  assign \A[16][213] [2] = 1'b1;
  assign \A[16][213] [0] = 1'b1;
  assign \A[16][214] [1] = 1'b1;
  assign \A[16][215] [0] = 1'b1;
  assign \A[16][216] [4] = 1'b1;
  assign \A[16][216] [3] = 1'b1;
  assign \A[16][216] [2] = 1'b1;
  assign \A[16][216] [1] = 1'b1;
  assign \A[16][217] [4] = 1'b1;
  assign \A[16][217] [3] = 1'b1;
  assign \A[16][217] [2] = 1'b1;
  assign \A[16][217] [1] = 1'b1;
  assign \A[16][217] [0] = 1'b1;
  assign \A[16][218] [4] = 1'b1;
  assign \A[16][218] [3] = 1'b1;
  assign \A[16][218] [2] = 1'b1;
  assign \A[16][218] [1] = 1'b1;
  assign \A[16][220] [0] = 1'b1;
  assign \A[16][222] [4] = 1'b1;
  assign \A[16][222] [3] = 1'b1;
  assign \A[16][222] [2] = 1'b1;
  assign \A[16][222] [1] = 1'b1;
  assign \A[16][222] [0] = 1'b1;
  assign \A[16][223] [4] = 1'b1;
  assign \A[16][223] [3] = 1'b1;
  assign \A[16][223] [2] = 1'b1;
  assign \A[16][223] [1] = 1'b1;
  assign \A[16][230] [1] = 1'b1;
  assign \A[16][231] [0] = 1'b1;
  assign \A[16][233] [4] = 1'b1;
  assign \A[16][233] [3] = 1'b1;
  assign \A[16][233] [2] = 1'b1;
  assign \A[16][233] [1] = 1'b1;
  assign \A[16][234] [1] = 1'b1;
  assign \A[16][235] [4] = 1'b1;
  assign \A[16][235] [3] = 1'b1;
  assign \A[16][235] [2] = 1'b1;
  assign \A[16][235] [1] = 1'b1;
  assign \A[16][235] [0] = 1'b1;
  assign \A[16][236] [4] = 1'b1;
  assign \A[16][236] [3] = 1'b1;
  assign \A[16][236] [2] = 1'b1;
  assign \A[16][236] [1] = 1'b1;
  assign \A[16][236] [0] = 1'b1;
  assign \A[16][239] [4] = 1'b1;
  assign \A[16][239] [3] = 1'b1;
  assign \A[16][239] [2] = 1'b1;
  assign \A[16][239] [0] = 1'b1;
  assign \A[16][241] [4] = 1'b1;
  assign \A[16][241] [3] = 1'b1;
  assign \A[16][241] [2] = 1'b1;
  assign \A[16][241] [1] = 1'b1;
  assign \A[16][242] [4] = 1'b1;
  assign \A[16][242] [3] = 1'b1;
  assign \A[16][242] [2] = 1'b1;
  assign \A[16][242] [1] = 1'b1;
  assign \A[16][243] [4] = 1'b1;
  assign \A[16][243] [3] = 1'b1;
  assign \A[16][243] [2] = 1'b1;
  assign \A[16][243] [1] = 1'b1;
  assign \A[16][243] [0] = 1'b1;
  assign \A[16][244] [4] = 1'b1;
  assign \A[16][244] [3] = 1'b1;
  assign \A[16][244] [2] = 1'b1;
  assign \A[16][244] [1] = 1'b1;
  assign \A[16][244] [0] = 1'b1;
  assign \A[16][245] [4] = 1'b1;
  assign \A[16][245] [3] = 1'b1;
  assign \A[16][245] [2] = 1'b1;
  assign \A[16][245] [1] = 1'b1;
  assign \A[16][246] [0] = 1'b1;
  assign \A[16][247] [0] = 1'b1;
  assign \A[16][249] [1] = 1'b1;
  assign \A[16][251] [1] = 1'b1;
  assign \A[16][252] [1] = 1'b1;
  assign \A[16][253] [0] = 1'b1;
  assign \A[16][254] [0] = 1'b1;
  assign \A[17][0] [4] = 1'b1;
  assign \A[17][0] [3] = 1'b1;
  assign \A[17][0] [2] = 1'b1;
  assign \A[17][0] [1] = 1'b1;
  assign \A[17][0] [0] = 1'b1;
  assign \A[17][1] [4] = 1'b1;
  assign \A[17][1] [3] = 1'b1;
  assign \A[17][1] [2] = 1'b1;
  assign \A[17][1] [0] = 1'b1;
  assign \A[17][2] [1] = 1'b1;
  assign \A[17][3] [0] = 1'b1;
  assign \A[17][4] [4] = 1'b1;
  assign \A[17][4] [3] = 1'b1;
  assign \A[17][4] [2] = 1'b1;
  assign \A[17][4] [0] = 1'b1;
  assign \A[17][5] [4] = 1'b1;
  assign \A[17][5] [3] = 1'b1;
  assign \A[17][5] [2] = 1'b1;
  assign \A[17][6] [1] = 1'b1;
  assign \A[17][7] [2] = 1'b1;
  assign \A[17][7] [1] = 1'b1;
  assign \A[17][9] [4] = 1'b1;
  assign \A[17][9] [3] = 1'b1;
  assign \A[17][9] [2] = 1'b1;
  assign \A[17][9] [1] = 1'b1;
  assign \A[17][11] [4] = 1'b1;
  assign \A[17][11] [3] = 1'b1;
  assign \A[17][11] [2] = 1'b1;
  assign \A[17][11] [0] = 1'b1;
  assign \A[17][12] [4] = 1'b1;
  assign \A[17][12] [3] = 1'b1;
  assign \A[17][12] [2] = 1'b1;
  assign \A[17][12] [0] = 1'b1;
  assign \A[17][13] [4] = 1'b1;
  assign \A[17][13] [3] = 1'b1;
  assign \A[17][13] [2] = 1'b1;
  assign \A[17][13] [1] = 1'b1;
  assign \A[17][13] [0] = 1'b1;
  assign \A[17][14] [4] = 1'b1;
  assign \A[17][14] [3] = 1'b1;
  assign \A[17][14] [2] = 1'b1;
  assign \A[17][14] [1] = 1'b1;
  assign \A[17][15] [4] = 1'b1;
  assign \A[17][15] [3] = 1'b1;
  assign \A[17][15] [1] = 1'b1;
  assign \A[17][15] [0] = 1'b1;
  assign \A[17][18] [1] = 1'b1;
  assign \A[17][19] [4] = 1'b1;
  assign \A[17][19] [3] = 1'b1;
  assign \A[17][19] [2] = 1'b1;
  assign \A[17][19] [1] = 1'b1;
  assign \A[17][19] [0] = 1'b1;
  assign \A[17][21] [0] = 1'b1;
  assign \A[17][22] [1] = 1'b1;
  assign \A[17][23] [0] = 1'b1;
  assign \A[17][24] [4] = 1'b1;
  assign \A[17][24] [3] = 1'b1;
  assign \A[17][24] [2] = 1'b1;
  assign \A[17][24] [1] = 1'b1;
  assign \A[17][25] [0] = 1'b1;
  assign \A[17][26] [0] = 1'b1;
  assign \A[17][27] [1] = 1'b1;
  assign \A[17][28] [4] = 1'b1;
  assign \A[17][28] [3] = 1'b1;
  assign \A[17][28] [2] = 1'b1;
  assign \A[17][28] [1] = 1'b1;
  assign \A[17][29] [0] = 1'b1;
  assign \A[17][30] [1] = 1'b1;
  assign \A[17][31] [4] = 1'b1;
  assign \A[17][31] [3] = 1'b1;
  assign \A[17][31] [2] = 1'b1;
  assign \A[17][31] [1] = 1'b1;
  assign \A[17][31] [0] = 1'b1;
  assign \A[17][32] [4] = 1'b1;
  assign \A[17][32] [3] = 1'b1;
  assign \A[17][32] [2] = 1'b1;
  assign \A[17][32] [1] = 1'b1;
  assign \A[17][32] [0] = 1'b1;
  assign \A[17][33] [4] = 1'b1;
  assign \A[17][33] [3] = 1'b1;
  assign \A[17][33] [2] = 1'b1;
  assign \A[17][33] [1] = 1'b1;
  assign \A[17][33] [0] = 1'b1;
  assign \A[17][35] [4] = 1'b1;
  assign \A[17][35] [3] = 1'b1;
  assign \A[17][35] [2] = 1'b1;
  assign \A[17][35] [1] = 1'b1;
  assign \A[17][35] [0] = 1'b1;
  assign \A[17][36] [4] = 1'b1;
  assign \A[17][36] [3] = 1'b1;
  assign \A[17][36] [2] = 1'b1;
  assign \A[17][36] [1] = 1'b1;
  assign \A[17][37] [4] = 1'b1;
  assign \A[17][37] [3] = 1'b1;
  assign \A[17][37] [2] = 1'b1;
  assign \A[17][37] [1] = 1'b1;
  assign \A[17][37] [0] = 1'b1;
  assign \A[17][39] [4] = 1'b1;
  assign \A[17][39] [3] = 1'b1;
  assign \A[17][39] [2] = 1'b1;
  assign \A[17][39] [1] = 1'b1;
  assign \A[17][39] [0] = 1'b1;
  assign \A[17][41] [4] = 1'b1;
  assign \A[17][41] [3] = 1'b1;
  assign \A[17][41] [2] = 1'b1;
  assign \A[17][41] [1] = 1'b1;
  assign \A[17][41] [0] = 1'b1;
  assign \A[17][42] [1] = 1'b1;
  assign \A[17][43] [4] = 1'b1;
  assign \A[17][43] [3] = 1'b1;
  assign \A[17][43] [2] = 1'b1;
  assign \A[17][43] [1] = 1'b1;
  assign \A[17][44] [0] = 1'b1;
  assign \A[17][45] [4] = 1'b1;
  assign \A[17][45] [3] = 1'b1;
  assign \A[17][45] [2] = 1'b1;
  assign \A[17][45] [0] = 1'b1;
  assign \A[17][46] [0] = 1'b1;
  assign \A[17][47] [2] = 1'b1;
  assign \A[17][47] [0] = 1'b1;
  assign \A[17][48] [4] = 1'b1;
  assign \A[17][48] [3] = 1'b1;
  assign \A[17][48] [2] = 1'b1;
  assign \A[17][48] [1] = 1'b1;
  assign \A[17][48] [0] = 1'b1;
  assign \A[17][49] [4] = 1'b1;
  assign \A[17][49] [3] = 1'b1;
  assign \A[17][49] [2] = 1'b1;
  assign \A[17][49] [0] = 1'b1;
  assign \A[17][50] [0] = 1'b1;
  assign \A[17][51] [4] = 1'b1;
  assign \A[17][51] [3] = 1'b1;
  assign \A[17][51] [2] = 1'b1;
  assign \A[17][51] [1] = 1'b1;
  assign \A[17][52] [4] = 1'b1;
  assign \A[17][52] [3] = 1'b1;
  assign \A[17][52] [2] = 1'b1;
  assign \A[17][52] [1] = 1'b1;
  assign \A[17][53] [4] = 1'b1;
  assign \A[17][53] [3] = 1'b1;
  assign \A[17][53] [2] = 1'b1;
  assign \A[17][53] [1] = 1'b1;
  assign \A[17][54] [4] = 1'b1;
  assign \A[17][54] [3] = 1'b1;
  assign \A[17][54] [2] = 1'b1;
  assign \A[17][54] [1] = 1'b1;
  assign \A[17][54] [0] = 1'b1;
  assign \A[17][55] [2] = 1'b1;
  assign \A[17][57] [1] = 1'b1;
  assign \A[17][58] [4] = 1'b1;
  assign \A[17][58] [3] = 1'b1;
  assign \A[17][58] [2] = 1'b1;
  assign \A[17][58] [1] = 1'b1;
  assign \A[17][58] [0] = 1'b1;
  assign \A[17][59] [0] = 1'b1;
  assign \A[17][60] [0] = 1'b1;
  assign \A[17][61] [4] = 1'b1;
  assign \A[17][61] [3] = 1'b1;
  assign \A[17][61] [2] = 1'b1;
  assign \A[17][61] [1] = 1'b1;
  assign \A[17][61] [0] = 1'b1;
  assign \A[17][62] [1] = 1'b1;
  assign \A[17][63] [1] = 1'b1;
  assign \A[17][63] [0] = 1'b1;
  assign \A[17][65] [4] = 1'b1;
  assign \A[17][65] [3] = 1'b1;
  assign \A[17][65] [2] = 1'b1;
  assign \A[17][66] [4] = 1'b1;
  assign \A[17][66] [3] = 1'b1;
  assign \A[17][66] [2] = 1'b1;
  assign \A[17][66] [0] = 1'b1;
  assign \A[17][67] [1] = 1'b1;
  assign \A[17][69] [0] = 1'b1;
  assign \A[17][70] [0] = 1'b1;
  assign \A[17][71] [0] = 1'b1;
  assign \A[17][72] [4] = 1'b1;
  assign \A[17][72] [3] = 1'b1;
  assign \A[17][72] [2] = 1'b1;
  assign \A[17][72] [1] = 1'b1;
  assign \A[17][73] [4] = 1'b1;
  assign \A[17][73] [3] = 1'b1;
  assign \A[17][73] [2] = 1'b1;
  assign \A[17][73] [1] = 1'b1;
  assign \A[17][73] [0] = 1'b1;
  assign \A[17][74] [1] = 1'b1;
  assign \A[17][76] [2] = 1'b1;
  assign \A[17][76] [0] = 1'b1;
  assign \A[17][77] [4] = 1'b1;
  assign \A[17][77] [3] = 1'b1;
  assign \A[17][77] [2] = 1'b1;
  assign \A[17][77] [1] = 1'b1;
  assign \A[17][77] [0] = 1'b1;
  assign \A[17][78] [2] = 1'b1;
  assign \A[17][80] [4] = 1'b1;
  assign \A[17][80] [3] = 1'b1;
  assign \A[17][80] [2] = 1'b1;
  assign \A[17][80] [1] = 1'b1;
  assign \A[17][80] [0] = 1'b1;
  assign \A[17][81] [4] = 1'b1;
  assign \A[17][81] [3] = 1'b1;
  assign \A[17][81] [2] = 1'b1;
  assign \A[17][81] [1] = 1'b1;
  assign \A[17][83] [4] = 1'b1;
  assign \A[17][83] [3] = 1'b1;
  assign \A[17][83] [2] = 1'b1;
  assign \A[17][83] [1] = 1'b1;
  assign \A[17][83] [0] = 1'b1;
  assign \A[17][84] [4] = 1'b1;
  assign \A[17][84] [3] = 1'b1;
  assign \A[17][84] [2] = 1'b1;
  assign \A[17][84] [1] = 1'b1;
  assign \A[17][85] [0] = 1'b1;
  assign \A[17][86] [0] = 1'b1;
  assign \A[17][87] [4] = 1'b1;
  assign \A[17][87] [3] = 1'b1;
  assign \A[17][87] [2] = 1'b1;
  assign \A[17][87] [1] = 1'b1;
  assign \A[17][87] [0] = 1'b1;
  assign \A[17][88] [2] = 1'b1;
  assign \A[17][89] [0] = 1'b1;
  assign \A[17][92] [4] = 1'b1;
  assign \A[17][92] [3] = 1'b1;
  assign \A[17][92] [2] = 1'b1;
  assign \A[17][92] [1] = 1'b1;
  assign \A[17][93] [0] = 1'b1;
  assign \A[17][94] [4] = 1'b1;
  assign \A[17][94] [3] = 1'b1;
  assign \A[17][94] [2] = 1'b1;
  assign \A[17][94] [1] = 1'b1;
  assign \A[17][98] [1] = 1'b1;
  assign \A[17][99] [4] = 1'b1;
  assign \A[17][99] [3] = 1'b1;
  assign \A[17][99] [2] = 1'b1;
  assign \A[17][99] [1] = 1'b1;
  assign \A[17][100] [1] = 1'b1;
  assign \A[17][101] [4] = 1'b1;
  assign \A[17][101] [3] = 1'b1;
  assign \A[17][101] [2] = 1'b1;
  assign \A[17][101] [0] = 1'b1;
  assign \A[17][102] [4] = 1'b1;
  assign \A[17][102] [3] = 1'b1;
  assign \A[17][102] [2] = 1'b1;
  assign \A[17][102] [0] = 1'b1;
  assign \A[17][104] [1] = 1'b1;
  assign \A[17][105] [4] = 1'b1;
  assign \A[17][105] [3] = 1'b1;
  assign \A[17][105] [2] = 1'b1;
  assign \A[17][105] [1] = 1'b1;
  assign \A[17][105] [0] = 1'b1;
  assign \A[17][108] [1] = 1'b1;
  assign \A[17][109] [4] = 1'b1;
  assign \A[17][109] [3] = 1'b1;
  assign \A[17][109] [2] = 1'b1;
  assign \A[17][109] [1] = 1'b1;
  assign \A[17][110] [4] = 1'b1;
  assign \A[17][110] [3] = 1'b1;
  assign \A[17][110] [2] = 1'b1;
  assign \A[17][110] [1] = 1'b1;
  assign \A[17][112] [4] = 1'b1;
  assign \A[17][112] [3] = 1'b1;
  assign \A[17][112] [2] = 1'b1;
  assign \A[17][113] [4] = 1'b1;
  assign \A[17][113] [3] = 1'b1;
  assign \A[17][113] [2] = 1'b1;
  assign \A[17][113] [1] = 1'b1;
  assign \A[17][115] [4] = 1'b1;
  assign \A[17][115] [3] = 1'b1;
  assign \A[17][115] [2] = 1'b1;
  assign \A[17][115] [1] = 1'b1;
  assign \A[17][115] [0] = 1'b1;
  assign \A[17][117] [4] = 1'b1;
  assign \A[17][117] [3] = 1'b1;
  assign \A[17][117] [2] = 1'b1;
  assign \A[17][117] [1] = 1'b1;
  assign \A[17][118] [4] = 1'b1;
  assign \A[17][118] [3] = 1'b1;
  assign \A[17][118] [2] = 1'b1;
  assign \A[17][118] [1] = 1'b1;
  assign \A[17][118] [0] = 1'b1;
  assign \A[17][119] [1] = 1'b1;
  assign \A[17][120] [4] = 1'b1;
  assign \A[17][120] [3] = 1'b1;
  assign \A[17][120] [2] = 1'b1;
  assign \A[17][120] [0] = 1'b1;
  assign \A[17][121] [0] = 1'b1;
  assign \A[17][122] [4] = 1'b1;
  assign \A[17][122] [3] = 1'b1;
  assign \A[17][122] [2] = 1'b1;
  assign \A[17][122] [1] = 1'b1;
  assign \A[17][122] [0] = 1'b1;
  assign \A[17][124] [4] = 1'b1;
  assign \A[17][124] [3] = 1'b1;
  assign \A[17][124] [2] = 1'b1;
  assign \A[17][124] [1] = 1'b1;
  assign \A[17][124] [0] = 1'b1;
  assign \A[17][125] [4] = 1'b1;
  assign \A[17][125] [3] = 1'b1;
  assign \A[17][125] [2] = 1'b1;
  assign \A[17][125] [0] = 1'b1;
  assign \A[17][126] [4] = 1'b1;
  assign \A[17][126] [3] = 1'b1;
  assign \A[17][126] [2] = 1'b1;
  assign \A[17][126] [1] = 1'b1;
  assign \A[17][127] [4] = 1'b1;
  assign \A[17][127] [3] = 1'b1;
  assign \A[17][127] [2] = 1'b1;
  assign \A[17][127] [1] = 1'b1;
  assign \A[17][128] [4] = 1'b1;
  assign \A[17][128] [3] = 1'b1;
  assign \A[17][128] [2] = 1'b1;
  assign \A[17][128] [1] = 1'b1;
  assign \A[17][129] [4] = 1'b1;
  assign \A[17][129] [3] = 1'b1;
  assign \A[17][129] [2] = 1'b1;
  assign \A[17][129] [1] = 1'b1;
  assign \A[17][129] [0] = 1'b1;
  assign \A[17][130] [0] = 1'b1;
  assign \A[17][131] [0] = 1'b1;
  assign \A[17][132] [1] = 1'b1;
  assign \A[17][133] [4] = 1'b1;
  assign \A[17][133] [3] = 1'b1;
  assign \A[17][133] [2] = 1'b1;
  assign \A[17][133] [1] = 1'b1;
  assign \A[17][134] [4] = 1'b1;
  assign \A[17][134] [3] = 1'b1;
  assign \A[17][134] [2] = 1'b1;
  assign \A[17][134] [1] = 1'b1;
  assign \A[17][134] [0] = 1'b1;
  assign \A[17][136] [4] = 1'b1;
  assign \A[17][136] [3] = 1'b1;
  assign \A[17][136] [2] = 1'b1;
  assign \A[17][136] [1] = 1'b1;
  assign \A[17][136] [0] = 1'b1;
  assign \A[17][137] [1] = 1'b1;
  assign \A[17][139] [4] = 1'b1;
  assign \A[17][139] [3] = 1'b1;
  assign \A[17][139] [2] = 1'b1;
  assign \A[17][139] [1] = 1'b1;
  assign \A[17][140] [0] = 1'b1;
  assign \A[17][142] [4] = 1'b1;
  assign \A[17][142] [3] = 1'b1;
  assign \A[17][142] [2] = 1'b1;
  assign \A[17][142] [1] = 1'b1;
  assign \A[17][142] [0] = 1'b1;
  assign \A[17][143] [4] = 1'b1;
  assign \A[17][143] [3] = 1'b1;
  assign \A[17][143] [2] = 1'b1;
  assign \A[17][143] [1] = 1'b1;
  assign \A[17][145] [4] = 1'b1;
  assign \A[17][145] [3] = 1'b1;
  assign \A[17][145] [2] = 1'b1;
  assign \A[17][145] [1] = 1'b1;
  assign \A[17][146] [4] = 1'b1;
  assign \A[17][146] [3] = 1'b1;
  assign \A[17][146] [2] = 1'b1;
  assign \A[17][146] [1] = 1'b1;
  assign \A[17][146] [0] = 1'b1;
  assign \A[17][148] [4] = 1'b1;
  assign \A[17][148] [3] = 1'b1;
  assign \A[17][148] [1] = 1'b1;
  assign \A[17][148] [0] = 1'b1;
  assign \A[17][149] [4] = 1'b1;
  assign \A[17][149] [3] = 1'b1;
  assign \A[17][149] [2] = 1'b1;
  assign \A[17][149] [1] = 1'b1;
  assign \A[17][149] [0] = 1'b1;
  assign \A[17][150] [0] = 1'b1;
  assign \A[17][151] [1] = 1'b1;
  assign \A[17][152] [4] = 1'b1;
  assign \A[17][152] [3] = 1'b1;
  assign \A[17][152] [2] = 1'b1;
  assign \A[17][152] [1] = 1'b1;
  assign \A[17][153] [0] = 1'b1;
  assign \A[17][154] [4] = 1'b1;
  assign \A[17][154] [3] = 1'b1;
  assign \A[17][154] [2] = 1'b1;
  assign \A[17][154] [1] = 1'b1;
  assign \A[17][154] [0] = 1'b1;
  assign \A[17][156] [4] = 1'b1;
  assign \A[17][156] [3] = 1'b1;
  assign \A[17][156] [2] = 1'b1;
  assign \A[17][157] [0] = 1'b1;
  assign \A[17][158] [4] = 1'b1;
  assign \A[17][158] [3] = 1'b1;
  assign \A[17][158] [2] = 1'b1;
  assign \A[17][158] [1] = 1'b1;
  assign \A[17][159] [4] = 1'b1;
  assign \A[17][159] [3] = 1'b1;
  assign \A[17][159] [2] = 1'b1;
  assign \A[17][159] [1] = 1'b1;
  assign \A[17][159] [0] = 1'b1;
  assign \A[17][161] [0] = 1'b1;
  assign \A[17][162] [1] = 1'b1;
  assign \A[17][163] [1] = 1'b1;
  assign \A[17][163] [0] = 1'b1;
  assign \A[17][164] [0] = 1'b1;
  assign \A[17][165] [1] = 1'b1;
  assign \A[17][166] [4] = 1'b1;
  assign \A[17][166] [3] = 1'b1;
  assign \A[17][166] [2] = 1'b1;
  assign \A[17][166] [1] = 1'b1;
  assign \A[17][166] [0] = 1'b1;
  assign \A[17][168] [4] = 1'b1;
  assign \A[17][168] [3] = 1'b1;
  assign \A[17][168] [2] = 1'b1;
  assign \A[17][168] [1] = 1'b1;
  assign \A[17][169] [4] = 1'b1;
  assign \A[17][169] [3] = 1'b1;
  assign \A[17][169] [2] = 1'b1;
  assign \A[17][169] [1] = 1'b1;
  assign \A[17][169] [0] = 1'b1;
  assign \A[17][170] [0] = 1'b1;
  assign \A[17][171] [4] = 1'b1;
  assign \A[17][171] [3] = 1'b1;
  assign \A[17][171] [2] = 1'b1;
  assign \A[17][172] [4] = 1'b1;
  assign \A[17][172] [3] = 1'b1;
  assign \A[17][172] [2] = 1'b1;
  assign \A[17][172] [1] = 1'b1;
  assign \A[17][174] [0] = 1'b1;
  assign \A[17][175] [4] = 1'b1;
  assign \A[17][175] [3] = 1'b1;
  assign \A[17][175] [2] = 1'b1;
  assign \A[17][175] [1] = 1'b1;
  assign \A[17][175] [0] = 1'b1;
  assign \A[17][177] [4] = 1'b1;
  assign \A[17][177] [3] = 1'b1;
  assign \A[17][177] [2] = 1'b1;
  assign \A[17][177] [0] = 1'b1;
  assign \A[17][178] [0] = 1'b1;
  assign \A[17][180] [4] = 1'b1;
  assign \A[17][180] [3] = 1'b1;
  assign \A[17][180] [2] = 1'b1;
  assign \A[17][180] [1] = 1'b1;
  assign \A[17][180] [0] = 1'b1;
  assign \A[17][181] [0] = 1'b1;
  assign \A[17][182] [1] = 1'b1;
  assign \A[17][182] [0] = 1'b1;
  assign \A[17][183] [0] = 1'b1;
  assign \A[17][185] [4] = 1'b1;
  assign \A[17][185] [3] = 1'b1;
  assign \A[17][185] [2] = 1'b1;
  assign \A[17][185] [1] = 1'b1;
  assign \A[17][185] [0] = 1'b1;
  assign \A[17][186] [4] = 1'b1;
  assign \A[17][186] [3] = 1'b1;
  assign \A[17][186] [2] = 1'b1;
  assign \A[17][186] [0] = 1'b1;
  assign \A[17][187] [4] = 1'b1;
  assign \A[17][187] [3] = 1'b1;
  assign \A[17][187] [2] = 1'b1;
  assign \A[17][187] [1] = 1'b1;
  assign \A[17][187] [0] = 1'b1;
  assign \A[17][188] [4] = 1'b1;
  assign \A[17][188] [3] = 1'b1;
  assign \A[17][188] [2] = 1'b1;
  assign \A[17][188] [1] = 1'b1;
  assign \A[17][189] [0] = 1'b1;
  assign \A[17][191] [1] = 1'b1;
  assign \A[17][192] [0] = 1'b1;
  assign \A[17][194] [4] = 1'b1;
  assign \A[17][194] [3] = 1'b1;
  assign \A[17][194] [2] = 1'b1;
  assign \A[17][194] [1] = 1'b1;
  assign \A[17][194] [0] = 1'b1;
  assign \A[17][195] [0] = 1'b1;
  assign \A[17][196] [4] = 1'b1;
  assign \A[17][196] [3] = 1'b1;
  assign \A[17][196] [2] = 1'b1;
  assign \A[17][196] [1] = 1'b1;
  assign \A[17][196] [0] = 1'b1;
  assign \A[17][199] [4] = 1'b1;
  assign \A[17][199] [3] = 1'b1;
  assign \A[17][199] [2] = 1'b1;
  assign \A[17][199] [0] = 1'b1;
  assign \A[17][200] [4] = 1'b1;
  assign \A[17][200] [3] = 1'b1;
  assign \A[17][200] [2] = 1'b1;
  assign \A[17][200] [1] = 1'b1;
  assign \A[17][201] [4] = 1'b1;
  assign \A[17][201] [3] = 1'b1;
  assign \A[17][201] [2] = 1'b1;
  assign \A[17][201] [1] = 1'b1;
  assign \A[17][201] [0] = 1'b1;
  assign \A[17][203] [1] = 1'b1;
  assign \A[17][204] [1] = 1'b1;
  assign \A[17][207] [0] = 1'b1;
  assign \A[17][208] [2] = 1'b1;
  assign \A[17][208] [0] = 1'b1;
  assign \A[17][209] [4] = 1'b1;
  assign \A[17][209] [3] = 1'b1;
  assign \A[17][209] [2] = 1'b1;
  assign \A[17][209] [1] = 1'b1;
  assign \A[17][209] [0] = 1'b1;
  assign \A[17][211] [4] = 1'b1;
  assign \A[17][211] [3] = 1'b1;
  assign \A[17][211] [2] = 1'b1;
  assign \A[17][211] [1] = 1'b1;
  assign \A[17][211] [0] = 1'b1;
  assign \A[17][212] [1] = 1'b1;
  assign \A[17][213] [4] = 1'b1;
  assign \A[17][213] [3] = 1'b1;
  assign \A[17][213] [2] = 1'b1;
  assign \A[17][213] [1] = 1'b1;
  assign \A[17][215] [4] = 1'b1;
  assign \A[17][215] [3] = 1'b1;
  assign \A[17][215] [2] = 1'b1;
  assign \A[17][215] [1] = 1'b1;
  assign \A[17][215] [0] = 1'b1;
  assign \A[17][219] [1] = 1'b1;
  assign \A[17][219] [0] = 1'b1;
  assign \A[17][220] [4] = 1'b1;
  assign \A[17][220] [3] = 1'b1;
  assign \A[17][220] [2] = 1'b1;
  assign \A[17][220] [1] = 1'b1;
  assign \A[17][221] [0] = 1'b1;
  assign \A[17][222] [2] = 1'b1;
  assign \A[17][222] [0] = 1'b1;
  assign \A[17][223] [4] = 1'b1;
  assign \A[17][223] [3] = 1'b1;
  assign \A[17][223] [2] = 1'b1;
  assign \A[17][223] [1] = 1'b1;
  assign \A[17][223] [0] = 1'b1;
  assign \A[17][224] [0] = 1'b1;
  assign \A[17][225] [4] = 1'b1;
  assign \A[17][225] [3] = 1'b1;
  assign \A[17][225] [2] = 1'b1;
  assign \A[17][225] [1] = 1'b1;
  assign \A[17][229] [1] = 1'b1;
  assign \A[17][230] [4] = 1'b1;
  assign \A[17][230] [3] = 1'b1;
  assign \A[17][230] [2] = 1'b1;
  assign \A[17][230] [0] = 1'b1;
  assign \A[17][231] [0] = 1'b1;
  assign \A[17][232] [0] = 1'b1;
  assign \A[17][233] [1] = 1'b1;
  assign \A[17][234] [0] = 1'b1;
  assign \A[17][235] [1] = 1'b1;
  assign \A[17][236] [0] = 1'b1;
  assign \A[17][237] [2] = 1'b1;
  assign \A[17][238] [4] = 1'b1;
  assign \A[17][238] [3] = 1'b1;
  assign \A[17][238] [2] = 1'b1;
  assign \A[17][238] [1] = 1'b1;
  assign \A[17][239] [0] = 1'b1;
  assign \A[17][240] [1] = 1'b1;
  assign \A[17][241] [0] = 1'b1;
  assign \A[17][245] [4] = 1'b1;
  assign \A[17][245] [3] = 1'b1;
  assign \A[17][245] [2] = 1'b1;
  assign \A[17][245] [1] = 1'b1;
  assign \A[17][245] [0] = 1'b1;
  assign \A[17][246] [4] = 1'b1;
  assign \A[17][246] [3] = 1'b1;
  assign \A[17][246] [2] = 1'b1;
  assign \A[17][246] [1] = 1'b1;
  assign \A[17][248] [4] = 1'b1;
  assign \A[17][248] [3] = 1'b1;
  assign \A[17][248] [2] = 1'b1;
  assign \A[17][248] [1] = 1'b1;
  assign \A[17][249] [4] = 1'b1;
  assign \A[17][249] [3] = 1'b1;
  assign \A[17][249] [2] = 1'b1;
  assign \A[17][250] [1] = 1'b1;
  assign \A[17][251] [1] = 1'b1;
  assign \A[17][251] [0] = 1'b1;
  assign \A[17][252] [0] = 1'b1;
  assign \A[17][253] [1] = 1'b1;
  assign \A[17][254] [0] = 1'b1;
  assign \A[17][255] [4] = 1'b1;
  assign \A[17][255] [3] = 1'b1;
  assign \A[17][255] [2] = 1'b1;
  assign \A[17][255] [1] = 1'b1;
  assign \A[17][255] [0] = 1'b1;
  assign \A[18][0] [0] = 1'b1;
  assign \A[18][1] [1] = 1'b1;
  assign \A[18][1] [0] = 1'b1;
  assign \A[18][2] [0] = 1'b1;
  assign \A[18][3] [0] = 1'b1;
  assign \A[18][7] [4] = 1'b1;
  assign \A[18][7] [3] = 1'b1;
  assign \A[18][7] [2] = 1'b1;
  assign \A[18][7] [1] = 1'b1;
  assign \A[18][7] [0] = 1'b1;
  assign \A[18][9] [0] = 1'b1;
  assign \A[18][10] [1] = 1'b1;
  assign \A[18][12] [1] = 1'b1;
  assign \A[18][13] [4] = 1'b1;
  assign \A[18][13] [3] = 1'b1;
  assign \A[18][13] [2] = 1'b1;
  assign \A[18][13] [1] = 1'b1;
  assign \A[18][13] [0] = 1'b1;
  assign \A[18][14] [4] = 1'b1;
  assign \A[18][14] [3] = 1'b1;
  assign \A[18][14] [2] = 1'b1;
  assign \A[18][14] [1] = 1'b1;
  assign \A[18][15] [0] = 1'b1;
  assign \A[18][16] [4] = 1'b1;
  assign \A[18][16] [3] = 1'b1;
  assign \A[18][16] [2] = 1'b1;
  assign \A[18][16] [0] = 1'b1;
  assign \A[18][17] [1] = 1'b1;
  assign \A[18][18] [4] = 1'b1;
  assign \A[18][18] [3] = 1'b1;
  assign \A[18][18] [2] = 1'b1;
  assign \A[18][18] [1] = 1'b1;
  assign \A[18][18] [0] = 1'b1;
  assign \A[18][19] [1] = 1'b1;
  assign \A[18][21] [0] = 1'b1;
  assign \A[18][22] [4] = 1'b1;
  assign \A[18][22] [3] = 1'b1;
  assign \A[18][22] [2] = 1'b1;
  assign \A[18][22] [1] = 1'b1;
  assign \A[18][22] [0] = 1'b1;
  assign \A[18][24] [1] = 1'b1;
  assign \A[18][25] [1] = 1'b1;
  assign \A[18][25] [0] = 1'b1;
  assign \A[18][28] [4] = 1'b1;
  assign \A[18][28] [3] = 1'b1;
  assign \A[18][28] [2] = 1'b1;
  assign \A[18][28] [1] = 1'b1;
  assign \A[18][28] [0] = 1'b1;
  assign \A[18][30] [2] = 1'b1;
  assign \A[18][31] [4] = 1'b1;
  assign \A[18][31] [3] = 1'b1;
  assign \A[18][31] [2] = 1'b1;
  assign \A[18][31] [1] = 1'b1;
  assign \A[18][32] [4] = 1'b1;
  assign \A[18][32] [3] = 1'b1;
  assign \A[18][32] [2] = 1'b1;
  assign \A[18][32] [1] = 1'b1;
  assign \A[18][32] [0] = 1'b1;
  assign \A[18][33] [4] = 1'b1;
  assign \A[18][33] [3] = 1'b1;
  assign \A[18][33] [2] = 1'b1;
  assign \A[18][33] [0] = 1'b1;
  assign \A[18][34] [4] = 1'b1;
  assign \A[18][34] [3] = 1'b1;
  assign \A[18][34] [2] = 1'b1;
  assign \A[18][34] [1] = 1'b1;
  assign \A[18][34] [0] = 1'b1;
  assign \A[18][35] [4] = 1'b1;
  assign \A[18][35] [3] = 1'b1;
  assign \A[18][35] [2] = 1'b1;
  assign \A[18][35] [1] = 1'b1;
  assign \A[18][35] [0] = 1'b1;
  assign \A[18][36] [4] = 1'b1;
  assign \A[18][36] [3] = 1'b1;
  assign \A[18][36] [2] = 1'b1;
  assign \A[18][36] [1] = 1'b1;
  assign \A[18][37] [4] = 1'b1;
  assign \A[18][37] [3] = 1'b1;
  assign \A[18][37] [2] = 1'b1;
  assign \A[18][37] [0] = 1'b1;
  assign \A[18][40] [4] = 1'b1;
  assign \A[18][40] [3] = 1'b1;
  assign \A[18][40] [2] = 1'b1;
  assign \A[18][40] [1] = 1'b1;
  assign \A[18][40] [0] = 1'b1;
  assign \A[18][41] [4] = 1'b1;
  assign \A[18][41] [3] = 1'b1;
  assign \A[18][41] [2] = 1'b1;
  assign \A[18][41] [1] = 1'b1;
  assign \A[18][42] [1] = 1'b1;
  assign \A[18][43] [1] = 1'b1;
  assign \A[18][44] [0] = 1'b1;
  assign \A[18][45] [0] = 1'b1;
  assign \A[18][47] [2] = 1'b1;
  assign \A[18][48] [1] = 1'b1;
  assign \A[18][48] [0] = 1'b1;
  assign \A[18][50] [4] = 1'b1;
  assign \A[18][50] [3] = 1'b1;
  assign \A[18][50] [2] = 1'b1;
  assign \A[18][50] [1] = 1'b1;
  assign \A[18][51] [0] = 1'b1;
  assign \A[18][52] [4] = 1'b1;
  assign \A[18][52] [3] = 1'b1;
  assign \A[18][52] [2] = 1'b1;
  assign \A[18][52] [1] = 1'b1;
  assign \A[18][52] [0] = 1'b1;
  assign \A[18][54] [4] = 1'b1;
  assign \A[18][54] [3] = 1'b1;
  assign \A[18][54] [2] = 1'b1;
  assign \A[18][54] [1] = 1'b1;
  assign \A[18][55] [4] = 1'b1;
  assign \A[18][55] [3] = 1'b1;
  assign \A[18][55] [2] = 1'b1;
  assign \A[18][55] [1] = 1'b1;
  assign \A[18][55] [0] = 1'b1;
  assign \A[18][56] [0] = 1'b1;
  assign \A[18][57] [0] = 1'b1;
  assign \A[18][58] [2] = 1'b1;
  assign \A[18][60] [0] = 1'b1;
  assign \A[18][61] [0] = 1'b1;
  assign \A[18][62] [0] = 1'b1;
  assign \A[18][63] [0] = 1'b1;
  assign \A[18][64] [4] = 1'b1;
  assign \A[18][64] [3] = 1'b1;
  assign \A[18][64] [2] = 1'b1;
  assign \A[18][64] [1] = 1'b1;
  assign \A[18][65] [4] = 1'b1;
  assign \A[18][65] [3] = 1'b1;
  assign \A[18][65] [2] = 1'b1;
  assign \A[18][65] [1] = 1'b1;
  assign \A[18][65] [0] = 1'b1;
  assign \A[18][66] [4] = 1'b1;
  assign \A[18][66] [3] = 1'b1;
  assign \A[18][66] [2] = 1'b1;
  assign \A[18][68] [0] = 1'b1;
  assign \A[18][69] [0] = 1'b1;
  assign \A[18][71] [4] = 1'b1;
  assign \A[18][71] [3] = 1'b1;
  assign \A[18][71] [2] = 1'b1;
  assign \A[18][71] [1] = 1'b1;
  assign \A[18][71] [0] = 1'b1;
  assign \A[18][72] [4] = 1'b1;
  assign \A[18][72] [3] = 1'b1;
  assign \A[18][72] [2] = 1'b1;
  assign \A[18][72] [1] = 1'b1;
  assign \A[18][72] [0] = 1'b1;
  assign \A[18][73] [4] = 1'b1;
  assign \A[18][73] [3] = 1'b1;
  assign \A[18][73] [2] = 1'b1;
  assign \A[18][73] [1] = 1'b1;
  assign \A[18][75] [4] = 1'b1;
  assign \A[18][75] [3] = 1'b1;
  assign \A[18][75] [2] = 1'b1;
  assign \A[18][75] [1] = 1'b1;
  assign \A[18][75] [0] = 1'b1;
  assign \A[18][76] [0] = 1'b1;
  assign \A[18][77] [4] = 1'b1;
  assign \A[18][77] [3] = 1'b1;
  assign \A[18][77] [2] = 1'b1;
  assign \A[18][77] [1] = 1'b1;
  assign \A[18][77] [0] = 1'b1;
  assign \A[18][78] [1] = 1'b1;
  assign \A[18][79] [4] = 1'b1;
  assign \A[18][79] [3] = 1'b1;
  assign \A[18][79] [2] = 1'b1;
  assign \A[18][79] [1] = 1'b1;
  assign \A[18][79] [0] = 1'b1;
  assign \A[18][80] [0] = 1'b1;
  assign \A[18][81] [0] = 1'b1;
  assign \A[18][83] [4] = 1'b1;
  assign \A[18][83] [3] = 1'b1;
  assign \A[18][83] [2] = 1'b1;
  assign \A[18][83] [1] = 1'b1;
  assign \A[18][83] [0] = 1'b1;
  assign \A[18][84] [4] = 1'b1;
  assign \A[18][84] [3] = 1'b1;
  assign \A[18][84] [2] = 1'b1;
  assign \A[18][84] [1] = 1'b1;
  assign \A[18][84] [0] = 1'b1;
  assign \A[18][86] [0] = 1'b1;
  assign \A[18][88] [4] = 1'b1;
  assign \A[18][88] [3] = 1'b1;
  assign \A[18][88] [2] = 1'b1;
  assign \A[18][88] [1] = 1'b1;
  assign \A[18][89] [4] = 1'b1;
  assign \A[18][89] [3] = 1'b1;
  assign \A[18][89] [2] = 1'b1;
  assign \A[18][90] [4] = 1'b1;
  assign \A[18][90] [3] = 1'b1;
  assign \A[18][90] [2] = 1'b1;
  assign \A[18][90] [1] = 1'b1;
  assign \A[18][90] [0] = 1'b1;
  assign \A[18][91] [4] = 1'b1;
  assign \A[18][91] [3] = 1'b1;
  assign \A[18][91] [2] = 1'b1;
  assign \A[18][91] [0] = 1'b1;
  assign \A[18][92] [4] = 1'b1;
  assign \A[18][92] [3] = 1'b1;
  assign \A[18][92] [2] = 1'b1;
  assign \A[18][92] [1] = 1'b1;
  assign \A[18][93] [4] = 1'b1;
  assign \A[18][93] [3] = 1'b1;
  assign \A[18][93] [2] = 1'b1;
  assign \A[18][93] [1] = 1'b1;
  assign \A[18][95] [1] = 1'b1;
  assign \A[18][95] [0] = 1'b1;
  assign \A[18][96] [4] = 1'b1;
  assign \A[18][96] [3] = 1'b1;
  assign \A[18][96] [2] = 1'b1;
  assign \A[18][96] [1] = 1'b1;
  assign \A[18][96] [0] = 1'b1;
  assign \A[18][97] [0] = 1'b1;
  assign \A[18][98] [4] = 1'b1;
  assign \A[18][98] [3] = 1'b1;
  assign \A[18][98] [2] = 1'b1;
  assign \A[18][98] [1] = 1'b1;
  assign \A[18][98] [0] = 1'b1;
  assign \A[18][99] [4] = 1'b1;
  assign \A[18][99] [3] = 1'b1;
  assign \A[18][99] [2] = 1'b1;
  assign \A[18][99] [1] = 1'b1;
  assign \A[18][100] [4] = 1'b1;
  assign \A[18][100] [3] = 1'b1;
  assign \A[18][100] [2] = 1'b1;
  assign \A[18][100] [1] = 1'b1;
  assign \A[18][100] [0] = 1'b1;
  assign \A[18][103] [4] = 1'b1;
  assign \A[18][103] [3] = 1'b1;
  assign \A[18][103] [2] = 1'b1;
  assign \A[18][103] [0] = 1'b1;
  assign \A[18][104] [4] = 1'b1;
  assign \A[18][104] [3] = 1'b1;
  assign \A[18][104] [2] = 1'b1;
  assign \A[18][104] [1] = 1'b1;
  assign \A[18][105] [4] = 1'b1;
  assign \A[18][105] [3] = 1'b1;
  assign \A[18][105] [2] = 1'b1;
  assign \A[18][105] [1] = 1'b1;
  assign \A[18][106] [0] = 1'b1;
  assign \A[18][108] [4] = 1'b1;
  assign \A[18][108] [3] = 1'b1;
  assign \A[18][108] [2] = 1'b1;
  assign \A[18][108] [1] = 1'b1;
  assign \A[18][108] [0] = 1'b1;
  assign \A[18][110] [1] = 1'b1;
  assign \A[18][110] [0] = 1'b1;
  assign \A[18][111] [0] = 1'b1;
  assign \A[18][112] [1] = 1'b1;
  assign \A[18][112] [0] = 1'b1;
  assign \A[18][113] [0] = 1'b1;
  assign \A[18][114] [4] = 1'b1;
  assign \A[18][114] [3] = 1'b1;
  assign \A[18][114] [2] = 1'b1;
  assign \A[18][114] [1] = 1'b1;
  assign \A[18][116] [0] = 1'b1;
  assign \A[18][117] [4] = 1'b1;
  assign \A[18][117] [3] = 1'b1;
  assign \A[18][117] [2] = 1'b1;
  assign \A[18][117] [1] = 1'b1;
  assign \A[18][118] [4] = 1'b1;
  assign \A[18][118] [3] = 1'b1;
  assign \A[18][118] [2] = 1'b1;
  assign \A[18][118] [1] = 1'b1;
  assign \A[18][118] [0] = 1'b1;
  assign \A[18][122] [4] = 1'b1;
  assign \A[18][122] [3] = 1'b1;
  assign \A[18][122] [2] = 1'b1;
  assign \A[18][122] [0] = 1'b1;
  assign \A[18][123] [4] = 1'b1;
  assign \A[18][123] [3] = 1'b1;
  assign \A[18][123] [2] = 1'b1;
  assign \A[18][123] [1] = 1'b1;
  assign \A[18][124] [4] = 1'b1;
  assign \A[18][124] [3] = 1'b1;
  assign \A[18][124] [2] = 1'b1;
  assign \A[18][124] [1] = 1'b1;
  assign \A[18][125] [1] = 1'b1;
  assign \A[18][126] [2] = 1'b1;
  assign \A[18][126] [0] = 1'b1;
  assign \A[18][127] [4] = 1'b1;
  assign \A[18][127] [3] = 1'b1;
  assign \A[18][127] [2] = 1'b1;
  assign \A[18][127] [1] = 1'b1;
  assign \A[18][127] [0] = 1'b1;
  assign \A[18][128] [4] = 1'b1;
  assign \A[18][128] [3] = 1'b1;
  assign \A[18][128] [2] = 1'b1;
  assign \A[18][128] [1] = 1'b1;
  assign \A[18][128] [0] = 1'b1;
  assign \A[18][129] [1] = 1'b1;
  assign \A[18][129] [0] = 1'b1;
  assign \A[18][130] [0] = 1'b1;
  assign \A[18][131] [4] = 1'b1;
  assign \A[18][131] [3] = 1'b1;
  assign \A[18][131] [2] = 1'b1;
  assign \A[18][131] [0] = 1'b1;
  assign \A[18][132] [4] = 1'b1;
  assign \A[18][132] [3] = 1'b1;
  assign \A[18][132] [2] = 1'b1;
  assign \A[18][132] [0] = 1'b1;
  assign \A[18][133] [4] = 1'b1;
  assign \A[18][133] [3] = 1'b1;
  assign \A[18][133] [2] = 1'b1;
  assign \A[18][133] [1] = 1'b1;
  assign \A[18][133] [0] = 1'b1;
  assign \A[18][134] [4] = 1'b1;
  assign \A[18][134] [3] = 1'b1;
  assign \A[18][134] [2] = 1'b1;
  assign \A[18][134] [1] = 1'b1;
  assign \A[18][134] [0] = 1'b1;
  assign \A[18][135] [4] = 1'b1;
  assign \A[18][135] [3] = 1'b1;
  assign \A[18][135] [2] = 1'b1;
  assign \A[18][135] [1] = 1'b1;
  assign \A[18][135] [0] = 1'b1;
  assign \A[18][136] [0] = 1'b1;
  assign \A[18][137] [4] = 1'b1;
  assign \A[18][137] [3] = 1'b1;
  assign \A[18][137] [2] = 1'b1;
  assign \A[18][137] [1] = 1'b1;
  assign \A[18][137] [0] = 1'b1;
  assign \A[18][138] [4] = 1'b1;
  assign \A[18][138] [3] = 1'b1;
  assign \A[18][138] [2] = 1'b1;
  assign \A[18][138] [1] = 1'b1;
  assign \A[18][138] [0] = 1'b1;
  assign \A[18][139] [4] = 1'b1;
  assign \A[18][139] [3] = 1'b1;
  assign \A[18][139] [2] = 1'b1;
  assign \A[18][139] [1] = 1'b1;
  assign \A[18][139] [0] = 1'b1;
  assign \A[18][141] [4] = 1'b1;
  assign \A[18][141] [3] = 1'b1;
  assign \A[18][141] [2] = 1'b1;
  assign \A[18][141] [1] = 1'b1;
  assign \A[18][141] [0] = 1'b1;
  assign \A[18][142] [0] = 1'b1;
  assign \A[18][143] [0] = 1'b1;
  assign \A[18][144] [0] = 1'b1;
  assign \A[18][145] [0] = 1'b1;
  assign \A[18][146] [4] = 1'b1;
  assign \A[18][146] [3] = 1'b1;
  assign \A[18][146] [2] = 1'b1;
  assign \A[18][146] [1] = 1'b1;
  assign \A[18][146] [0] = 1'b1;
  assign \A[18][148] [0] = 1'b1;
  assign \A[18][149] [4] = 1'b1;
  assign \A[18][149] [3] = 1'b1;
  assign \A[18][149] [2] = 1'b1;
  assign \A[18][149] [1] = 1'b1;
  assign \A[18][149] [0] = 1'b1;
  assign \A[18][151] [4] = 1'b1;
  assign \A[18][151] [3] = 1'b1;
  assign \A[18][151] [2] = 1'b1;
  assign \A[18][151] [0] = 1'b1;
  assign \A[18][152] [4] = 1'b1;
  assign \A[18][152] [3] = 1'b1;
  assign \A[18][152] [2] = 1'b1;
  assign \A[18][152] [1] = 1'b1;
  assign \A[18][153] [1] = 1'b1;
  assign \A[18][153] [0] = 1'b1;
  assign \A[18][155] [1] = 1'b1;
  assign \A[18][156] [4] = 1'b1;
  assign \A[18][156] [3] = 1'b1;
  assign \A[18][156] [2] = 1'b1;
  assign \A[18][156] [1] = 1'b1;
  assign \A[18][156] [0] = 1'b1;
  assign \A[18][157] [0] = 1'b1;
  assign \A[18][158] [0] = 1'b1;
  assign \A[18][159] [2] = 1'b1;
  assign \A[18][160] [1] = 1'b1;
  assign \A[18][162] [1] = 1'b1;
  assign \A[18][163] [4] = 1'b1;
  assign \A[18][163] [3] = 1'b1;
  assign \A[18][163] [2] = 1'b1;
  assign \A[18][163] [1] = 1'b1;
  assign \A[18][165] [4] = 1'b1;
  assign \A[18][165] [3] = 1'b1;
  assign \A[18][165] [2] = 1'b1;
  assign \A[18][165] [0] = 1'b1;
  assign \A[18][166] [4] = 1'b1;
  assign \A[18][166] [3] = 1'b1;
  assign \A[18][166] [2] = 1'b1;
  assign \A[18][166] [1] = 1'b1;
  assign \A[18][166] [0] = 1'b1;
  assign \A[18][167] [4] = 1'b1;
  assign \A[18][167] [3] = 1'b1;
  assign \A[18][167] [2] = 1'b1;
  assign \A[18][167] [0] = 1'b1;
  assign \A[18][171] [4] = 1'b1;
  assign \A[18][171] [3] = 1'b1;
  assign \A[18][171] [2] = 1'b1;
  assign \A[18][171] [0] = 1'b1;
  assign \A[18][172] [4] = 1'b1;
  assign \A[18][172] [3] = 1'b1;
  assign \A[18][172] [2] = 1'b1;
  assign \A[18][172] [1] = 1'b1;
  assign \A[18][172] [0] = 1'b1;
  assign \A[18][173] [4] = 1'b1;
  assign \A[18][173] [3] = 1'b1;
  assign \A[18][173] [2] = 1'b1;
  assign \A[18][173] [1] = 1'b1;
  assign \A[18][173] [0] = 1'b1;
  assign \A[18][175] [0] = 1'b1;
  assign \A[18][176] [4] = 1'b1;
  assign \A[18][176] [3] = 1'b1;
  assign \A[18][176] [2] = 1'b1;
  assign \A[18][176] [1] = 1'b1;
  assign \A[18][176] [0] = 1'b1;
  assign \A[18][177] [4] = 1'b1;
  assign \A[18][177] [3] = 1'b1;
  assign \A[18][177] [2] = 1'b1;
  assign \A[18][177] [0] = 1'b1;
  assign \A[18][179] [0] = 1'b1;
  assign \A[18][180] [1] = 1'b1;
  assign \A[18][180] [0] = 1'b1;
  assign \A[18][181] [1] = 1'b1;
  assign \A[18][183] [4] = 1'b1;
  assign \A[18][183] [3] = 1'b1;
  assign \A[18][183] [2] = 1'b1;
  assign \A[18][183] [1] = 1'b1;
  assign \A[18][185] [1] = 1'b1;
  assign \A[18][186] [1] = 1'b1;
  assign \A[18][186] [0] = 1'b1;
  assign \A[18][188] [4] = 1'b1;
  assign \A[18][188] [3] = 1'b1;
  assign \A[18][188] [2] = 1'b1;
  assign \A[18][188] [1] = 1'b1;
  assign \A[18][188] [0] = 1'b1;
  assign \A[18][189] [4] = 1'b1;
  assign \A[18][189] [3] = 1'b1;
  assign \A[18][189] [2] = 1'b1;
  assign \A[18][189] [1] = 1'b1;
  assign \A[18][189] [0] = 1'b1;
  assign \A[18][190] [0] = 1'b1;
  assign \A[18][191] [4] = 1'b1;
  assign \A[18][191] [3] = 1'b1;
  assign \A[18][191] [2] = 1'b1;
  assign \A[18][191] [1] = 1'b1;
  assign \A[18][191] [0] = 1'b1;
  assign \A[18][192] [1] = 1'b1;
  assign \A[18][192] [0] = 1'b1;
  assign \A[18][194] [4] = 1'b1;
  assign \A[18][194] [3] = 1'b1;
  assign \A[18][194] [2] = 1'b1;
  assign \A[18][194] [1] = 1'b1;
  assign \A[18][194] [0] = 1'b1;
  assign \A[18][197] [0] = 1'b1;
  assign \A[18][198] [0] = 1'b1;
  assign \A[18][199] [0] = 1'b1;
  assign \A[18][201] [0] = 1'b1;
  assign \A[18][202] [0] = 1'b1;
  assign \A[18][203] [1] = 1'b1;
  assign \A[18][204] [1] = 1'b1;
  assign \A[18][205] [0] = 1'b1;
  assign \A[18][206] [4] = 1'b1;
  assign \A[18][206] [3] = 1'b1;
  assign \A[18][206] [2] = 1'b1;
  assign \A[18][206] [1] = 1'b1;
  assign \A[18][206] [0] = 1'b1;
  assign \A[18][207] [4] = 1'b1;
  assign \A[18][207] [3] = 1'b1;
  assign \A[18][207] [2] = 1'b1;
  assign \A[18][207] [1] = 1'b1;
  assign \A[18][207] [0] = 1'b1;
  assign \A[18][208] [0] = 1'b1;
  assign \A[18][209] [1] = 1'b1;
  assign \A[18][209] [0] = 1'b1;
  assign \A[18][210] [0] = 1'b1;
  assign \A[18][211] [1] = 1'b1;
  assign \A[18][212] [1] = 1'b1;
  assign \A[18][212] [0] = 1'b1;
  assign \A[18][214] [4] = 1'b1;
  assign \A[18][214] [3] = 1'b1;
  assign \A[18][214] [2] = 1'b1;
  assign \A[18][214] [1] = 1'b1;
  assign \A[18][214] [0] = 1'b1;
  assign \A[18][215] [1] = 1'b1;
  assign \A[18][215] [0] = 1'b1;
  assign \A[18][217] [4] = 1'b1;
  assign \A[18][217] [3] = 1'b1;
  assign \A[18][217] [2] = 1'b1;
  assign \A[18][217] [1] = 1'b1;
  assign \A[18][217] [0] = 1'b1;
  assign \A[18][219] [4] = 1'b1;
  assign \A[18][219] [3] = 1'b1;
  assign \A[18][219] [2] = 1'b1;
  assign \A[18][219] [1] = 1'b1;
  assign \A[18][221] [4] = 1'b1;
  assign \A[18][221] [3] = 1'b1;
  assign \A[18][221] [2] = 1'b1;
  assign \A[18][221] [1] = 1'b1;
  assign \A[18][221] [0] = 1'b1;
  assign \A[18][223] [4] = 1'b1;
  assign \A[18][223] [3] = 1'b1;
  assign \A[18][223] [2] = 1'b1;
  assign \A[18][223] [1] = 1'b1;
  assign \A[18][224] [1] = 1'b1;
  assign \A[18][225] [1] = 1'b1;
  assign \A[18][226] [0] = 1'b1;
  assign \A[18][228] [4] = 1'b1;
  assign \A[18][228] [3] = 1'b1;
  assign \A[18][228] [2] = 1'b1;
  assign \A[18][228] [1] = 1'b1;
  assign \A[18][228] [0] = 1'b1;
  assign \A[18][229] [1] = 1'b1;
  assign \A[18][230] [4] = 1'b1;
  assign \A[18][230] [3] = 1'b1;
  assign \A[18][230] [2] = 1'b1;
  assign \A[18][230] [1] = 1'b1;
  assign \A[18][230] [0] = 1'b1;
  assign \A[18][231] [1] = 1'b1;
  assign \A[18][231] [0] = 1'b1;
  assign \A[18][233] [1] = 1'b1;
  assign \A[18][235] [4] = 1'b1;
  assign \A[18][235] [3] = 1'b1;
  assign \A[18][235] [2] = 1'b1;
  assign \A[18][235] [1] = 1'b1;
  assign \A[18][237] [4] = 1'b1;
  assign \A[18][237] [3] = 1'b1;
  assign \A[18][237] [2] = 1'b1;
  assign \A[18][237] [1] = 1'b1;
  assign \A[18][238] [4] = 1'b1;
  assign \A[18][238] [3] = 1'b1;
  assign \A[18][238] [2] = 1'b1;
  assign \A[18][238] [1] = 1'b1;
  assign \A[18][238] [0] = 1'b1;
  assign \A[18][239] [4] = 1'b1;
  assign \A[18][239] [3] = 1'b1;
  assign \A[18][239] [2] = 1'b1;
  assign \A[18][239] [1] = 1'b1;
  assign \A[18][239] [0] = 1'b1;
  assign \A[18][240] [0] = 1'b1;
  assign \A[18][241] [1] = 1'b1;
  assign \A[18][242] [0] = 1'b1;
  assign \A[18][244] [4] = 1'b1;
  assign \A[18][244] [3] = 1'b1;
  assign \A[18][244] [2] = 1'b1;
  assign \A[18][244] [1] = 1'b1;
  assign \A[18][245] [4] = 1'b1;
  assign \A[18][245] [3] = 1'b1;
  assign \A[18][245] [2] = 1'b1;
  assign \A[18][245] [1] = 1'b1;
  assign \A[18][245] [0] = 1'b1;
  assign \A[18][246] [1] = 1'b1;
  assign \A[18][246] [0] = 1'b1;
  assign \A[18][247] [1] = 1'b1;
  assign \A[18][250] [4] = 1'b1;
  assign \A[18][250] [3] = 1'b1;
  assign \A[18][250] [2] = 1'b1;
  assign \A[18][250] [1] = 1'b1;
  assign \A[18][250] [0] = 1'b1;
  assign \A[18][251] [0] = 1'b1;
  assign \A[18][253] [4] = 1'b1;
  assign \A[18][253] [3] = 1'b1;
  assign \A[18][253] [2] = 1'b1;
  assign \A[18][253] [1] = 1'b1;
  assign \A[18][253] [0] = 1'b1;
  assign \A[18][254] [4] = 1'b1;
  assign \A[18][254] [3] = 1'b1;
  assign \A[18][254] [2] = 1'b1;
  assign \A[18][254] [1] = 1'b1;
  assign \A[18][254] [0] = 1'b1;
  assign \A[18][255] [0] = 1'b1;
  assign \A[19][0] [2] = 1'b1;
  assign \A[19][1] [4] = 1'b1;
  assign \A[19][1] [3] = 1'b1;
  assign \A[19][1] [2] = 1'b1;
  assign \A[19][1] [1] = 1'b1;
  assign \A[19][1] [0] = 1'b1;
  assign \A[19][2] [1] = 1'b1;
  assign \A[19][2] [0] = 1'b1;
  assign \A[19][3] [0] = 1'b1;
  assign \A[19][4] [4] = 1'b1;
  assign \A[19][4] [3] = 1'b1;
  assign \A[19][4] [2] = 1'b1;
  assign \A[19][4] [1] = 1'b1;
  assign \A[19][4] [0] = 1'b1;
  assign \A[19][5] [0] = 1'b1;
  assign \A[19][6] [2] = 1'b1;
  assign \A[19][7] [1] = 1'b1;
  assign \A[19][11] [1] = 1'b1;
  assign \A[19][12] [1] = 1'b1;
  assign \A[19][12] [0] = 1'b1;
  assign \A[19][13] [0] = 1'b1;
  assign \A[19][15] [2] = 1'b1;
  assign \A[19][16] [0] = 1'b1;
  assign \A[19][17] [4] = 1'b1;
  assign \A[19][17] [3] = 1'b1;
  assign \A[19][17] [2] = 1'b1;
  assign \A[19][17] [1] = 1'b1;
  assign \A[19][18] [0] = 1'b1;
  assign \A[19][19] [0] = 1'b1;
  assign \A[19][21] [1] = 1'b1;
  assign \A[19][22] [1] = 1'b1;
  assign \A[19][23] [4] = 1'b1;
  assign \A[19][23] [3] = 1'b1;
  assign \A[19][23] [2] = 1'b1;
  assign \A[19][23] [1] = 1'b1;
  assign \A[19][23] [0] = 1'b1;
  assign \A[19][24] [0] = 1'b1;
  assign \A[19][25] [1] = 1'b1;
  assign \A[19][26] [4] = 1'b1;
  assign \A[19][26] [3] = 1'b1;
  assign \A[19][26] [2] = 1'b1;
  assign \A[19][27] [1] = 1'b1;
  assign \A[19][28] [4] = 1'b1;
  assign \A[19][28] [3] = 1'b1;
  assign \A[19][28] [2] = 1'b1;
  assign \A[19][28] [1] = 1'b1;
  assign \A[19][28] [0] = 1'b1;
  assign \A[19][29] [4] = 1'b1;
  assign \A[19][29] [3] = 1'b1;
  assign \A[19][29] [2] = 1'b1;
  assign \A[19][29] [1] = 1'b1;
  assign \A[19][29] [0] = 1'b1;
  assign \A[19][30] [0] = 1'b1;
  assign \A[19][31] [4] = 1'b1;
  assign \A[19][31] [3] = 1'b1;
  assign \A[19][31] [2] = 1'b1;
  assign \A[19][31] [0] = 1'b1;
  assign \A[19][32] [0] = 1'b1;
  assign \A[19][33] [4] = 1'b1;
  assign \A[19][33] [3] = 1'b1;
  assign \A[19][33] [2] = 1'b1;
  assign \A[19][33] [1] = 1'b1;
  assign \A[19][33] [0] = 1'b1;
  assign \A[19][34] [4] = 1'b1;
  assign \A[19][34] [3] = 1'b1;
  assign \A[19][34] [2] = 1'b1;
  assign \A[19][34] [1] = 1'b1;
  assign \A[19][34] [0] = 1'b1;
  assign \A[19][36] [0] = 1'b1;
  assign \A[19][37] [4] = 1'b1;
  assign \A[19][37] [3] = 1'b1;
  assign \A[19][37] [2] = 1'b1;
  assign \A[19][37] [0] = 1'b1;
  assign \A[19][39] [2] = 1'b1;
  assign \A[19][41] [4] = 1'b1;
  assign \A[19][41] [3] = 1'b1;
  assign \A[19][41] [2] = 1'b1;
  assign \A[19][41] [1] = 1'b1;
  assign \A[19][41] [0] = 1'b1;
  assign \A[19][44] [4] = 1'b1;
  assign \A[19][44] [3] = 1'b1;
  assign \A[19][44] [2] = 1'b1;
  assign \A[19][44] [0] = 1'b1;
  assign \A[19][45] [1] = 1'b1;
  assign \A[19][46] [4] = 1'b1;
  assign \A[19][46] [3] = 1'b1;
  assign \A[19][46] [2] = 1'b1;
  assign \A[19][47] [4] = 1'b1;
  assign \A[19][47] [3] = 1'b1;
  assign \A[19][47] [2] = 1'b1;
  assign \A[19][47] [1] = 1'b1;
  assign \A[19][48] [4] = 1'b1;
  assign \A[19][48] [3] = 1'b1;
  assign \A[19][48] [2] = 1'b1;
  assign \A[19][48] [1] = 1'b1;
  assign \A[19][49] [4] = 1'b1;
  assign \A[19][49] [3] = 1'b1;
  assign \A[19][49] [2] = 1'b1;
  assign \A[19][49] [1] = 1'b1;
  assign \A[19][52] [4] = 1'b1;
  assign \A[19][52] [3] = 1'b1;
  assign \A[19][52] [2] = 1'b1;
  assign \A[19][52] [1] = 1'b1;
  assign \A[19][52] [0] = 1'b1;
  assign \A[19][54] [4] = 1'b1;
  assign \A[19][54] [3] = 1'b1;
  assign \A[19][54] [2] = 1'b1;
  assign \A[19][54] [1] = 1'b1;
  assign \A[19][56] [4] = 1'b1;
  assign \A[19][56] [3] = 1'b1;
  assign \A[19][56] [2] = 1'b1;
  assign \A[19][56] [0] = 1'b1;
  assign \A[19][57] [4] = 1'b1;
  assign \A[19][57] [3] = 1'b1;
  assign \A[19][57] [2] = 1'b1;
  assign \A[19][58] [4] = 1'b1;
  assign \A[19][58] [3] = 1'b1;
  assign \A[19][58] [2] = 1'b1;
  assign \A[19][58] [1] = 1'b1;
  assign \A[19][59] [4] = 1'b1;
  assign \A[19][59] [3] = 1'b1;
  assign \A[19][59] [1] = 1'b1;
  assign \A[19][60] [4] = 1'b1;
  assign \A[19][60] [3] = 1'b1;
  assign \A[19][60] [2] = 1'b1;
  assign \A[19][61] [4] = 1'b1;
  assign \A[19][61] [3] = 1'b1;
  assign \A[19][61] [2] = 1'b1;
  assign \A[19][61] [1] = 1'b1;
  assign \A[19][62] [4] = 1'b1;
  assign \A[19][62] [3] = 1'b1;
  assign \A[19][62] [2] = 1'b1;
  assign \A[19][62] [1] = 1'b1;
  assign \A[19][65] [4] = 1'b1;
  assign \A[19][65] [3] = 1'b1;
  assign \A[19][65] [2] = 1'b1;
  assign \A[19][65] [1] = 1'b1;
  assign \A[19][65] [0] = 1'b1;
  assign \A[19][66] [4] = 1'b1;
  assign \A[19][66] [3] = 1'b1;
  assign \A[19][66] [2] = 1'b1;
  assign \A[19][66] [1] = 1'b1;
  assign \A[19][66] [0] = 1'b1;
  assign \A[19][68] [4] = 1'b1;
  assign \A[19][68] [3] = 1'b1;
  assign \A[19][68] [2] = 1'b1;
  assign \A[19][68] [1] = 1'b1;
  assign \A[19][68] [0] = 1'b1;
  assign \A[19][69] [4] = 1'b1;
  assign \A[19][69] [3] = 1'b1;
  assign \A[19][69] [2] = 1'b1;
  assign \A[19][69] [1] = 1'b1;
  assign \A[19][69] [0] = 1'b1;
  assign \A[19][70] [4] = 1'b1;
  assign \A[19][70] [3] = 1'b1;
  assign \A[19][70] [2] = 1'b1;
  assign \A[19][70] [1] = 1'b1;
  assign \A[19][70] [0] = 1'b1;
  assign \A[19][71] [4] = 1'b1;
  assign \A[19][71] [3] = 1'b1;
  assign \A[19][71] [2] = 1'b1;
  assign \A[19][71] [1] = 1'b1;
  assign \A[19][71] [0] = 1'b1;
  assign \A[19][72] [4] = 1'b1;
  assign \A[19][72] [3] = 1'b1;
  assign \A[19][72] [2] = 1'b1;
  assign \A[19][72] [1] = 1'b1;
  assign \A[19][72] [0] = 1'b1;
  assign \A[19][73] [4] = 1'b1;
  assign \A[19][73] [3] = 1'b1;
  assign \A[19][73] [2] = 1'b1;
  assign \A[19][73] [0] = 1'b1;
  assign \A[19][74] [1] = 1'b1;
  assign \A[19][75] [4] = 1'b1;
  assign \A[19][75] [3] = 1'b1;
  assign \A[19][75] [2] = 1'b1;
  assign \A[19][75] [1] = 1'b1;
  assign \A[19][75] [0] = 1'b1;
  assign \A[19][76] [4] = 1'b1;
  assign \A[19][76] [3] = 1'b1;
  assign \A[19][76] [2] = 1'b1;
  assign \A[19][76] [0] = 1'b1;
  assign \A[19][77] [4] = 1'b1;
  assign \A[19][77] [3] = 1'b1;
  assign \A[19][77] [1] = 1'b1;
  assign \A[19][77] [0] = 1'b1;
  assign \A[19][78] [4] = 1'b1;
  assign \A[19][78] [3] = 1'b1;
  assign \A[19][78] [0] = 1'b1;
  assign \A[19][79] [4] = 1'b1;
  assign \A[19][79] [3] = 1'b1;
  assign \A[19][79] [1] = 1'b1;
  assign \A[19][79] [0] = 1'b1;
  assign \A[19][80] [4] = 1'b1;
  assign \A[19][80] [3] = 1'b1;
  assign \A[19][80] [2] = 1'b1;
  assign \A[19][80] [1] = 1'b1;
  assign \A[19][81] [4] = 1'b1;
  assign \A[19][81] [3] = 1'b1;
  assign \A[19][81] [2] = 1'b1;
  assign \A[19][81] [1] = 1'b1;
  assign \A[19][81] [0] = 1'b1;
  assign \A[19][82] [4] = 1'b1;
  assign \A[19][82] [3] = 1'b1;
  assign \A[19][82] [2] = 1'b1;
  assign \A[19][83] [4] = 1'b1;
  assign \A[19][83] [3] = 1'b1;
  assign \A[19][83] [2] = 1'b1;
  assign \A[19][83] [1] = 1'b1;
  assign \A[19][84] [0] = 1'b1;
  assign \A[19][85] [4] = 1'b1;
  assign \A[19][85] [3] = 1'b1;
  assign \A[19][85] [2] = 1'b1;
  assign \A[19][85] [1] = 1'b1;
  assign \A[19][85] [0] = 1'b1;
  assign \A[19][86] [1] = 1'b1;
  assign \A[19][87] [4] = 1'b1;
  assign \A[19][87] [3] = 1'b1;
  assign \A[19][87] [1] = 1'b1;
  assign \A[19][87] [0] = 1'b1;
  assign \A[19][88] [4] = 1'b1;
  assign \A[19][88] [3] = 1'b1;
  assign \A[19][88] [2] = 1'b1;
  assign \A[19][88] [1] = 1'b1;
  assign \A[19][88] [0] = 1'b1;
  assign \A[19][90] [4] = 1'b1;
  assign \A[19][90] [3] = 1'b1;
  assign \A[19][90] [2] = 1'b1;
  assign \A[19][90] [1] = 1'b1;
  assign \A[19][90] [0] = 1'b1;
  assign \A[19][91] [4] = 1'b1;
  assign \A[19][91] [3] = 1'b1;
  assign \A[19][91] [2] = 1'b1;
  assign \A[19][91] [1] = 1'b1;
  assign \A[19][92] [4] = 1'b1;
  assign \A[19][92] [3] = 1'b1;
  assign \A[19][92] [2] = 1'b1;
  assign \A[19][92] [1] = 1'b1;
  assign \A[19][92] [0] = 1'b1;
  assign \A[19][93] [4] = 1'b1;
  assign \A[19][93] [3] = 1'b1;
  assign \A[19][93] [2] = 1'b1;
  assign \A[19][93] [1] = 1'b1;
  assign \A[19][94] [4] = 1'b1;
  assign \A[19][94] [3] = 1'b1;
  assign \A[19][95] [4] = 1'b1;
  assign \A[19][95] [3] = 1'b1;
  assign \A[19][95] [2] = 1'b1;
  assign \A[19][96] [4] = 1'b1;
  assign \A[19][96] [3] = 1'b1;
  assign \A[19][96] [2] = 1'b1;
  assign \A[19][96] [1] = 1'b1;
  assign \A[19][96] [0] = 1'b1;
  assign \A[19][97] [0] = 1'b1;
  assign \A[19][100] [4] = 1'b1;
  assign \A[19][100] [3] = 1'b1;
  assign \A[19][100] [2] = 1'b1;
  assign \A[19][100] [1] = 1'b1;
  assign \A[19][102] [4] = 1'b1;
  assign \A[19][102] [3] = 1'b1;
  assign \A[19][102] [2] = 1'b1;
  assign \A[19][102] [1] = 1'b1;
  assign \A[19][102] [0] = 1'b1;
  assign \A[19][104] [4] = 1'b1;
  assign \A[19][104] [3] = 1'b1;
  assign \A[19][104] [2] = 1'b1;
  assign \A[19][104] [1] = 1'b1;
  assign \A[19][104] [0] = 1'b1;
  assign \A[19][106] [4] = 1'b1;
  assign \A[19][106] [3] = 1'b1;
  assign \A[19][106] [2] = 1'b1;
  assign \A[19][106] [1] = 1'b1;
  assign \A[19][106] [0] = 1'b1;
  assign \A[19][108] [4] = 1'b1;
  assign \A[19][108] [3] = 1'b1;
  assign \A[19][108] [2] = 1'b1;
  assign \A[19][108] [1] = 1'b1;
  assign \A[19][108] [0] = 1'b1;
  assign \A[19][110] [4] = 1'b1;
  assign \A[19][110] [3] = 1'b1;
  assign \A[19][110] [2] = 1'b1;
  assign \A[19][111] [4] = 1'b1;
  assign \A[19][111] [3] = 1'b1;
  assign \A[19][111] [0] = 1'b1;
  assign \A[19][114] [0] = 1'b1;
  assign \A[19][115] [4] = 1'b1;
  assign \A[19][115] [3] = 1'b1;
  assign \A[19][115] [2] = 1'b1;
  assign \A[19][115] [1] = 1'b1;
  assign \A[19][115] [0] = 1'b1;
  assign \A[19][117] [0] = 1'b1;
  assign \A[19][118] [4] = 1'b1;
  assign \A[19][118] [3] = 1'b1;
  assign \A[19][118] [2] = 1'b1;
  assign \A[19][118] [1] = 1'b1;
  assign \A[19][118] [0] = 1'b1;
  assign \A[19][119] [4] = 1'b1;
  assign \A[19][119] [3] = 1'b1;
  assign \A[19][119] [2] = 1'b1;
  assign \A[19][119] [1] = 1'b1;
  assign \A[19][120] [4] = 1'b1;
  assign \A[19][120] [3] = 1'b1;
  assign \A[19][120] [2] = 1'b1;
  assign \A[19][120] [1] = 1'b1;
  assign \A[19][123] [4] = 1'b1;
  assign \A[19][123] [3] = 1'b1;
  assign \A[19][123] [2] = 1'b1;
  assign \A[19][123] [1] = 1'b1;
  assign \A[19][123] [0] = 1'b1;
  assign \A[19][125] [0] = 1'b1;
  assign \A[19][127] [4] = 1'b1;
  assign \A[19][127] [3] = 1'b1;
  assign \A[19][127] [2] = 1'b1;
  assign \A[19][127] [1] = 1'b1;
  assign \A[19][127] [0] = 1'b1;
  assign \A[19][128] [4] = 1'b1;
  assign \A[19][128] [3] = 1'b1;
  assign \A[19][128] [2] = 1'b1;
  assign \A[19][128] [0] = 1'b1;
  assign \A[19][130] [0] = 1'b1;
  assign \A[19][131] [0] = 1'b1;
  assign \A[19][132] [4] = 1'b1;
  assign \A[19][132] [3] = 1'b1;
  assign \A[19][132] [2] = 1'b1;
  assign \A[19][132] [1] = 1'b1;
  assign \A[19][133] [4] = 1'b1;
  assign \A[19][133] [3] = 1'b1;
  assign \A[19][133] [2] = 1'b1;
  assign \A[19][133] [1] = 1'b1;
  assign \A[19][133] [0] = 1'b1;
  assign \A[19][134] [4] = 1'b1;
  assign \A[19][134] [3] = 1'b1;
  assign \A[19][134] [2] = 1'b1;
  assign \A[19][134] [1] = 1'b1;
  assign \A[19][136] [4] = 1'b1;
  assign \A[19][136] [3] = 1'b1;
  assign \A[19][136] [2] = 1'b1;
  assign \A[19][136] [1] = 1'b1;
  assign \A[19][138] [1] = 1'b1;
  assign \A[19][138] [0] = 1'b1;
  assign \A[19][139] [4] = 1'b1;
  assign \A[19][139] [3] = 1'b1;
  assign \A[19][139] [2] = 1'b1;
  assign \A[19][139] [1] = 1'b1;
  assign \A[19][139] [0] = 1'b1;
  assign \A[19][140] [0] = 1'b1;
  assign \A[19][141] [4] = 1'b1;
  assign \A[19][141] [3] = 1'b1;
  assign \A[19][141] [2] = 1'b1;
  assign \A[19][141] [1] = 1'b1;
  assign \A[19][141] [0] = 1'b1;
  assign \A[19][143] [4] = 1'b1;
  assign \A[19][143] [3] = 1'b1;
  assign \A[19][143] [2] = 1'b1;
  assign \A[19][143] [1] = 1'b1;
  assign \A[19][143] [0] = 1'b1;
  assign \A[19][144] [4] = 1'b1;
  assign \A[19][144] [3] = 1'b1;
  assign \A[19][144] [1] = 1'b1;
  assign \A[19][144] [0] = 1'b1;
  assign \A[19][145] [4] = 1'b1;
  assign \A[19][145] [3] = 1'b1;
  assign \A[19][145] [2] = 1'b1;
  assign \A[19][145] [0] = 1'b1;
  assign \A[19][146] [0] = 1'b1;
  assign \A[19][147] [4] = 1'b1;
  assign \A[19][147] [3] = 1'b1;
  assign \A[19][147] [2] = 1'b1;
  assign \A[19][147] [1] = 1'b1;
  assign \A[19][150] [0] = 1'b1;
  assign \A[19][151] [4] = 1'b1;
  assign \A[19][151] [3] = 1'b1;
  assign \A[19][151] [2] = 1'b1;
  assign \A[19][151] [1] = 1'b1;
  assign \A[19][151] [0] = 1'b1;
  assign \A[19][152] [4] = 1'b1;
  assign \A[19][152] [3] = 1'b1;
  assign \A[19][152] [2] = 1'b1;
  assign \A[19][152] [1] = 1'b1;
  assign \A[19][152] [0] = 1'b1;
  assign \A[19][154] [4] = 1'b1;
  assign \A[19][154] [3] = 1'b1;
  assign \A[19][154] [2] = 1'b1;
  assign \A[19][154] [1] = 1'b1;
  assign \A[19][154] [0] = 1'b1;
  assign \A[19][155] [4] = 1'b1;
  assign \A[19][155] [3] = 1'b1;
  assign \A[19][155] [2] = 1'b1;
  assign \A[19][155] [1] = 1'b1;
  assign \A[19][155] [0] = 1'b1;
  assign \A[19][157] [4] = 1'b1;
  assign \A[19][157] [3] = 1'b1;
  assign \A[19][157] [2] = 1'b1;
  assign \A[19][157] [1] = 1'b1;
  assign \A[19][157] [0] = 1'b1;
  assign \A[19][160] [4] = 1'b1;
  assign \A[19][160] [3] = 1'b1;
  assign \A[19][160] [2] = 1'b1;
  assign \A[19][160] [1] = 1'b1;
  assign \A[19][161] [4] = 1'b1;
  assign \A[19][161] [3] = 1'b1;
  assign \A[19][161] [2] = 1'b1;
  assign \A[19][161] [1] = 1'b1;
  assign \A[19][162] [4] = 1'b1;
  assign \A[19][162] [3] = 1'b1;
  assign \A[19][162] [2] = 1'b1;
  assign \A[19][162] [1] = 1'b1;
  assign \A[19][162] [0] = 1'b1;
  assign \A[19][165] [0] = 1'b1;
  assign \A[19][168] [4] = 1'b1;
  assign \A[19][168] [3] = 1'b1;
  assign \A[19][168] [2] = 1'b1;
  assign \A[19][168] [1] = 1'b1;
  assign \A[19][168] [0] = 1'b1;
  assign \A[19][170] [0] = 1'b1;
  assign \A[19][173] [4] = 1'b1;
  assign \A[19][173] [3] = 1'b1;
  assign \A[19][173] [2] = 1'b1;
  assign \A[19][173] [0] = 1'b1;
  assign \A[19][174] [4] = 1'b1;
  assign \A[19][174] [3] = 1'b1;
  assign \A[19][174] [2] = 1'b1;
  assign \A[19][174] [1] = 1'b1;
  assign \A[19][176] [4] = 1'b1;
  assign \A[19][176] [3] = 1'b1;
  assign \A[19][176] [2] = 1'b1;
  assign \A[19][176] [1] = 1'b1;
  assign \A[19][178] [4] = 1'b1;
  assign \A[19][178] [3] = 1'b1;
  assign \A[19][178] [2] = 1'b1;
  assign \A[19][178] [1] = 1'b1;
  assign \A[19][179] [4] = 1'b1;
  assign \A[19][179] [3] = 1'b1;
  assign \A[19][179] [2] = 1'b1;
  assign \A[19][179] [1] = 1'b1;
  assign \A[19][181] [4] = 1'b1;
  assign \A[19][181] [3] = 1'b1;
  assign \A[19][181] [2] = 1'b1;
  assign \A[19][181] [1] = 1'b1;
  assign \A[19][181] [0] = 1'b1;
  assign \A[19][182] [4] = 1'b1;
  assign \A[19][182] [3] = 1'b1;
  assign \A[19][182] [2] = 1'b1;
  assign \A[19][182] [1] = 1'b1;
  assign \A[19][182] [0] = 1'b1;
  assign \A[19][183] [4] = 1'b1;
  assign \A[19][183] [3] = 1'b1;
  assign \A[19][183] [2] = 1'b1;
  assign \A[19][183] [1] = 1'b1;
  assign \A[19][183] [0] = 1'b1;
  assign \A[19][184] [4] = 1'b1;
  assign \A[19][184] [3] = 1'b1;
  assign \A[19][184] [2] = 1'b1;
  assign \A[19][184] [0] = 1'b1;
  assign \A[19][187] [1] = 1'b1;
  assign \A[19][188] [4] = 1'b1;
  assign \A[19][188] [3] = 1'b1;
  assign \A[19][188] [2] = 1'b1;
  assign \A[19][188] [1] = 1'b1;
  assign \A[19][189] [0] = 1'b1;
  assign \A[19][190] [1] = 1'b1;
  assign \A[19][191] [1] = 1'b1;
  assign \A[19][192] [1] = 1'b1;
  assign \A[19][193] [0] = 1'b1;
  assign \A[19][195] [4] = 1'b1;
  assign \A[19][195] [3] = 1'b1;
  assign \A[19][195] [2] = 1'b1;
  assign \A[19][195] [0] = 1'b1;
  assign \A[19][197] [4] = 1'b1;
  assign \A[19][197] [3] = 1'b1;
  assign \A[19][197] [2] = 1'b1;
  assign \A[19][197] [1] = 1'b1;
  assign \A[19][197] [0] = 1'b1;
  assign \A[19][198] [1] = 1'b1;
  assign \A[19][199] [4] = 1'b1;
  assign \A[19][199] [3] = 1'b1;
  assign \A[19][199] [2] = 1'b1;
  assign \A[19][199] [1] = 1'b1;
  assign \A[19][199] [0] = 1'b1;
  assign \A[19][201] [4] = 1'b1;
  assign \A[19][201] [3] = 1'b1;
  assign \A[19][201] [2] = 1'b1;
  assign \A[19][202] [4] = 1'b1;
  assign \A[19][202] [3] = 1'b1;
  assign \A[19][202] [2] = 1'b1;
  assign \A[19][202] [1] = 1'b1;
  assign \A[19][204] [0] = 1'b1;
  assign \A[19][205] [1] = 1'b1;
  assign \A[19][206] [4] = 1'b1;
  assign \A[19][206] [3] = 1'b1;
  assign \A[19][206] [2] = 1'b1;
  assign \A[19][206] [1] = 1'b1;
  assign \A[19][206] [0] = 1'b1;
  assign \A[19][207] [1] = 1'b1;
  assign \A[19][208] [4] = 1'b1;
  assign \A[19][208] [3] = 1'b1;
  assign \A[19][208] [2] = 1'b1;
  assign \A[19][208] [1] = 1'b1;
  assign \A[19][208] [0] = 1'b1;
  assign \A[19][210] [4] = 1'b1;
  assign \A[19][210] [3] = 1'b1;
  assign \A[19][210] [2] = 1'b1;
  assign \A[19][210] [1] = 1'b1;
  assign \A[19][211] [1] = 1'b1;
  assign \A[19][212] [0] = 1'b1;
  assign \A[19][213] [0] = 1'b1;
  assign \A[19][214] [4] = 1'b1;
  assign \A[19][214] [3] = 1'b1;
  assign \A[19][214] [2] = 1'b1;
  assign \A[19][214] [1] = 1'b1;
  assign \A[19][215] [1] = 1'b1;
  assign \A[19][215] [0] = 1'b1;
  assign \A[19][217] [0] = 1'b1;
  assign \A[19][218] [4] = 1'b1;
  assign \A[19][218] [3] = 1'b1;
  assign \A[19][218] [2] = 1'b1;
  assign \A[19][218] [1] = 1'b1;
  assign \A[19][218] [0] = 1'b1;
  assign \A[19][219] [4] = 1'b1;
  assign \A[19][219] [3] = 1'b1;
  assign \A[19][219] [2] = 1'b1;
  assign \A[19][219] [1] = 1'b1;
  assign \A[19][221] [4] = 1'b1;
  assign \A[19][221] [3] = 1'b1;
  assign \A[19][221] [2] = 1'b1;
  assign \A[19][221] [1] = 1'b1;
  assign \A[19][221] [0] = 1'b1;
  assign \A[19][222] [4] = 1'b1;
  assign \A[19][222] [3] = 1'b1;
  assign \A[19][222] [2] = 1'b1;
  assign \A[19][222] [1] = 1'b1;
  assign \A[19][222] [0] = 1'b1;
  assign \A[19][224] [4] = 1'b1;
  assign \A[19][224] [3] = 1'b1;
  assign \A[19][224] [2] = 1'b1;
  assign \A[19][224] [1] = 1'b1;
  assign \A[19][227] [1] = 1'b1;
  assign \A[19][227] [0] = 1'b1;
  assign \A[19][229] [4] = 1'b1;
  assign \A[19][229] [3] = 1'b1;
  assign \A[19][229] [2] = 1'b1;
  assign \A[19][229] [1] = 1'b1;
  assign \A[19][231] [1] = 1'b1;
  assign \A[19][232] [4] = 1'b1;
  assign \A[19][232] [3] = 1'b1;
  assign \A[19][232] [2] = 1'b1;
  assign \A[19][232] [0] = 1'b1;
  assign \A[19][233] [0] = 1'b1;
  assign \A[19][234] [1] = 1'b1;
  assign \A[19][235] [4] = 1'b1;
  assign \A[19][235] [3] = 1'b1;
  assign \A[19][235] [2] = 1'b1;
  assign \A[19][235] [1] = 1'b1;
  assign \A[19][235] [0] = 1'b1;
  assign \A[19][236] [0] = 1'b1;
  assign \A[19][237] [0] = 1'b1;
  assign \A[19][238] [4] = 1'b1;
  assign \A[19][238] [3] = 1'b1;
  assign \A[19][238] [2] = 1'b1;
  assign \A[19][238] [0] = 1'b1;
  assign \A[19][242] [1] = 1'b1;
  assign \A[19][244] [4] = 1'b1;
  assign \A[19][244] [3] = 1'b1;
  assign \A[19][244] [2] = 1'b1;
  assign \A[19][244] [1] = 1'b1;
  assign \A[19][246] [0] = 1'b1;
  assign \A[19][248] [4] = 1'b1;
  assign \A[19][248] [3] = 1'b1;
  assign \A[19][248] [2] = 1'b1;
  assign \A[19][248] [0] = 1'b1;
  assign \A[19][250] [0] = 1'b1;
  assign \A[19][252] [0] = 1'b1;
  assign \A[19][253] [4] = 1'b1;
  assign \A[19][253] [3] = 1'b1;
  assign \A[19][253] [2] = 1'b1;
  assign \A[19][253] [1] = 1'b1;
  assign \A[19][254] [4] = 1'b1;
  assign \A[19][254] [3] = 1'b1;
  assign \A[19][254] [2] = 1'b1;
  assign \A[19][254] [1] = 1'b1;
  assign \A[19][254] [0] = 1'b1;
  VDW_WMUX5 U$1(.Z({ \dot_product_and_ReLU[19].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$2(.Z({ \dot_product_and_ReLU[19].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$3(.Z({ \dot_product_and_ReLU[19].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$4(.Z({ \dot_product_and_ReLU[19].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$5(.Z({ \dot_product_and_ReLU[19].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$6(.Z({ \dot_product_and_ReLU[19].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$7(.Z({ \dot_product_and_ReLU[19].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$8(.Z({ \dot_product_and_ReLU[19].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$9(.Z({ \dot_product_and_ReLU[19].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$10(.Z({ \dot_product_and_ReLU[19].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$11(.Z({ \dot_product_and_ReLU[19].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$12(.Z({ \dot_product_and_ReLU[19].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$13(.Z({ \dot_product_and_ReLU[19].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$14(.Z({ \dot_product_and_ReLU[19].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$15(.Z({ \dot_product_and_ReLU[19].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$16(.Z({ \dot_product_and_ReLU[19].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$17(.Z({ \dot_product_and_ReLU[19].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$18(.Z({ \dot_product_and_ReLU[19].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$19(.Z({ \dot_product_and_ReLU[19].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$20(.Z({ \dot_product_and_ReLU[19].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$21(.Z({ \dot_product_and_ReLU[19].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$22(.Z({ \dot_product_and_ReLU[19].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$23(.Z({ \dot_product_and_ReLU[19].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$24(.Z({ \dot_product_and_ReLU[19].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$25(.Z({ \dot_product_and_ReLU[19].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$26(.Z({ \dot_product_and_ReLU[19].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$27(.Z({ \dot_product_and_ReLU[19].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$28(.Z({ \dot_product_and_ReLU[19].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$29(.Z({ \dot_product_and_ReLU[19].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$30(.Z({ \dot_product_and_ReLU[19].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$31(.Z({ \dot_product_and_ReLU[19].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$32(.Z({ \dot_product_and_ReLU[19].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$33(.Z({ \dot_product_and_ReLU[19].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$34(.Z({ \dot_product_and_ReLU[19].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$35(.Z({ \dot_product_and_ReLU[19].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$36(.Z({ \dot_product_and_ReLU[19].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$37(.Z({ \dot_product_and_ReLU[19].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$38(.Z({ \dot_product_and_ReLU[19].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$39(.Z({ \dot_product_and_ReLU[19].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$40(.Z({ \dot_product_and_ReLU[19].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$41(.Z({ \dot_product_and_ReLU[19].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$42(.Z({ \dot_product_and_ReLU[19].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$43(.Z({ \dot_product_and_ReLU[19].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$44(.Z({ \dot_product_and_ReLU[19].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$45(.Z({ \dot_product_and_ReLU[19].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$46(.Z({ \dot_product_and_ReLU[19].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$47(.Z({ \dot_product_and_ReLU[19].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$48(.Z({ \dot_product_and_ReLU[19].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$49(.Z({ \dot_product_and_ReLU[19].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$50(.Z({ \dot_product_and_ReLU[19].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$51(.Z({ \dot_product_and_ReLU[19].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$52(.Z({ \dot_product_and_ReLU[19].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$53(.Z({ \dot_product_and_ReLU[19].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$54(.Z({ \dot_product_and_ReLU[19].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$55(.Z({ \dot_product_and_ReLU[19].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$56(.Z({ \dot_product_and_ReLU[19].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$57(.Z({ \dot_product_and_ReLU[19].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$58(.Z({ \dot_product_and_ReLU[19].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$59(.Z({ \dot_product_and_ReLU[19].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$60(.Z({ \dot_product_and_ReLU[19].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$61(.Z({ \dot_product_and_ReLU[19].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$62(.Z({ \dot_product_and_ReLU[19].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$63(.Z({ \dot_product_and_ReLU[19].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$64(.Z({ \dot_product_and_ReLU[19].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$65(.Z({ \dot_product_and_ReLU[19].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$66(.Z({ \dot_product_and_ReLU[19].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$67(.Z({ \dot_product_and_ReLU[19].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$68(.Z({ \dot_product_and_ReLU[19].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$69(.Z({ \dot_product_and_ReLU[19].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$70(.Z({ \dot_product_and_ReLU[19].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$71(.Z({ \dot_product_and_ReLU[19].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$72(.Z({ \dot_product_and_ReLU[19].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$73(.Z({ \dot_product_and_ReLU[19].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$74(.Z({ \dot_product_and_ReLU[19].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$75(.Z({ \dot_product_and_ReLU[19].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$76(.Z({ \dot_product_and_ReLU[19].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$77(.Z({ \dot_product_and_ReLU[19].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$78(.Z({ \dot_product_and_ReLU[19].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$79(.Z({ \dot_product_and_ReLU[19].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$80(.Z({ \dot_product_and_ReLU[19].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$81(.Z({ \dot_product_and_ReLU[19].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$82(.Z({ \dot_product_and_ReLU[19].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$83(.Z({ \dot_product_and_ReLU[19].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$84(.Z({ \dot_product_and_ReLU[19].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$85(.Z({ \dot_product_and_ReLU[19].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$86(.Z({ \dot_product_and_ReLU[19].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$87(.Z({ \dot_product_and_ReLU[19].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$88(.Z({ \dot_product_and_ReLU[19].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$89(.Z({ \dot_product_and_ReLU[19].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$90(.Z({ \dot_product_and_ReLU[19].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$91(.Z({ \dot_product_and_ReLU[19].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$92(.Z({ \dot_product_and_ReLU[19].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$93(.Z({ \dot_product_and_ReLU[19].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$94(.Z({ \dot_product_and_ReLU[19].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$95(.Z({ \dot_product_and_ReLU[19].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$96(.Z({ \dot_product_and_ReLU[19].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$97(.Z({ \dot_product_and_ReLU[19].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$98(.Z({ \dot_product_and_ReLU[19].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$99(.Z({ \dot_product_and_ReLU[19].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$100(.Z({ \dot_product_and_ReLU[19].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$101(.Z({ \dot_product_and_ReLU[19].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$102(.Z({ \dot_product_and_ReLU[19].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$103(.Z({ \dot_product_and_ReLU[19].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$104(.Z({ \dot_product_and_ReLU[19].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$105(.Z({ \dot_product_and_ReLU[19].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$106(.Z({ \dot_product_and_ReLU[19].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$107(.Z({ \dot_product_and_ReLU[19].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$108(.Z({ \dot_product_and_ReLU[19].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$109(.Z({ \dot_product_and_ReLU[19].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$110(.Z({ \dot_product_and_ReLU[19].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$111(.Z({ \dot_product_and_ReLU[19].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$112(.Z({ \dot_product_and_ReLU[19].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$113(.Z({ \dot_product_and_ReLU[19].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$114(.Z({ \dot_product_and_ReLU[19].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$115(.Z({ \dot_product_and_ReLU[19].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$116(.Z({ \dot_product_and_ReLU[19].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$117(.Z({ \dot_product_and_ReLU[19].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$118(.Z({ \dot_product_and_ReLU[19].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$119(.Z({ \dot_product_and_ReLU[19].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$120(.Z({ \dot_product_and_ReLU[19].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$121(.Z({ \dot_product_and_ReLU[19].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$122(.Z({ \dot_product_and_ReLU[19].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$123(.Z({ \dot_product_and_ReLU[19].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$124(.Z({ \dot_product_and_ReLU[19].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$125(.Z({ \dot_product_and_ReLU[19].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$126(.Z({ \dot_product_and_ReLU[19].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$127(.Z({ \dot_product_and_ReLU[19].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$128(.Z({ \dot_product_and_ReLU[19].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$129(.Z({ \dot_product_and_ReLU[19].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$130(.Z({ \dot_product_and_ReLU[19].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$131(.Z({ \dot_product_and_ReLU[19].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$132(.Z({ \dot_product_and_ReLU[19].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$133(.Z({ \dot_product_and_ReLU[19].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$134(.Z({ \dot_product_and_ReLU[19].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$135(.Z({ \dot_product_and_ReLU[19].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$136(.Z({ \dot_product_and_ReLU[19].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$137(.Z({ \dot_product_and_ReLU[19].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$138(.Z({ \dot_product_and_ReLU[19].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$139(.Z({ \dot_product_and_ReLU[19].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$140(.Z({ \dot_product_and_ReLU[19].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$141(.Z({ \dot_product_and_ReLU[19].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$142(.Z({ \dot_product_and_ReLU[19].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$143(.Z({ \dot_product_and_ReLU[19].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$144(.Z({ \dot_product_and_ReLU[19].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$145(.Z({ \dot_product_and_ReLU[19].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$146(.Z({ \dot_product_and_ReLU[19].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$147(.Z({ \dot_product_and_ReLU[19].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$148(.Z({ \dot_product_and_ReLU[19].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$149(.Z({ \dot_product_and_ReLU[19].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$150(.Z({ \dot_product_and_ReLU[19].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$151(.Z({ \dot_product_and_ReLU[19].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$152(.Z({ \dot_product_and_ReLU[19].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$153(.Z({ \dot_product_and_ReLU[19].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$154(.Z({ \dot_product_and_ReLU[19].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$155(.Z({ \dot_product_and_ReLU[19].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$156(.Z({ \dot_product_and_ReLU[19].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$157(.Z({ \dot_product_and_ReLU[19].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$158(.Z({ \dot_product_and_ReLU[19].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$159(.Z({ \dot_product_and_ReLU[19].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$160(.Z({ \dot_product_and_ReLU[19].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$161(.Z({ \dot_product_and_ReLU[19].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$162(.Z({ \dot_product_and_ReLU[19].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$163(.Z({ \dot_product_and_ReLU[19].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$164(.Z({ \dot_product_and_ReLU[19].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$165(.Z({ \dot_product_and_ReLU[19].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$166(.Z({ \dot_product_and_ReLU[19].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$167(.Z({ \dot_product_and_ReLU[19].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$168(.Z({ \dot_product_and_ReLU[19].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$169(.Z({ \dot_product_and_ReLU[19].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$170(.Z({ \dot_product_and_ReLU[19].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$171(.Z({ \dot_product_and_ReLU[19].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$172(.Z({ \dot_product_and_ReLU[19].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$173(.Z({ \dot_product_and_ReLU[19].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$174(.Z({ \dot_product_and_ReLU[19].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$175(.Z({ \dot_product_and_ReLU[19].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$176(.Z({ \dot_product_and_ReLU[19].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$177(.Z({ \dot_product_and_ReLU[19].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$178(.Z({ \dot_product_and_ReLU[19].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$179(.Z({ \dot_product_and_ReLU[19].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$180(.Z({ \dot_product_and_ReLU[19].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$181(.Z({ \dot_product_and_ReLU[19].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$182(.Z({ \dot_product_and_ReLU[19].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$183(.Z({ \dot_product_and_ReLU[19].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$184(.Z({ \dot_product_and_ReLU[19].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$185(.Z({ \dot_product_and_ReLU[19].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$186(.Z({ \dot_product_and_ReLU[19].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$187(.Z({ \dot_product_and_ReLU[19].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$188(.Z({ \dot_product_and_ReLU[19].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$189(.Z({ \dot_product_and_ReLU[19].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$190(.Z({ \dot_product_and_ReLU[19].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$191(.Z({ \dot_product_and_ReLU[19].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$192(.Z({ \dot_product_and_ReLU[19].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$193(.Z({ \dot_product_and_ReLU[19].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$194(.Z({ \dot_product_and_ReLU[19].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$195(.Z({ \dot_product_and_ReLU[19].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$196(.Z({ \dot_product_and_ReLU[19].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$197(.Z({ \dot_product_and_ReLU[19].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$198(.Z({ \dot_product_and_ReLU[19].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$199(.Z({ \dot_product_and_ReLU[19].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$200(.Z({ \dot_product_and_ReLU[19].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$201(.Z({ \dot_product_and_ReLU[19].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$202(.Z({ \dot_product_and_ReLU[19].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$203(.Z({ \dot_product_and_ReLU[19].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$204(.Z({ \dot_product_and_ReLU[19].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$205(.Z({ \dot_product_and_ReLU[19].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$206(.Z({ \dot_product_and_ReLU[19].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$207(.Z({ \dot_product_and_ReLU[19].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$208(.Z({ \dot_product_and_ReLU[19].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$209(.Z({ \dot_product_and_ReLU[19].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$210(.Z({ \dot_product_and_ReLU[19].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$211(.Z({ \dot_product_and_ReLU[19].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$212(.Z({ \dot_product_and_ReLU[19].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$213(.Z({ \dot_product_and_ReLU[19].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$214(.Z({ \dot_product_and_ReLU[19].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$215(.Z({ \dot_product_and_ReLU[19].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$216(.Z({ \dot_product_and_ReLU[19].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$217(.Z({ \dot_product_and_ReLU[19].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$218(.Z({ \dot_product_and_ReLU[19].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$219(.Z({ \dot_product_and_ReLU[19].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$220(.Z({ \dot_product_and_ReLU[19].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$221(.Z({ \dot_product_and_ReLU[19].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$222(.Z({ \dot_product_and_ReLU[19].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$223(.Z({ \dot_product_and_ReLU[19].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$224(.Z({ \dot_product_and_ReLU[19].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$225(.Z({ \dot_product_and_ReLU[19].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$226(.Z({ \dot_product_and_ReLU[19].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$227(.Z({ \dot_product_and_ReLU[19].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$228(.Z({ \dot_product_and_ReLU[19].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$229(.Z({ \dot_product_and_ReLU[19].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$230(.Z({ \dot_product_and_ReLU[19].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$231(.Z({ \dot_product_and_ReLU[19].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$232(.Z({ \dot_product_and_ReLU[19].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$233(.Z({ \dot_product_and_ReLU[19].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$234(.Z({ \dot_product_and_ReLU[19].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$235(.Z({ \dot_product_and_ReLU[19].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$236(.Z({ \dot_product_and_ReLU[19].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$237(.Z({ \dot_product_and_ReLU[19].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$238(.Z({ \dot_product_and_ReLU[19].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$239(.Z({ \dot_product_and_ReLU[19].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$240(.Z({ \dot_product_and_ReLU[19].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$241(.Z({ \dot_product_and_ReLU[19].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$242(.Z({ \dot_product_and_ReLU[19].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$243(.Z({ \dot_product_and_ReLU[19].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$244(.Z({ \dot_product_and_ReLU[19].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$245(.Z({ \dot_product_and_ReLU[19].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$246(.Z({ \dot_product_and_ReLU[19].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$247(.Z({ \dot_product_and_ReLU[19].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$248(.Z({ \dot_product_and_ReLU[19].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$249(.Z({ \dot_product_and_ReLU[19].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$250(.Z({ \dot_product_and_ReLU[19].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$251(.Z({ \dot_product_and_ReLU[19].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$252(.Z({ \dot_product_and_ReLU[19].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$253(.Z({ \dot_product_and_ReLU[19].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$254(.Z({ \dot_product_and_ReLU[19].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$255(.Z({ \dot_product_and_ReLU[19].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$256(.Z({ \dot_product_and_ReLU[19].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[19][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$257(.Z({ \dot_product_and_ReLU[18].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$258(.Z({ \dot_product_and_ReLU[18].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$259(.Z({ \dot_product_and_ReLU[18].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$260(.Z({ \dot_product_and_ReLU[18].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$261(.Z({ \dot_product_and_ReLU[18].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$262(.Z({ \dot_product_and_ReLU[18].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$263(.Z({ \dot_product_and_ReLU[18].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$264(.Z({ \dot_product_and_ReLU[18].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$265(.Z({ \dot_product_and_ReLU[18].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$266(.Z({ \dot_product_and_ReLU[18].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$267(.Z({ \dot_product_and_ReLU[18].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$268(.Z({ \dot_product_and_ReLU[18].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$269(.Z({ \dot_product_and_ReLU[18].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$270(.Z({ \dot_product_and_ReLU[18].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$271(.Z({ \dot_product_and_ReLU[18].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$272(.Z({ \dot_product_and_ReLU[18].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$273(.Z({ \dot_product_and_ReLU[18].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$274(.Z({ \dot_product_and_ReLU[18].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$275(.Z({ \dot_product_and_ReLU[18].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$276(.Z({ \dot_product_and_ReLU[18].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$277(.Z({ \dot_product_and_ReLU[18].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$278(.Z({ \dot_product_and_ReLU[18].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$279(.Z({ \dot_product_and_ReLU[18].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$280(.Z({ \dot_product_and_ReLU[18].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$281(.Z({ \dot_product_and_ReLU[18].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$282(.Z({ \dot_product_and_ReLU[18].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$283(.Z({ \dot_product_and_ReLU[18].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$284(.Z({ \dot_product_and_ReLU[18].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$285(.Z({ \dot_product_and_ReLU[18].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$286(.Z({ \dot_product_and_ReLU[18].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$287(.Z({ \dot_product_and_ReLU[18].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$288(.Z({ \dot_product_and_ReLU[18].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$289(.Z({ \dot_product_and_ReLU[18].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$290(.Z({ \dot_product_and_ReLU[18].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$291(.Z({ \dot_product_and_ReLU[18].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$292(.Z({ \dot_product_and_ReLU[18].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$293(.Z({ \dot_product_and_ReLU[18].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$294(.Z({ \dot_product_and_ReLU[18].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$295(.Z({ \dot_product_and_ReLU[18].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$296(.Z({ \dot_product_and_ReLU[18].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$297(.Z({ \dot_product_and_ReLU[18].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$298(.Z({ \dot_product_and_ReLU[18].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$299(.Z({ \dot_product_and_ReLU[18].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$300(.Z({ \dot_product_and_ReLU[18].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$301(.Z({ \dot_product_and_ReLU[18].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$302(.Z({ \dot_product_and_ReLU[18].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$303(.Z({ \dot_product_and_ReLU[18].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$304(.Z({ \dot_product_and_ReLU[18].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$305(.Z({ \dot_product_and_ReLU[18].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$306(.Z({ \dot_product_and_ReLU[18].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$307(.Z({ \dot_product_and_ReLU[18].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$308(.Z({ \dot_product_and_ReLU[18].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$309(.Z({ \dot_product_and_ReLU[18].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$310(.Z({ \dot_product_and_ReLU[18].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$311(.Z({ \dot_product_and_ReLU[18].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$312(.Z({ \dot_product_and_ReLU[18].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$313(.Z({ \dot_product_and_ReLU[18].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$314(.Z({ \dot_product_and_ReLU[18].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$315(.Z({ \dot_product_and_ReLU[18].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$316(.Z({ \dot_product_and_ReLU[18].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$317(.Z({ \dot_product_and_ReLU[18].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$318(.Z({ \dot_product_and_ReLU[18].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$319(.Z({ \dot_product_and_ReLU[18].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$320(.Z({ \dot_product_and_ReLU[18].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$321(.Z({ \dot_product_and_ReLU[18].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$322(.Z({ \dot_product_and_ReLU[18].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$323(.Z({ \dot_product_and_ReLU[18].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$324(.Z({ \dot_product_and_ReLU[18].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$325(.Z({ \dot_product_and_ReLU[18].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$326(.Z({ \dot_product_and_ReLU[18].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$327(.Z({ \dot_product_and_ReLU[18].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$328(.Z({ \dot_product_and_ReLU[18].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$329(.Z({ \dot_product_and_ReLU[18].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$330(.Z({ \dot_product_and_ReLU[18].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$331(.Z({ \dot_product_and_ReLU[18].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$332(.Z({ \dot_product_and_ReLU[18].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$333(.Z({ \dot_product_and_ReLU[18].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$334(.Z({ \dot_product_and_ReLU[18].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$335(.Z({ \dot_product_and_ReLU[18].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$336(.Z({ \dot_product_and_ReLU[18].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$337(.Z({ \dot_product_and_ReLU[18].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$338(.Z({ \dot_product_and_ReLU[18].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$339(.Z({ \dot_product_and_ReLU[18].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$340(.Z({ \dot_product_and_ReLU[18].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$341(.Z({ \dot_product_and_ReLU[18].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$342(.Z({ \dot_product_and_ReLU[18].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$343(.Z({ \dot_product_and_ReLU[18].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$344(.Z({ \dot_product_and_ReLU[18].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$345(.Z({ \dot_product_and_ReLU[18].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$346(.Z({ \dot_product_and_ReLU[18].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$347(.Z({ \dot_product_and_ReLU[18].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$348(.Z({ \dot_product_and_ReLU[18].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$349(.Z({ \dot_product_and_ReLU[18].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$350(.Z({ \dot_product_and_ReLU[18].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$351(.Z({ \dot_product_and_ReLU[18].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$352(.Z({ \dot_product_and_ReLU[18].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$353(.Z({ \dot_product_and_ReLU[18].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$354(.Z({ \dot_product_and_ReLU[18].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$355(.Z({ \dot_product_and_ReLU[18].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$356(.Z({ \dot_product_and_ReLU[18].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$357(.Z({ \dot_product_and_ReLU[18].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$358(.Z({ \dot_product_and_ReLU[18].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$359(.Z({ \dot_product_and_ReLU[18].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$360(.Z({ \dot_product_and_ReLU[18].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$361(.Z({ \dot_product_and_ReLU[18].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$362(.Z({ \dot_product_and_ReLU[18].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$363(.Z({ \dot_product_and_ReLU[18].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$364(.Z({ \dot_product_and_ReLU[18].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$365(.Z({ \dot_product_and_ReLU[18].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$366(.Z({ \dot_product_and_ReLU[18].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$367(.Z({ \dot_product_and_ReLU[18].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$368(.Z({ \dot_product_and_ReLU[18].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$369(.Z({ \dot_product_and_ReLU[18].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$370(.Z({ \dot_product_and_ReLU[18].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$371(.Z({ \dot_product_and_ReLU[18].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$372(.Z({ \dot_product_and_ReLU[18].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$373(.Z({ \dot_product_and_ReLU[18].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$374(.Z({ \dot_product_and_ReLU[18].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$375(.Z({ \dot_product_and_ReLU[18].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$376(.Z({ \dot_product_and_ReLU[18].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$377(.Z({ \dot_product_and_ReLU[18].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$378(.Z({ \dot_product_and_ReLU[18].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$379(.Z({ \dot_product_and_ReLU[18].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$380(.Z({ \dot_product_and_ReLU[18].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$381(.Z({ \dot_product_and_ReLU[18].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$382(.Z({ \dot_product_and_ReLU[18].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$383(.Z({ \dot_product_and_ReLU[18].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$384(.Z({ \dot_product_and_ReLU[18].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$385(.Z({ \dot_product_and_ReLU[18].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$386(.Z({ \dot_product_and_ReLU[18].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$387(.Z({ \dot_product_and_ReLU[18].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$388(.Z({ \dot_product_and_ReLU[18].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$389(.Z({ \dot_product_and_ReLU[18].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$390(.Z({ \dot_product_and_ReLU[18].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$391(.Z({ \dot_product_and_ReLU[18].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$392(.Z({ \dot_product_and_ReLU[18].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$393(.Z({ \dot_product_and_ReLU[18].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$394(.Z({ \dot_product_and_ReLU[18].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$395(.Z({ \dot_product_and_ReLU[18].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$396(.Z({ \dot_product_and_ReLU[18].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$397(.Z({ \dot_product_and_ReLU[18].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$398(.Z({ \dot_product_and_ReLU[18].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$399(.Z({ \dot_product_and_ReLU[18].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$400(.Z({ \dot_product_and_ReLU[18].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$401(.Z({ \dot_product_and_ReLU[18].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$402(.Z({ \dot_product_and_ReLU[18].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$403(.Z({ \dot_product_and_ReLU[18].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$404(.Z({ \dot_product_and_ReLU[18].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$405(.Z({ \dot_product_and_ReLU[18].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$406(.Z({ \dot_product_and_ReLU[18].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$407(.Z({ \dot_product_and_ReLU[18].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$408(.Z({ \dot_product_and_ReLU[18].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$409(.Z({ \dot_product_and_ReLU[18].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$410(.Z({ \dot_product_and_ReLU[18].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$411(.Z({ \dot_product_and_ReLU[18].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$412(.Z({ \dot_product_and_ReLU[18].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$413(.Z({ \dot_product_and_ReLU[18].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$414(.Z({ \dot_product_and_ReLU[18].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$415(.Z({ \dot_product_and_ReLU[18].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$416(.Z({ \dot_product_and_ReLU[18].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$417(.Z({ \dot_product_and_ReLU[18].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$418(.Z({ \dot_product_and_ReLU[18].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$419(.Z({ \dot_product_and_ReLU[18].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$420(.Z({ \dot_product_and_ReLU[18].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$421(.Z({ \dot_product_and_ReLU[18].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$422(.Z({ \dot_product_and_ReLU[18].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$423(.Z({ \dot_product_and_ReLU[18].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$424(.Z({ \dot_product_and_ReLU[18].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$425(.Z({ \dot_product_and_ReLU[18].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$426(.Z({ \dot_product_and_ReLU[18].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$427(.Z({ \dot_product_and_ReLU[18].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$428(.Z({ \dot_product_and_ReLU[18].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$429(.Z({ \dot_product_and_ReLU[18].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$430(.Z({ \dot_product_and_ReLU[18].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$431(.Z({ \dot_product_and_ReLU[18].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$432(.Z({ \dot_product_and_ReLU[18].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$433(.Z({ \dot_product_and_ReLU[18].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$434(.Z({ \dot_product_and_ReLU[18].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$435(.Z({ \dot_product_and_ReLU[18].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$436(.Z({ \dot_product_and_ReLU[18].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$437(.Z({ \dot_product_and_ReLU[18].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$438(.Z({ \dot_product_and_ReLU[18].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$439(.Z({ \dot_product_and_ReLU[18].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$440(.Z({ \dot_product_and_ReLU[18].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$441(.Z({ \dot_product_and_ReLU[18].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$442(.Z({ \dot_product_and_ReLU[18].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$443(.Z({ \dot_product_and_ReLU[18].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$444(.Z({ \dot_product_and_ReLU[18].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$445(.Z({ \dot_product_and_ReLU[18].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$446(.Z({ \dot_product_and_ReLU[18].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$447(.Z({ \dot_product_and_ReLU[18].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$448(.Z({ \dot_product_and_ReLU[18].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$449(.Z({ \dot_product_and_ReLU[18].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$450(.Z({ \dot_product_and_ReLU[18].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$451(.Z({ \dot_product_and_ReLU[18].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$452(.Z({ \dot_product_and_ReLU[18].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$453(.Z({ \dot_product_and_ReLU[18].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$454(.Z({ \dot_product_and_ReLU[18].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$455(.Z({ \dot_product_and_ReLU[18].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$456(.Z({ \dot_product_and_ReLU[18].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$457(.Z({ \dot_product_and_ReLU[18].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$458(.Z({ \dot_product_and_ReLU[18].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$459(.Z({ \dot_product_and_ReLU[18].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$460(.Z({ \dot_product_and_ReLU[18].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$461(.Z({ \dot_product_and_ReLU[18].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$462(.Z({ \dot_product_and_ReLU[18].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$463(.Z({ \dot_product_and_ReLU[18].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$464(.Z({ \dot_product_and_ReLU[18].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$465(.Z({ \dot_product_and_ReLU[18].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$466(.Z({ \dot_product_and_ReLU[18].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$467(.Z({ \dot_product_and_ReLU[18].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$468(.Z({ \dot_product_and_ReLU[18].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$469(.Z({ \dot_product_and_ReLU[18].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$470(.Z({ \dot_product_and_ReLU[18].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$471(.Z({ \dot_product_and_ReLU[18].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$472(.Z({ \dot_product_and_ReLU[18].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$473(.Z({ \dot_product_and_ReLU[18].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$474(.Z({ \dot_product_and_ReLU[18].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$475(.Z({ \dot_product_and_ReLU[18].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$476(.Z({ \dot_product_and_ReLU[18].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$477(.Z({ \dot_product_and_ReLU[18].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$478(.Z({ \dot_product_and_ReLU[18].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$479(.Z({ \dot_product_and_ReLU[18].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$480(.Z({ \dot_product_and_ReLU[18].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$481(.Z({ \dot_product_and_ReLU[18].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$482(.Z({ \dot_product_and_ReLU[18].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$483(.Z({ \dot_product_and_ReLU[18].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$484(.Z({ \dot_product_and_ReLU[18].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$485(.Z({ \dot_product_and_ReLU[18].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$486(.Z({ \dot_product_and_ReLU[18].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$487(.Z({ \dot_product_and_ReLU[18].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$488(.Z({ \dot_product_and_ReLU[18].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$489(.Z({ \dot_product_and_ReLU[18].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$490(.Z({ \dot_product_and_ReLU[18].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$491(.Z({ \dot_product_and_ReLU[18].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$492(.Z({ \dot_product_and_ReLU[18].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$493(.Z({ \dot_product_and_ReLU[18].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$494(.Z({ \dot_product_and_ReLU[18].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$495(.Z({ \dot_product_and_ReLU[18].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$496(.Z({ \dot_product_and_ReLU[18].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$497(.Z({ \dot_product_and_ReLU[18].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$498(.Z({ \dot_product_and_ReLU[18].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$499(.Z({ \dot_product_and_ReLU[18].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$500(.Z({ \dot_product_and_ReLU[18].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$501(.Z({ \dot_product_and_ReLU[18].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$502(.Z({ \dot_product_and_ReLU[18].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$503(.Z({ \dot_product_and_ReLU[18].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$504(.Z({ \dot_product_and_ReLU[18].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$505(.Z({ \dot_product_and_ReLU[18].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$506(.Z({ \dot_product_and_ReLU[18].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$507(.Z({ \dot_product_and_ReLU[18].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$508(.Z({ \dot_product_and_ReLU[18].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$509(.Z({ \dot_product_and_ReLU[18].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$510(.Z({ \dot_product_and_ReLU[18].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$511(.Z({ \dot_product_and_ReLU[18].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$512(.Z({ \dot_product_and_ReLU[18].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[18][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$513(.Z({ \dot_product_and_ReLU[17].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$514(.Z({ \dot_product_and_ReLU[17].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$515(.Z({ \dot_product_and_ReLU[17].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$516(.Z({ \dot_product_and_ReLU[17].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$517(.Z({ \dot_product_and_ReLU[17].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$518(.Z({ \dot_product_and_ReLU[17].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$519(.Z({ \dot_product_and_ReLU[17].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$520(.Z({ \dot_product_and_ReLU[17].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$521(.Z({ \dot_product_and_ReLU[17].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$522(.Z({ \dot_product_and_ReLU[17].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$523(.Z({ \dot_product_and_ReLU[17].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$524(.Z({ \dot_product_and_ReLU[17].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$525(.Z({ \dot_product_and_ReLU[17].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$526(.Z({ \dot_product_and_ReLU[17].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$527(.Z({ \dot_product_and_ReLU[17].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$528(.Z({ \dot_product_and_ReLU[17].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$529(.Z({ \dot_product_and_ReLU[17].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$530(.Z({ \dot_product_and_ReLU[17].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$531(.Z({ \dot_product_and_ReLU[17].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$532(.Z({ \dot_product_and_ReLU[17].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$533(.Z({ \dot_product_and_ReLU[17].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$534(.Z({ \dot_product_and_ReLU[17].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$535(.Z({ \dot_product_and_ReLU[17].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$536(.Z({ \dot_product_and_ReLU[17].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$537(.Z({ \dot_product_and_ReLU[17].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$538(.Z({ \dot_product_and_ReLU[17].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$539(.Z({ \dot_product_and_ReLU[17].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$540(.Z({ \dot_product_and_ReLU[17].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$541(.Z({ \dot_product_and_ReLU[17].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$542(.Z({ \dot_product_and_ReLU[17].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$543(.Z({ \dot_product_and_ReLU[17].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$544(.Z({ \dot_product_and_ReLU[17].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$545(.Z({ \dot_product_and_ReLU[17].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$546(.Z({ \dot_product_and_ReLU[17].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$547(.Z({ \dot_product_and_ReLU[17].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$548(.Z({ \dot_product_and_ReLU[17].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$549(.Z({ \dot_product_and_ReLU[17].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$550(.Z({ \dot_product_and_ReLU[17].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$551(.Z({ \dot_product_and_ReLU[17].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$552(.Z({ \dot_product_and_ReLU[17].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$553(.Z({ \dot_product_and_ReLU[17].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$554(.Z({ \dot_product_and_ReLU[17].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$555(.Z({ \dot_product_and_ReLU[17].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$556(.Z({ \dot_product_and_ReLU[17].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$557(.Z({ \dot_product_and_ReLU[17].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$558(.Z({ \dot_product_and_ReLU[17].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$559(.Z({ \dot_product_and_ReLU[17].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$560(.Z({ \dot_product_and_ReLU[17].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$561(.Z({ \dot_product_and_ReLU[17].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$562(.Z({ \dot_product_and_ReLU[17].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$563(.Z({ \dot_product_and_ReLU[17].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$564(.Z({ \dot_product_and_ReLU[17].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$565(.Z({ \dot_product_and_ReLU[17].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$566(.Z({ \dot_product_and_ReLU[17].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$567(.Z({ \dot_product_and_ReLU[17].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$568(.Z({ \dot_product_and_ReLU[17].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$569(.Z({ \dot_product_and_ReLU[17].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$570(.Z({ \dot_product_and_ReLU[17].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$571(.Z({ \dot_product_and_ReLU[17].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$572(.Z({ \dot_product_and_ReLU[17].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$573(.Z({ \dot_product_and_ReLU[17].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$574(.Z({ \dot_product_and_ReLU[17].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$575(.Z({ \dot_product_and_ReLU[17].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$576(.Z({ \dot_product_and_ReLU[17].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$577(.Z({ \dot_product_and_ReLU[17].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$578(.Z({ \dot_product_and_ReLU[17].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$579(.Z({ \dot_product_and_ReLU[17].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$580(.Z({ \dot_product_and_ReLU[17].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$581(.Z({ \dot_product_and_ReLU[17].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$582(.Z({ \dot_product_and_ReLU[17].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$583(.Z({ \dot_product_and_ReLU[17].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$584(.Z({ \dot_product_and_ReLU[17].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$585(.Z({ \dot_product_and_ReLU[17].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$586(.Z({ \dot_product_and_ReLU[17].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$587(.Z({ \dot_product_and_ReLU[17].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$588(.Z({ \dot_product_and_ReLU[17].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$589(.Z({ \dot_product_and_ReLU[17].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$590(.Z({ \dot_product_and_ReLU[17].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$591(.Z({ \dot_product_and_ReLU[17].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$592(.Z({ \dot_product_and_ReLU[17].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$593(.Z({ \dot_product_and_ReLU[17].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$594(.Z({ \dot_product_and_ReLU[17].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$595(.Z({ \dot_product_and_ReLU[17].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$596(.Z({ \dot_product_and_ReLU[17].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$597(.Z({ \dot_product_and_ReLU[17].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$598(.Z({ \dot_product_and_ReLU[17].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$599(.Z({ \dot_product_and_ReLU[17].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$600(.Z({ \dot_product_and_ReLU[17].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$601(.Z({ \dot_product_and_ReLU[17].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$602(.Z({ \dot_product_and_ReLU[17].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$603(.Z({ \dot_product_and_ReLU[17].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$604(.Z({ \dot_product_and_ReLU[17].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$605(.Z({ \dot_product_and_ReLU[17].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$606(.Z({ \dot_product_and_ReLU[17].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$607(.Z({ \dot_product_and_ReLU[17].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$608(.Z({ \dot_product_and_ReLU[17].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$609(.Z({ \dot_product_and_ReLU[17].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$610(.Z({ \dot_product_and_ReLU[17].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$611(.Z({ \dot_product_and_ReLU[17].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$612(.Z({ \dot_product_and_ReLU[17].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$613(.Z({ \dot_product_and_ReLU[17].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$614(.Z({ \dot_product_and_ReLU[17].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$615(.Z({ \dot_product_and_ReLU[17].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$616(.Z({ \dot_product_and_ReLU[17].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$617(.Z({ \dot_product_and_ReLU[17].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$618(.Z({ \dot_product_and_ReLU[17].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$619(.Z({ \dot_product_and_ReLU[17].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$620(.Z({ \dot_product_and_ReLU[17].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$621(.Z({ \dot_product_and_ReLU[17].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$622(.Z({ \dot_product_and_ReLU[17].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$623(.Z({ \dot_product_and_ReLU[17].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$624(.Z({ \dot_product_and_ReLU[17].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$625(.Z({ \dot_product_and_ReLU[17].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$626(.Z({ \dot_product_and_ReLU[17].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$627(.Z({ \dot_product_and_ReLU[17].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$628(.Z({ \dot_product_and_ReLU[17].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$629(.Z({ \dot_product_and_ReLU[17].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$630(.Z({ \dot_product_and_ReLU[17].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$631(.Z({ \dot_product_and_ReLU[17].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$632(.Z({ \dot_product_and_ReLU[17].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$633(.Z({ \dot_product_and_ReLU[17].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$634(.Z({ \dot_product_and_ReLU[17].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$635(.Z({ \dot_product_and_ReLU[17].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$636(.Z({ \dot_product_and_ReLU[17].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$637(.Z({ \dot_product_and_ReLU[17].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$638(.Z({ \dot_product_and_ReLU[17].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$639(.Z({ \dot_product_and_ReLU[17].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$640(.Z({ \dot_product_and_ReLU[17].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$641(.Z({ \dot_product_and_ReLU[17].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$642(.Z({ \dot_product_and_ReLU[17].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$643(.Z({ \dot_product_and_ReLU[17].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$644(.Z({ \dot_product_and_ReLU[17].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$645(.Z({ \dot_product_and_ReLU[17].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$646(.Z({ \dot_product_and_ReLU[17].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$647(.Z({ \dot_product_and_ReLU[17].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$648(.Z({ \dot_product_and_ReLU[17].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$649(.Z({ \dot_product_and_ReLU[17].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$650(.Z({ \dot_product_and_ReLU[17].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$651(.Z({ \dot_product_and_ReLU[17].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$652(.Z({ \dot_product_and_ReLU[17].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$653(.Z({ \dot_product_and_ReLU[17].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$654(.Z({ \dot_product_and_ReLU[17].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$655(.Z({ \dot_product_and_ReLU[17].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$656(.Z({ \dot_product_and_ReLU[17].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$657(.Z({ \dot_product_and_ReLU[17].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$658(.Z({ \dot_product_and_ReLU[17].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$659(.Z({ \dot_product_and_ReLU[17].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$660(.Z({ \dot_product_and_ReLU[17].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$661(.Z({ \dot_product_and_ReLU[17].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$662(.Z({ \dot_product_and_ReLU[17].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$663(.Z({ \dot_product_and_ReLU[17].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$664(.Z({ \dot_product_and_ReLU[17].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$665(.Z({ \dot_product_and_ReLU[17].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$666(.Z({ \dot_product_and_ReLU[17].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$667(.Z({ \dot_product_and_ReLU[17].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$668(.Z({ \dot_product_and_ReLU[17].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$669(.Z({ \dot_product_and_ReLU[17].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$670(.Z({ \dot_product_and_ReLU[17].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$671(.Z({ \dot_product_and_ReLU[17].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$672(.Z({ \dot_product_and_ReLU[17].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$673(.Z({ \dot_product_and_ReLU[17].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$674(.Z({ \dot_product_and_ReLU[17].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$675(.Z({ \dot_product_and_ReLU[17].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$676(.Z({ \dot_product_and_ReLU[17].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$677(.Z({ \dot_product_and_ReLU[17].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$678(.Z({ \dot_product_and_ReLU[17].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$679(.Z({ \dot_product_and_ReLU[17].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$680(.Z({ \dot_product_and_ReLU[17].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$681(.Z({ \dot_product_and_ReLU[17].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$682(.Z({ \dot_product_and_ReLU[17].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$683(.Z({ \dot_product_and_ReLU[17].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$684(.Z({ \dot_product_and_ReLU[17].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$685(.Z({ \dot_product_and_ReLU[17].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$686(.Z({ \dot_product_and_ReLU[17].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$687(.Z({ \dot_product_and_ReLU[17].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$688(.Z({ \dot_product_and_ReLU[17].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$689(.Z({ \dot_product_and_ReLU[17].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$690(.Z({ \dot_product_and_ReLU[17].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$691(.Z({ \dot_product_and_ReLU[17].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$692(.Z({ \dot_product_and_ReLU[17].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$693(.Z({ \dot_product_and_ReLU[17].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$694(.Z({ \dot_product_and_ReLU[17].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$695(.Z({ \dot_product_and_ReLU[17].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$696(.Z({ \dot_product_and_ReLU[17].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$697(.Z({ \dot_product_and_ReLU[17].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$698(.Z({ \dot_product_and_ReLU[17].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$699(.Z({ \dot_product_and_ReLU[17].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$700(.Z({ \dot_product_and_ReLU[17].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$701(.Z({ \dot_product_and_ReLU[17].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$702(.Z({ \dot_product_and_ReLU[17].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$703(.Z({ \dot_product_and_ReLU[17].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$704(.Z({ \dot_product_and_ReLU[17].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$705(.Z({ \dot_product_and_ReLU[17].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$706(.Z({ \dot_product_and_ReLU[17].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$707(.Z({ \dot_product_and_ReLU[17].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$708(.Z({ \dot_product_and_ReLU[17].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$709(.Z({ \dot_product_and_ReLU[17].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$710(.Z({ \dot_product_and_ReLU[17].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$711(.Z({ \dot_product_and_ReLU[17].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$712(.Z({ \dot_product_and_ReLU[17].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$713(.Z({ \dot_product_and_ReLU[17].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$714(.Z({ \dot_product_and_ReLU[17].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$715(.Z({ \dot_product_and_ReLU[17].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$716(.Z({ \dot_product_and_ReLU[17].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$717(.Z({ \dot_product_and_ReLU[17].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$718(.Z({ \dot_product_and_ReLU[17].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$719(.Z({ \dot_product_and_ReLU[17].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$720(.Z({ \dot_product_and_ReLU[17].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$721(.Z({ \dot_product_and_ReLU[17].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$722(.Z({ \dot_product_and_ReLU[17].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$723(.Z({ \dot_product_and_ReLU[17].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$724(.Z({ \dot_product_and_ReLU[17].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$725(.Z({ \dot_product_and_ReLU[17].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$726(.Z({ \dot_product_and_ReLU[17].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$727(.Z({ \dot_product_and_ReLU[17].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$728(.Z({ \dot_product_and_ReLU[17].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$729(.Z({ \dot_product_and_ReLU[17].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$730(.Z({ \dot_product_and_ReLU[17].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$731(.Z({ \dot_product_and_ReLU[17].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$732(.Z({ \dot_product_and_ReLU[17].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$733(.Z({ \dot_product_and_ReLU[17].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$734(.Z({ \dot_product_and_ReLU[17].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$735(.Z({ \dot_product_and_ReLU[17].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$736(.Z({ \dot_product_and_ReLU[17].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$737(.Z({ \dot_product_and_ReLU[17].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$738(.Z({ \dot_product_and_ReLU[17].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$739(.Z({ \dot_product_and_ReLU[17].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$740(.Z({ \dot_product_and_ReLU[17].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$741(.Z({ \dot_product_and_ReLU[17].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$742(.Z({ \dot_product_and_ReLU[17].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$743(.Z({ \dot_product_and_ReLU[17].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$744(.Z({ \dot_product_and_ReLU[17].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$745(.Z({ \dot_product_and_ReLU[17].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$746(.Z({ \dot_product_and_ReLU[17].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$747(.Z({ \dot_product_and_ReLU[17].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$748(.Z({ \dot_product_and_ReLU[17].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$749(.Z({ \dot_product_and_ReLU[17].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$750(.Z({ \dot_product_and_ReLU[17].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$751(.Z({ \dot_product_and_ReLU[17].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$752(.Z({ \dot_product_and_ReLU[17].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$753(.Z({ \dot_product_and_ReLU[17].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$754(.Z({ \dot_product_and_ReLU[17].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$755(.Z({ \dot_product_and_ReLU[17].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$756(.Z({ \dot_product_and_ReLU[17].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$757(.Z({ \dot_product_and_ReLU[17].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$758(.Z({ \dot_product_and_ReLU[17].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$759(.Z({ \dot_product_and_ReLU[17].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$760(.Z({ \dot_product_and_ReLU[17].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$761(.Z({ \dot_product_and_ReLU[17].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$762(.Z({ \dot_product_and_ReLU[17].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$763(.Z({ \dot_product_and_ReLU[17].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$764(.Z({ \dot_product_and_ReLU[17].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$765(.Z({ \dot_product_and_ReLU[17].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$766(.Z({ \dot_product_and_ReLU[17].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$767(.Z({ \dot_product_and_ReLU[17].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$768(.Z({ \dot_product_and_ReLU[17].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[17][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$769(.Z({ \dot_product_and_ReLU[16].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$770(.Z({ \dot_product_and_ReLU[16].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$771(.Z({ \dot_product_and_ReLU[16].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$772(.Z({ \dot_product_and_ReLU[16].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$773(.Z({ \dot_product_and_ReLU[16].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$774(.Z({ \dot_product_and_ReLU[16].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$775(.Z({ \dot_product_and_ReLU[16].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$776(.Z({ \dot_product_and_ReLU[16].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$777(.Z({ \dot_product_and_ReLU[16].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$778(.Z({ \dot_product_and_ReLU[16].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$779(.Z({ \dot_product_and_ReLU[16].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$780(.Z({ \dot_product_and_ReLU[16].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$781(.Z({ \dot_product_and_ReLU[16].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$782(.Z({ \dot_product_and_ReLU[16].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$783(.Z({ \dot_product_and_ReLU[16].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$784(.Z({ \dot_product_and_ReLU[16].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$785(.Z({ \dot_product_and_ReLU[16].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$786(.Z({ \dot_product_and_ReLU[16].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$787(.Z({ \dot_product_and_ReLU[16].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$788(.Z({ \dot_product_and_ReLU[16].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$789(.Z({ \dot_product_and_ReLU[16].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$790(.Z({ \dot_product_and_ReLU[16].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$791(.Z({ \dot_product_and_ReLU[16].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$792(.Z({ \dot_product_and_ReLU[16].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$793(.Z({ \dot_product_and_ReLU[16].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$794(.Z({ \dot_product_and_ReLU[16].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$795(.Z({ \dot_product_and_ReLU[16].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$796(.Z({ \dot_product_and_ReLU[16].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$797(.Z({ \dot_product_and_ReLU[16].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$798(.Z({ \dot_product_and_ReLU[16].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$799(.Z({ \dot_product_and_ReLU[16].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$800(.Z({ \dot_product_and_ReLU[16].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$801(.Z({ \dot_product_and_ReLU[16].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$802(.Z({ \dot_product_and_ReLU[16].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$803(.Z({ \dot_product_and_ReLU[16].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$804(.Z({ \dot_product_and_ReLU[16].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$805(.Z({ \dot_product_and_ReLU[16].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$806(.Z({ \dot_product_and_ReLU[16].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$807(.Z({ \dot_product_and_ReLU[16].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$808(.Z({ \dot_product_and_ReLU[16].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$809(.Z({ \dot_product_and_ReLU[16].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$810(.Z({ \dot_product_and_ReLU[16].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$811(.Z({ \dot_product_and_ReLU[16].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$812(.Z({ \dot_product_and_ReLU[16].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$813(.Z({ \dot_product_and_ReLU[16].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$814(.Z({ \dot_product_and_ReLU[16].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$815(.Z({ \dot_product_and_ReLU[16].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$816(.Z({ \dot_product_and_ReLU[16].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$817(.Z({ \dot_product_and_ReLU[16].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$818(.Z({ \dot_product_and_ReLU[16].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$819(.Z({ \dot_product_and_ReLU[16].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$820(.Z({ \dot_product_and_ReLU[16].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$821(.Z({ \dot_product_and_ReLU[16].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$822(.Z({ \dot_product_and_ReLU[16].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$823(.Z({ \dot_product_and_ReLU[16].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$824(.Z({ \dot_product_and_ReLU[16].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$825(.Z({ \dot_product_and_ReLU[16].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$826(.Z({ \dot_product_and_ReLU[16].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$827(.Z({ \dot_product_and_ReLU[16].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$828(.Z({ \dot_product_and_ReLU[16].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$829(.Z({ \dot_product_and_ReLU[16].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$830(.Z({ \dot_product_and_ReLU[16].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$831(.Z({ \dot_product_and_ReLU[16].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$832(.Z({ \dot_product_and_ReLU[16].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$833(.Z({ \dot_product_and_ReLU[16].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$834(.Z({ \dot_product_and_ReLU[16].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$835(.Z({ \dot_product_and_ReLU[16].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$836(.Z({ \dot_product_and_ReLU[16].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$837(.Z({ \dot_product_and_ReLU[16].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$838(.Z({ \dot_product_and_ReLU[16].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$839(.Z({ \dot_product_and_ReLU[16].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$840(.Z({ \dot_product_and_ReLU[16].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$841(.Z({ \dot_product_and_ReLU[16].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$842(.Z({ \dot_product_and_ReLU[16].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$843(.Z({ \dot_product_and_ReLU[16].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$844(.Z({ \dot_product_and_ReLU[16].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$845(.Z({ \dot_product_and_ReLU[16].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$846(.Z({ \dot_product_and_ReLU[16].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$847(.Z({ \dot_product_and_ReLU[16].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$848(.Z({ \dot_product_and_ReLU[16].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$849(.Z({ \dot_product_and_ReLU[16].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$850(.Z({ \dot_product_and_ReLU[16].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$851(.Z({ \dot_product_and_ReLU[16].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$852(.Z({ \dot_product_and_ReLU[16].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$853(.Z({ \dot_product_and_ReLU[16].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$854(.Z({ \dot_product_and_ReLU[16].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$855(.Z({ \dot_product_and_ReLU[16].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$856(.Z({ \dot_product_and_ReLU[16].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$857(.Z({ \dot_product_and_ReLU[16].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$858(.Z({ \dot_product_and_ReLU[16].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$859(.Z({ \dot_product_and_ReLU[16].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$860(.Z({ \dot_product_and_ReLU[16].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$861(.Z({ \dot_product_and_ReLU[16].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$862(.Z({ \dot_product_and_ReLU[16].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$863(.Z({ \dot_product_and_ReLU[16].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$864(.Z({ \dot_product_and_ReLU[16].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$865(.Z({ \dot_product_and_ReLU[16].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$866(.Z({ \dot_product_and_ReLU[16].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$867(.Z({ \dot_product_and_ReLU[16].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$868(.Z({ \dot_product_and_ReLU[16].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$869(.Z({ \dot_product_and_ReLU[16].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$870(.Z({ \dot_product_and_ReLU[16].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$871(.Z({ \dot_product_and_ReLU[16].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$872(.Z({ \dot_product_and_ReLU[16].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$873(.Z({ \dot_product_and_ReLU[16].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$874(.Z({ \dot_product_and_ReLU[16].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$875(.Z({ \dot_product_and_ReLU[16].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$876(.Z({ \dot_product_and_ReLU[16].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$877(.Z({ \dot_product_and_ReLU[16].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$878(.Z({ \dot_product_and_ReLU[16].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$879(.Z({ \dot_product_and_ReLU[16].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$880(.Z({ \dot_product_and_ReLU[16].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$881(.Z({ \dot_product_and_ReLU[16].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$882(.Z({ \dot_product_and_ReLU[16].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$883(.Z({ \dot_product_and_ReLU[16].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$884(.Z({ \dot_product_and_ReLU[16].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$885(.Z({ \dot_product_and_ReLU[16].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$886(.Z({ \dot_product_and_ReLU[16].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$887(.Z({ \dot_product_and_ReLU[16].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$888(.Z({ \dot_product_and_ReLU[16].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$889(.Z({ \dot_product_and_ReLU[16].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$890(.Z({ \dot_product_and_ReLU[16].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$891(.Z({ \dot_product_and_ReLU[16].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$892(.Z({ \dot_product_and_ReLU[16].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$893(.Z({ \dot_product_and_ReLU[16].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$894(.Z({ \dot_product_and_ReLU[16].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$895(.Z({ \dot_product_and_ReLU[16].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$896(.Z({ \dot_product_and_ReLU[16].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$897(.Z({ \dot_product_and_ReLU[16].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$898(.Z({ \dot_product_and_ReLU[16].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$899(.Z({ \dot_product_and_ReLU[16].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$900(.Z({ \dot_product_and_ReLU[16].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$901(.Z({ \dot_product_and_ReLU[16].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$902(.Z({ \dot_product_and_ReLU[16].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$903(.Z({ \dot_product_and_ReLU[16].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$904(.Z({ \dot_product_and_ReLU[16].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$905(.Z({ \dot_product_and_ReLU[16].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$906(.Z({ \dot_product_and_ReLU[16].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$907(.Z({ \dot_product_and_ReLU[16].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$908(.Z({ \dot_product_and_ReLU[16].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$909(.Z({ \dot_product_and_ReLU[16].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$910(.Z({ \dot_product_and_ReLU[16].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$911(.Z({ \dot_product_and_ReLU[16].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$912(.Z({ \dot_product_and_ReLU[16].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$913(.Z({ \dot_product_and_ReLU[16].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$914(.Z({ \dot_product_and_ReLU[16].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$915(.Z({ \dot_product_and_ReLU[16].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$916(.Z({ \dot_product_and_ReLU[16].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$917(.Z({ \dot_product_and_ReLU[16].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$918(.Z({ \dot_product_and_ReLU[16].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$919(.Z({ \dot_product_and_ReLU[16].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$920(.Z({ \dot_product_and_ReLU[16].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$921(.Z({ \dot_product_and_ReLU[16].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$922(.Z({ \dot_product_and_ReLU[16].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$923(.Z({ \dot_product_and_ReLU[16].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$924(.Z({ \dot_product_and_ReLU[16].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$925(.Z({ \dot_product_and_ReLU[16].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$926(.Z({ \dot_product_and_ReLU[16].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$927(.Z({ \dot_product_and_ReLU[16].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$928(.Z({ \dot_product_and_ReLU[16].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$929(.Z({ \dot_product_and_ReLU[16].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$930(.Z({ \dot_product_and_ReLU[16].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$931(.Z({ \dot_product_and_ReLU[16].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$932(.Z({ \dot_product_and_ReLU[16].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$933(.Z({ \dot_product_and_ReLU[16].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$934(.Z({ \dot_product_and_ReLU[16].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$935(.Z({ \dot_product_and_ReLU[16].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$936(.Z({ \dot_product_and_ReLU[16].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$937(.Z({ \dot_product_and_ReLU[16].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$938(.Z({ \dot_product_and_ReLU[16].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$939(.Z({ \dot_product_and_ReLU[16].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$940(.Z({ \dot_product_and_ReLU[16].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$941(.Z({ \dot_product_and_ReLU[16].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$942(.Z({ \dot_product_and_ReLU[16].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$943(.Z({ \dot_product_and_ReLU[16].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$944(.Z({ \dot_product_and_ReLU[16].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$945(.Z({ \dot_product_and_ReLU[16].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$946(.Z({ \dot_product_and_ReLU[16].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$947(.Z({ \dot_product_and_ReLU[16].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$948(.Z({ \dot_product_and_ReLU[16].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$949(.Z({ \dot_product_and_ReLU[16].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$950(.Z({ \dot_product_and_ReLU[16].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$951(.Z({ \dot_product_and_ReLU[16].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$952(.Z({ \dot_product_and_ReLU[16].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$953(.Z({ \dot_product_and_ReLU[16].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$954(.Z({ \dot_product_and_ReLU[16].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$955(.Z({ \dot_product_and_ReLU[16].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$956(.Z({ \dot_product_and_ReLU[16].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$957(.Z({ \dot_product_and_ReLU[16].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$958(.Z({ \dot_product_and_ReLU[16].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$959(.Z({ \dot_product_and_ReLU[16].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$960(.Z({ \dot_product_and_ReLU[16].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$961(.Z({ \dot_product_and_ReLU[16].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$962(.Z({ \dot_product_and_ReLU[16].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$963(.Z({ \dot_product_and_ReLU[16].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$964(.Z({ \dot_product_and_ReLU[16].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$965(.Z({ \dot_product_and_ReLU[16].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$966(.Z({ \dot_product_and_ReLU[16].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$967(.Z({ \dot_product_and_ReLU[16].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$968(.Z({ \dot_product_and_ReLU[16].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$969(.Z({ \dot_product_and_ReLU[16].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$970(.Z({ \dot_product_and_ReLU[16].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$971(.Z({ \dot_product_and_ReLU[16].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$972(.Z({ \dot_product_and_ReLU[16].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$973(.Z({ \dot_product_and_ReLU[16].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$974(.Z({ \dot_product_and_ReLU[16].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$975(.Z({ \dot_product_and_ReLU[16].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$976(.Z({ \dot_product_and_ReLU[16].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$977(.Z({ \dot_product_and_ReLU[16].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$978(.Z({ \dot_product_and_ReLU[16].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$979(.Z({ \dot_product_and_ReLU[16].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$980(.Z({ \dot_product_and_ReLU[16].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$981(.Z({ \dot_product_and_ReLU[16].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$982(.Z({ \dot_product_and_ReLU[16].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$983(.Z({ \dot_product_and_ReLU[16].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$984(.Z({ \dot_product_and_ReLU[16].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$985(.Z({ \dot_product_and_ReLU[16].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$986(.Z({ \dot_product_and_ReLU[16].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$987(.Z({ \dot_product_and_ReLU[16].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$988(.Z({ \dot_product_and_ReLU[16].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$989(.Z({ \dot_product_and_ReLU[16].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$990(.Z({ \dot_product_and_ReLU[16].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$991(.Z({ \dot_product_and_ReLU[16].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$992(.Z({ \dot_product_and_ReLU[16].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$993(.Z({ \dot_product_and_ReLU[16].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$994(.Z({ \dot_product_and_ReLU[16].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$995(.Z({ \dot_product_and_ReLU[16].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$996(.Z({ \dot_product_and_ReLU[16].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$997(.Z({ \dot_product_and_ReLU[16].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$998(.Z({ \dot_product_and_ReLU[16].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$999(.Z({ \dot_product_and_ReLU[16].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$1000(.Z({ \dot_product_and_ReLU[16].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$1001(.Z({ \dot_product_and_ReLU[16].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$1002(.Z({ \dot_product_and_ReLU[16].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$1003(.Z({ \dot_product_and_ReLU[16].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$1004(.Z({ \dot_product_and_ReLU[16].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$1005(.Z({ \dot_product_and_ReLU[16].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$1006(.Z({ \dot_product_and_ReLU[16].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$1007(.Z({ \dot_product_and_ReLU[16].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$1008(.Z({ \dot_product_and_ReLU[16].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$1009(.Z({ \dot_product_and_ReLU[16].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$1010(.Z({ \dot_product_and_ReLU[16].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$1011(.Z({ \dot_product_and_ReLU[16].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$1012(.Z({ \dot_product_and_ReLU[16].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$1013(.Z({ \dot_product_and_ReLU[16].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$1014(.Z({ \dot_product_and_ReLU[16].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$1015(.Z({ \dot_product_and_ReLU[16].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$1016(.Z({ \dot_product_and_ReLU[16].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$1017(.Z({ \dot_product_and_ReLU[16].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$1018(.Z({ \dot_product_and_ReLU[16].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$1019(.Z({ \dot_product_and_ReLU[16].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$1020(.Z({ \dot_product_and_ReLU[16].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$1021(.Z({ \dot_product_and_ReLU[16].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$1022(.Z({ \dot_product_and_ReLU[16].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$1023(.Z({ \dot_product_and_ReLU[16].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$1024(.Z({ \dot_product_and_ReLU[16].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[16][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$1025(.Z({ \dot_product_and_ReLU[15].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$1026(.Z({ \dot_product_and_ReLU[15].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$1027(.Z({ \dot_product_and_ReLU[15].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$1028(.Z({ \dot_product_and_ReLU[15].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$1029(.Z({ \dot_product_and_ReLU[15].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$1030(.Z({ \dot_product_and_ReLU[15].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$1031(.Z({ \dot_product_and_ReLU[15].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$1032(.Z({ \dot_product_and_ReLU[15].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$1033(.Z({ \dot_product_and_ReLU[15].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$1034(.Z({ \dot_product_and_ReLU[15].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$1035(.Z({ \dot_product_and_ReLU[15].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$1036(.Z({ \dot_product_and_ReLU[15].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$1037(.Z({ \dot_product_and_ReLU[15].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$1038(.Z({ \dot_product_and_ReLU[15].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$1039(.Z({ \dot_product_and_ReLU[15].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$1040(.Z({ \dot_product_and_ReLU[15].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$1041(.Z({ \dot_product_and_ReLU[15].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$1042(.Z({ \dot_product_and_ReLU[15].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$1043(.Z({ \dot_product_and_ReLU[15].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$1044(.Z({ \dot_product_and_ReLU[15].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$1045(.Z({ \dot_product_and_ReLU[15].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$1046(.Z({ \dot_product_and_ReLU[15].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$1047(.Z({ \dot_product_and_ReLU[15].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$1048(.Z({ \dot_product_and_ReLU[15].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$1049(.Z({ \dot_product_and_ReLU[15].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$1050(.Z({ \dot_product_and_ReLU[15].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$1051(.Z({ \dot_product_and_ReLU[15].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$1052(.Z({ \dot_product_and_ReLU[15].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$1053(.Z({ \dot_product_and_ReLU[15].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$1054(.Z({ \dot_product_and_ReLU[15].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$1055(.Z({ \dot_product_and_ReLU[15].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$1056(.Z({ \dot_product_and_ReLU[15].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$1057(.Z({ \dot_product_and_ReLU[15].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$1058(.Z({ \dot_product_and_ReLU[15].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$1059(.Z({ \dot_product_and_ReLU[15].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$1060(.Z({ \dot_product_and_ReLU[15].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$1061(.Z({ \dot_product_and_ReLU[15].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$1062(.Z({ \dot_product_and_ReLU[15].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$1063(.Z({ \dot_product_and_ReLU[15].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$1064(.Z({ \dot_product_and_ReLU[15].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$1065(.Z({ \dot_product_and_ReLU[15].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$1066(.Z({ \dot_product_and_ReLU[15].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$1067(.Z({ \dot_product_and_ReLU[15].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$1068(.Z({ \dot_product_and_ReLU[15].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$1069(.Z({ \dot_product_and_ReLU[15].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$1070(.Z({ \dot_product_and_ReLU[15].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$1071(.Z({ \dot_product_and_ReLU[15].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$1072(.Z({ \dot_product_and_ReLU[15].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$1073(.Z({ \dot_product_and_ReLU[15].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$1074(.Z({ \dot_product_and_ReLU[15].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$1075(.Z({ \dot_product_and_ReLU[15].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$1076(.Z({ \dot_product_and_ReLU[15].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$1077(.Z({ \dot_product_and_ReLU[15].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$1078(.Z({ \dot_product_and_ReLU[15].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$1079(.Z({ \dot_product_and_ReLU[15].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$1080(.Z({ \dot_product_and_ReLU[15].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$1081(.Z({ \dot_product_and_ReLU[15].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$1082(.Z({ \dot_product_and_ReLU[15].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$1083(.Z({ \dot_product_and_ReLU[15].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$1084(.Z({ \dot_product_and_ReLU[15].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$1085(.Z({ \dot_product_and_ReLU[15].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$1086(.Z({ \dot_product_and_ReLU[15].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$1087(.Z({ \dot_product_and_ReLU[15].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$1088(.Z({ \dot_product_and_ReLU[15].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$1089(.Z({ \dot_product_and_ReLU[15].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$1090(.Z({ \dot_product_and_ReLU[15].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$1091(.Z({ \dot_product_and_ReLU[15].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$1092(.Z({ \dot_product_and_ReLU[15].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$1093(.Z({ \dot_product_and_ReLU[15].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$1094(.Z({ \dot_product_and_ReLU[15].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$1095(.Z({ \dot_product_and_ReLU[15].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$1096(.Z({ \dot_product_and_ReLU[15].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$1097(.Z({ \dot_product_and_ReLU[15].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$1098(.Z({ \dot_product_and_ReLU[15].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$1099(.Z({ \dot_product_and_ReLU[15].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$1100(.Z({ \dot_product_and_ReLU[15].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$1101(.Z({ \dot_product_and_ReLU[15].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$1102(.Z({ \dot_product_and_ReLU[15].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$1103(.Z({ \dot_product_and_ReLU[15].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$1104(.Z({ \dot_product_and_ReLU[15].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$1105(.Z({ \dot_product_and_ReLU[15].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$1106(.Z({ \dot_product_and_ReLU[15].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$1107(.Z({ \dot_product_and_ReLU[15].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$1108(.Z({ \dot_product_and_ReLU[15].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$1109(.Z({ \dot_product_and_ReLU[15].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$1110(.Z({ \dot_product_and_ReLU[15].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$1111(.Z({ \dot_product_and_ReLU[15].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$1112(.Z({ \dot_product_and_ReLU[15].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$1113(.Z({ \dot_product_and_ReLU[15].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$1114(.Z({ \dot_product_and_ReLU[15].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$1115(.Z({ \dot_product_and_ReLU[15].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$1116(.Z({ \dot_product_and_ReLU[15].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$1117(.Z({ \dot_product_and_ReLU[15].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$1118(.Z({ \dot_product_and_ReLU[15].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$1119(.Z({ \dot_product_and_ReLU[15].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$1120(.Z({ \dot_product_and_ReLU[15].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$1121(.Z({ \dot_product_and_ReLU[15].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$1122(.Z({ \dot_product_and_ReLU[15].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$1123(.Z({ \dot_product_and_ReLU[15].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$1124(.Z({ \dot_product_and_ReLU[15].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$1125(.Z({ \dot_product_and_ReLU[15].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$1126(.Z({ \dot_product_and_ReLU[15].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$1127(.Z({ \dot_product_and_ReLU[15].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$1128(.Z({ \dot_product_and_ReLU[15].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$1129(.Z({ \dot_product_and_ReLU[15].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$1130(.Z({ \dot_product_and_ReLU[15].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$1131(.Z({ \dot_product_and_ReLU[15].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$1132(.Z({ \dot_product_and_ReLU[15].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$1133(.Z({ \dot_product_and_ReLU[15].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$1134(.Z({ \dot_product_and_ReLU[15].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$1135(.Z({ \dot_product_and_ReLU[15].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$1136(.Z({ \dot_product_and_ReLU[15].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$1137(.Z({ \dot_product_and_ReLU[15].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$1138(.Z({ \dot_product_and_ReLU[15].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$1139(.Z({ \dot_product_and_ReLU[15].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$1140(.Z({ \dot_product_and_ReLU[15].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$1141(.Z({ \dot_product_and_ReLU[15].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$1142(.Z({ \dot_product_and_ReLU[15].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$1143(.Z({ \dot_product_and_ReLU[15].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$1144(.Z({ \dot_product_and_ReLU[15].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$1145(.Z({ \dot_product_and_ReLU[15].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$1146(.Z({ \dot_product_and_ReLU[15].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$1147(.Z({ \dot_product_and_ReLU[15].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$1148(.Z({ \dot_product_and_ReLU[15].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$1149(.Z({ \dot_product_and_ReLU[15].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$1150(.Z({ \dot_product_and_ReLU[15].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$1151(.Z({ \dot_product_and_ReLU[15].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$1152(.Z({ \dot_product_and_ReLU[15].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$1153(.Z({ \dot_product_and_ReLU[15].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$1154(.Z({ \dot_product_and_ReLU[15].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$1155(.Z({ \dot_product_and_ReLU[15].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$1156(.Z({ \dot_product_and_ReLU[15].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$1157(.Z({ \dot_product_and_ReLU[15].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$1158(.Z({ \dot_product_and_ReLU[15].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$1159(.Z({ \dot_product_and_ReLU[15].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$1160(.Z({ \dot_product_and_ReLU[15].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$1161(.Z({ \dot_product_and_ReLU[15].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$1162(.Z({ \dot_product_and_ReLU[15].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$1163(.Z({ \dot_product_and_ReLU[15].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$1164(.Z({ \dot_product_and_ReLU[15].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$1165(.Z({ \dot_product_and_ReLU[15].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$1166(.Z({ \dot_product_and_ReLU[15].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$1167(.Z({ \dot_product_and_ReLU[15].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$1168(.Z({ \dot_product_and_ReLU[15].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$1169(.Z({ \dot_product_and_ReLU[15].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$1170(.Z({ \dot_product_and_ReLU[15].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$1171(.Z({ \dot_product_and_ReLU[15].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$1172(.Z({ \dot_product_and_ReLU[15].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$1173(.Z({ \dot_product_and_ReLU[15].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$1174(.Z({ \dot_product_and_ReLU[15].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$1175(.Z({ \dot_product_and_ReLU[15].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$1176(.Z({ \dot_product_and_ReLU[15].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$1177(.Z({ \dot_product_and_ReLU[15].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$1178(.Z({ \dot_product_and_ReLU[15].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$1179(.Z({ \dot_product_and_ReLU[15].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$1180(.Z({ \dot_product_and_ReLU[15].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$1181(.Z({ \dot_product_and_ReLU[15].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$1182(.Z({ \dot_product_and_ReLU[15].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$1183(.Z({ \dot_product_and_ReLU[15].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$1184(.Z({ \dot_product_and_ReLU[15].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$1185(.Z({ \dot_product_and_ReLU[15].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$1186(.Z({ \dot_product_and_ReLU[15].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$1187(.Z({ \dot_product_and_ReLU[15].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$1188(.Z({ \dot_product_and_ReLU[15].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$1189(.Z({ \dot_product_and_ReLU[15].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$1190(.Z({ \dot_product_and_ReLU[15].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$1191(.Z({ \dot_product_and_ReLU[15].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$1192(.Z({ \dot_product_and_ReLU[15].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$1193(.Z({ \dot_product_and_ReLU[15].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$1194(.Z({ \dot_product_and_ReLU[15].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$1195(.Z({ \dot_product_and_ReLU[15].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$1196(.Z({ \dot_product_and_ReLU[15].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$1197(.Z({ \dot_product_and_ReLU[15].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$1198(.Z({ \dot_product_and_ReLU[15].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$1199(.Z({ \dot_product_and_ReLU[15].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$1200(.Z({ \dot_product_and_ReLU[15].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$1201(.Z({ \dot_product_and_ReLU[15].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$1202(.Z({ \dot_product_and_ReLU[15].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$1203(.Z({ \dot_product_and_ReLU[15].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$1204(.Z({ \dot_product_and_ReLU[15].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$1205(.Z({ \dot_product_and_ReLU[15].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$1206(.Z({ \dot_product_and_ReLU[15].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$1207(.Z({ \dot_product_and_ReLU[15].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$1208(.Z({ \dot_product_and_ReLU[15].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$1209(.Z({ \dot_product_and_ReLU[15].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$1210(.Z({ \dot_product_and_ReLU[15].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$1211(.Z({ \dot_product_and_ReLU[15].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$1212(.Z({ \dot_product_and_ReLU[15].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$1213(.Z({ \dot_product_and_ReLU[15].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$1214(.Z({ \dot_product_and_ReLU[15].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$1215(.Z({ \dot_product_and_ReLU[15].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$1216(.Z({ \dot_product_and_ReLU[15].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$1217(.Z({ \dot_product_and_ReLU[15].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$1218(.Z({ \dot_product_and_ReLU[15].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$1219(.Z({ \dot_product_and_ReLU[15].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$1220(.Z({ \dot_product_and_ReLU[15].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$1221(.Z({ \dot_product_and_ReLU[15].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$1222(.Z({ \dot_product_and_ReLU[15].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$1223(.Z({ \dot_product_and_ReLU[15].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$1224(.Z({ \dot_product_and_ReLU[15].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$1225(.Z({ \dot_product_and_ReLU[15].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$1226(.Z({ \dot_product_and_ReLU[15].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$1227(.Z({ \dot_product_and_ReLU[15].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$1228(.Z({ \dot_product_and_ReLU[15].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$1229(.Z({ \dot_product_and_ReLU[15].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$1230(.Z({ \dot_product_and_ReLU[15].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$1231(.Z({ \dot_product_and_ReLU[15].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$1232(.Z({ \dot_product_and_ReLU[15].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$1233(.Z({ \dot_product_and_ReLU[15].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$1234(.Z({ \dot_product_and_ReLU[15].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$1235(.Z({ \dot_product_and_ReLU[15].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$1236(.Z({ \dot_product_and_ReLU[15].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$1237(.Z({ \dot_product_and_ReLU[15].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$1238(.Z({ \dot_product_and_ReLU[15].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$1239(.Z({ \dot_product_and_ReLU[15].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$1240(.Z({ \dot_product_and_ReLU[15].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$1241(.Z({ \dot_product_and_ReLU[15].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$1242(.Z({ \dot_product_and_ReLU[15].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$1243(.Z({ \dot_product_and_ReLU[15].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$1244(.Z({ \dot_product_and_ReLU[15].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$1245(.Z({ \dot_product_and_ReLU[15].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$1246(.Z({ \dot_product_and_ReLU[15].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$1247(.Z({ \dot_product_and_ReLU[15].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$1248(.Z({ \dot_product_and_ReLU[15].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$1249(.Z({ \dot_product_and_ReLU[15].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$1250(.Z({ \dot_product_and_ReLU[15].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$1251(.Z({ \dot_product_and_ReLU[15].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$1252(.Z({ \dot_product_and_ReLU[15].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$1253(.Z({ \dot_product_and_ReLU[15].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$1254(.Z({ \dot_product_and_ReLU[15].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$1255(.Z({ \dot_product_and_ReLU[15].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$1256(.Z({ \dot_product_and_ReLU[15].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$1257(.Z({ \dot_product_and_ReLU[15].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$1258(.Z({ \dot_product_and_ReLU[15].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$1259(.Z({ \dot_product_and_ReLU[15].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$1260(.Z({ \dot_product_and_ReLU[15].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$1261(.Z({ \dot_product_and_ReLU[15].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$1262(.Z({ \dot_product_and_ReLU[15].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$1263(.Z({ \dot_product_and_ReLU[15].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$1264(.Z({ \dot_product_and_ReLU[15].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$1265(.Z({ \dot_product_and_ReLU[15].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$1266(.Z({ \dot_product_and_ReLU[15].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$1267(.Z({ \dot_product_and_ReLU[15].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$1268(.Z({ \dot_product_and_ReLU[15].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$1269(.Z({ \dot_product_and_ReLU[15].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$1270(.Z({ \dot_product_and_ReLU[15].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$1271(.Z({ \dot_product_and_ReLU[15].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$1272(.Z({ \dot_product_and_ReLU[15].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$1273(.Z({ \dot_product_and_ReLU[15].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$1274(.Z({ \dot_product_and_ReLU[15].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$1275(.Z({ \dot_product_and_ReLU[15].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$1276(.Z({ \dot_product_and_ReLU[15].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$1277(.Z({ \dot_product_and_ReLU[15].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$1278(.Z({ \dot_product_and_ReLU[15].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$1279(.Z({ \dot_product_and_ReLU[15].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$1280(.Z({ \dot_product_and_ReLU[15].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[15][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$1281(.Z({ \dot_product_and_ReLU[14].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$1282(.Z({ \dot_product_and_ReLU[14].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$1283(.Z({ \dot_product_and_ReLU[14].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$1284(.Z({ \dot_product_and_ReLU[14].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$1285(.Z({ \dot_product_and_ReLU[14].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$1286(.Z({ \dot_product_and_ReLU[14].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$1287(.Z({ \dot_product_and_ReLU[14].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$1288(.Z({ \dot_product_and_ReLU[14].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$1289(.Z({ \dot_product_and_ReLU[14].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$1290(.Z({ \dot_product_and_ReLU[14].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$1291(.Z({ \dot_product_and_ReLU[14].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$1292(.Z({ \dot_product_and_ReLU[14].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$1293(.Z({ \dot_product_and_ReLU[14].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$1294(.Z({ \dot_product_and_ReLU[14].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$1295(.Z({ \dot_product_and_ReLU[14].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$1296(.Z({ \dot_product_and_ReLU[14].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$1297(.Z({ \dot_product_and_ReLU[14].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$1298(.Z({ \dot_product_and_ReLU[14].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$1299(.Z({ \dot_product_and_ReLU[14].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$1300(.Z({ \dot_product_and_ReLU[14].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$1301(.Z({ \dot_product_and_ReLU[14].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$1302(.Z({ \dot_product_and_ReLU[14].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$1303(.Z({ \dot_product_and_ReLU[14].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$1304(.Z({ \dot_product_and_ReLU[14].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$1305(.Z({ \dot_product_and_ReLU[14].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$1306(.Z({ \dot_product_and_ReLU[14].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$1307(.Z({ \dot_product_and_ReLU[14].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$1308(.Z({ \dot_product_and_ReLU[14].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$1309(.Z({ \dot_product_and_ReLU[14].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$1310(.Z({ \dot_product_and_ReLU[14].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$1311(.Z({ \dot_product_and_ReLU[14].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$1312(.Z({ \dot_product_and_ReLU[14].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$1313(.Z({ \dot_product_and_ReLU[14].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$1314(.Z({ \dot_product_and_ReLU[14].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$1315(.Z({ \dot_product_and_ReLU[14].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$1316(.Z({ \dot_product_and_ReLU[14].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$1317(.Z({ \dot_product_and_ReLU[14].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$1318(.Z({ \dot_product_and_ReLU[14].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$1319(.Z({ \dot_product_and_ReLU[14].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$1320(.Z({ \dot_product_and_ReLU[14].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$1321(.Z({ \dot_product_and_ReLU[14].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$1322(.Z({ \dot_product_and_ReLU[14].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$1323(.Z({ \dot_product_and_ReLU[14].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$1324(.Z({ \dot_product_and_ReLU[14].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$1325(.Z({ \dot_product_and_ReLU[14].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$1326(.Z({ \dot_product_and_ReLU[14].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$1327(.Z({ \dot_product_and_ReLU[14].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$1328(.Z({ \dot_product_and_ReLU[14].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$1329(.Z({ \dot_product_and_ReLU[14].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$1330(.Z({ \dot_product_and_ReLU[14].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$1331(.Z({ \dot_product_and_ReLU[14].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$1332(.Z({ \dot_product_and_ReLU[14].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$1333(.Z({ \dot_product_and_ReLU[14].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$1334(.Z({ \dot_product_and_ReLU[14].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$1335(.Z({ \dot_product_and_ReLU[14].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$1336(.Z({ \dot_product_and_ReLU[14].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$1337(.Z({ \dot_product_and_ReLU[14].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$1338(.Z({ \dot_product_and_ReLU[14].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$1339(.Z({ \dot_product_and_ReLU[14].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$1340(.Z({ \dot_product_and_ReLU[14].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$1341(.Z({ \dot_product_and_ReLU[14].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$1342(.Z({ \dot_product_and_ReLU[14].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$1343(.Z({ \dot_product_and_ReLU[14].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$1344(.Z({ \dot_product_and_ReLU[14].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$1345(.Z({ \dot_product_and_ReLU[14].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$1346(.Z({ \dot_product_and_ReLU[14].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$1347(.Z({ \dot_product_and_ReLU[14].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$1348(.Z({ \dot_product_and_ReLU[14].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$1349(.Z({ \dot_product_and_ReLU[14].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$1350(.Z({ \dot_product_and_ReLU[14].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$1351(.Z({ \dot_product_and_ReLU[14].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$1352(.Z({ \dot_product_and_ReLU[14].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$1353(.Z({ \dot_product_and_ReLU[14].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$1354(.Z({ \dot_product_and_ReLU[14].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$1355(.Z({ \dot_product_and_ReLU[14].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$1356(.Z({ \dot_product_and_ReLU[14].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$1357(.Z({ \dot_product_and_ReLU[14].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$1358(.Z({ \dot_product_and_ReLU[14].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$1359(.Z({ \dot_product_and_ReLU[14].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$1360(.Z({ \dot_product_and_ReLU[14].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$1361(.Z({ \dot_product_and_ReLU[14].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$1362(.Z({ \dot_product_and_ReLU[14].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$1363(.Z({ \dot_product_and_ReLU[14].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$1364(.Z({ \dot_product_and_ReLU[14].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$1365(.Z({ \dot_product_and_ReLU[14].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$1366(.Z({ \dot_product_and_ReLU[14].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$1367(.Z({ \dot_product_and_ReLU[14].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$1368(.Z({ \dot_product_and_ReLU[14].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$1369(.Z({ \dot_product_and_ReLU[14].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$1370(.Z({ \dot_product_and_ReLU[14].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$1371(.Z({ \dot_product_and_ReLU[14].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$1372(.Z({ \dot_product_and_ReLU[14].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$1373(.Z({ \dot_product_and_ReLU[14].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$1374(.Z({ \dot_product_and_ReLU[14].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$1375(.Z({ \dot_product_and_ReLU[14].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$1376(.Z({ \dot_product_and_ReLU[14].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$1377(.Z({ \dot_product_and_ReLU[14].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$1378(.Z({ \dot_product_and_ReLU[14].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$1379(.Z({ \dot_product_and_ReLU[14].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$1380(.Z({ \dot_product_and_ReLU[14].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$1381(.Z({ \dot_product_and_ReLU[14].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$1382(.Z({ \dot_product_and_ReLU[14].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$1383(.Z({ \dot_product_and_ReLU[14].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$1384(.Z({ \dot_product_and_ReLU[14].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$1385(.Z({ \dot_product_and_ReLU[14].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$1386(.Z({ \dot_product_and_ReLU[14].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$1387(.Z({ \dot_product_and_ReLU[14].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$1388(.Z({ \dot_product_and_ReLU[14].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$1389(.Z({ \dot_product_and_ReLU[14].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$1390(.Z({ \dot_product_and_ReLU[14].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$1391(.Z({ \dot_product_and_ReLU[14].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$1392(.Z({ \dot_product_and_ReLU[14].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$1393(.Z({ \dot_product_and_ReLU[14].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$1394(.Z({ \dot_product_and_ReLU[14].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$1395(.Z({ \dot_product_and_ReLU[14].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$1396(.Z({ \dot_product_and_ReLU[14].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$1397(.Z({ \dot_product_and_ReLU[14].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$1398(.Z({ \dot_product_and_ReLU[14].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$1399(.Z({ \dot_product_and_ReLU[14].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$1400(.Z({ \dot_product_and_ReLU[14].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$1401(.Z({ \dot_product_and_ReLU[14].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$1402(.Z({ \dot_product_and_ReLU[14].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$1403(.Z({ \dot_product_and_ReLU[14].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$1404(.Z({ \dot_product_and_ReLU[14].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$1405(.Z({ \dot_product_and_ReLU[14].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$1406(.Z({ \dot_product_and_ReLU[14].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$1407(.Z({ \dot_product_and_ReLU[14].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$1408(.Z({ \dot_product_and_ReLU[14].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$1409(.Z({ \dot_product_and_ReLU[14].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$1410(.Z({ \dot_product_and_ReLU[14].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$1411(.Z({ \dot_product_and_ReLU[14].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$1412(.Z({ \dot_product_and_ReLU[14].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$1413(.Z({ \dot_product_and_ReLU[14].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$1414(.Z({ \dot_product_and_ReLU[14].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$1415(.Z({ \dot_product_and_ReLU[14].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$1416(.Z({ \dot_product_and_ReLU[14].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$1417(.Z({ \dot_product_and_ReLU[14].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$1418(.Z({ \dot_product_and_ReLU[14].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$1419(.Z({ \dot_product_and_ReLU[14].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$1420(.Z({ \dot_product_and_ReLU[14].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$1421(.Z({ \dot_product_and_ReLU[14].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$1422(.Z({ \dot_product_and_ReLU[14].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$1423(.Z({ \dot_product_and_ReLU[14].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$1424(.Z({ \dot_product_and_ReLU[14].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$1425(.Z({ \dot_product_and_ReLU[14].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$1426(.Z({ \dot_product_and_ReLU[14].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$1427(.Z({ \dot_product_and_ReLU[14].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$1428(.Z({ \dot_product_and_ReLU[14].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$1429(.Z({ \dot_product_and_ReLU[14].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$1430(.Z({ \dot_product_and_ReLU[14].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$1431(.Z({ \dot_product_and_ReLU[14].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$1432(.Z({ \dot_product_and_ReLU[14].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$1433(.Z({ \dot_product_and_ReLU[14].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$1434(.Z({ \dot_product_and_ReLU[14].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$1435(.Z({ \dot_product_and_ReLU[14].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$1436(.Z({ \dot_product_and_ReLU[14].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$1437(.Z({ \dot_product_and_ReLU[14].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$1438(.Z({ \dot_product_and_ReLU[14].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$1439(.Z({ \dot_product_and_ReLU[14].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$1440(.Z({ \dot_product_and_ReLU[14].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$1441(.Z({ \dot_product_and_ReLU[14].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$1442(.Z({ \dot_product_and_ReLU[14].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$1443(.Z({ \dot_product_and_ReLU[14].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$1444(.Z({ \dot_product_and_ReLU[14].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$1445(.Z({ \dot_product_and_ReLU[14].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$1446(.Z({ \dot_product_and_ReLU[14].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$1447(.Z({ \dot_product_and_ReLU[14].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$1448(.Z({ \dot_product_and_ReLU[14].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$1449(.Z({ \dot_product_and_ReLU[14].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$1450(.Z({ \dot_product_and_ReLU[14].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$1451(.Z({ \dot_product_and_ReLU[14].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$1452(.Z({ \dot_product_and_ReLU[14].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$1453(.Z({ \dot_product_and_ReLU[14].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$1454(.Z({ \dot_product_and_ReLU[14].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$1455(.Z({ \dot_product_and_ReLU[14].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$1456(.Z({ \dot_product_and_ReLU[14].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$1457(.Z({ \dot_product_and_ReLU[14].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$1458(.Z({ \dot_product_and_ReLU[14].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$1459(.Z({ \dot_product_and_ReLU[14].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$1460(.Z({ \dot_product_and_ReLU[14].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$1461(.Z({ \dot_product_and_ReLU[14].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$1462(.Z({ \dot_product_and_ReLU[14].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$1463(.Z({ \dot_product_and_ReLU[14].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$1464(.Z({ \dot_product_and_ReLU[14].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$1465(.Z({ \dot_product_and_ReLU[14].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$1466(.Z({ \dot_product_and_ReLU[14].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$1467(.Z({ \dot_product_and_ReLU[14].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$1468(.Z({ \dot_product_and_ReLU[14].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$1469(.Z({ \dot_product_and_ReLU[14].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$1470(.Z({ \dot_product_and_ReLU[14].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$1471(.Z({ \dot_product_and_ReLU[14].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$1472(.Z({ \dot_product_and_ReLU[14].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$1473(.Z({ \dot_product_and_ReLU[14].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$1474(.Z({ \dot_product_and_ReLU[14].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$1475(.Z({ \dot_product_and_ReLU[14].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$1476(.Z({ \dot_product_and_ReLU[14].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$1477(.Z({ \dot_product_and_ReLU[14].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$1478(.Z({ \dot_product_and_ReLU[14].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$1479(.Z({ \dot_product_and_ReLU[14].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$1480(.Z({ \dot_product_and_ReLU[14].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$1481(.Z({ \dot_product_and_ReLU[14].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$1482(.Z({ \dot_product_and_ReLU[14].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$1483(.Z({ \dot_product_and_ReLU[14].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$1484(.Z({ \dot_product_and_ReLU[14].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$1485(.Z({ \dot_product_and_ReLU[14].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$1486(.Z({ \dot_product_and_ReLU[14].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$1487(.Z({ \dot_product_and_ReLU[14].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$1488(.Z({ \dot_product_and_ReLU[14].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$1489(.Z({ \dot_product_and_ReLU[14].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$1490(.Z({ \dot_product_and_ReLU[14].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$1491(.Z({ \dot_product_and_ReLU[14].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$1492(.Z({ \dot_product_and_ReLU[14].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$1493(.Z({ \dot_product_and_ReLU[14].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$1494(.Z({ \dot_product_and_ReLU[14].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$1495(.Z({ \dot_product_and_ReLU[14].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$1496(.Z({ \dot_product_and_ReLU[14].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$1497(.Z({ \dot_product_and_ReLU[14].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$1498(.Z({ \dot_product_and_ReLU[14].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$1499(.Z({ \dot_product_and_ReLU[14].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$1500(.Z({ \dot_product_and_ReLU[14].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$1501(.Z({ \dot_product_and_ReLU[14].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$1502(.Z({ \dot_product_and_ReLU[14].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$1503(.Z({ \dot_product_and_ReLU[14].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$1504(.Z({ \dot_product_and_ReLU[14].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$1505(.Z({ \dot_product_and_ReLU[14].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$1506(.Z({ \dot_product_and_ReLU[14].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$1507(.Z({ \dot_product_and_ReLU[14].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$1508(.Z({ \dot_product_and_ReLU[14].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$1509(.Z({ \dot_product_and_ReLU[14].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$1510(.Z({ \dot_product_and_ReLU[14].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$1511(.Z({ \dot_product_and_ReLU[14].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$1512(.Z({ \dot_product_and_ReLU[14].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$1513(.Z({ \dot_product_and_ReLU[14].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$1514(.Z({ \dot_product_and_ReLU[14].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$1515(.Z({ \dot_product_and_ReLU[14].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$1516(.Z({ \dot_product_and_ReLU[14].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$1517(.Z({ \dot_product_and_ReLU[14].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$1518(.Z({ \dot_product_and_ReLU[14].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$1519(.Z({ \dot_product_and_ReLU[14].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$1520(.Z({ \dot_product_and_ReLU[14].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$1521(.Z({ \dot_product_and_ReLU[14].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$1522(.Z({ \dot_product_and_ReLU[14].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$1523(.Z({ \dot_product_and_ReLU[14].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$1524(.Z({ \dot_product_and_ReLU[14].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$1525(.Z({ \dot_product_and_ReLU[14].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$1526(.Z({ \dot_product_and_ReLU[14].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$1527(.Z({ \dot_product_and_ReLU[14].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$1528(.Z({ \dot_product_and_ReLU[14].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$1529(.Z({ \dot_product_and_ReLU[14].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$1530(.Z({ \dot_product_and_ReLU[14].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$1531(.Z({ \dot_product_and_ReLU[14].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$1532(.Z({ \dot_product_and_ReLU[14].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$1533(.Z({ \dot_product_and_ReLU[14].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$1534(.Z({ \dot_product_and_ReLU[14].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$1535(.Z({ \dot_product_and_ReLU[14].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$1536(.Z({ \dot_product_and_ReLU[14].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[14][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$1537(.Z({ \dot_product_and_ReLU[13].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$1538(.Z({ \dot_product_and_ReLU[13].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$1539(.Z({ \dot_product_and_ReLU[13].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$1540(.Z({ \dot_product_and_ReLU[13].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$1541(.Z({ \dot_product_and_ReLU[13].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$1542(.Z({ \dot_product_and_ReLU[13].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$1543(.Z({ \dot_product_and_ReLU[13].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$1544(.Z({ \dot_product_and_ReLU[13].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$1545(.Z({ \dot_product_and_ReLU[13].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$1546(.Z({ \dot_product_and_ReLU[13].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$1547(.Z({ \dot_product_and_ReLU[13].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$1548(.Z({ \dot_product_and_ReLU[13].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$1549(.Z({ \dot_product_and_ReLU[13].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$1550(.Z({ \dot_product_and_ReLU[13].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$1551(.Z({ \dot_product_and_ReLU[13].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$1552(.Z({ \dot_product_and_ReLU[13].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$1553(.Z({ \dot_product_and_ReLU[13].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$1554(.Z({ \dot_product_and_ReLU[13].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$1555(.Z({ \dot_product_and_ReLU[13].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$1556(.Z({ \dot_product_and_ReLU[13].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$1557(.Z({ \dot_product_and_ReLU[13].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$1558(.Z({ \dot_product_and_ReLU[13].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$1559(.Z({ \dot_product_and_ReLU[13].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$1560(.Z({ \dot_product_and_ReLU[13].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$1561(.Z({ \dot_product_and_ReLU[13].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$1562(.Z({ \dot_product_and_ReLU[13].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$1563(.Z({ \dot_product_and_ReLU[13].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$1564(.Z({ \dot_product_and_ReLU[13].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$1565(.Z({ \dot_product_and_ReLU[13].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$1566(.Z({ \dot_product_and_ReLU[13].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$1567(.Z({ \dot_product_and_ReLU[13].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$1568(.Z({ \dot_product_and_ReLU[13].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$1569(.Z({ \dot_product_and_ReLU[13].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$1570(.Z({ \dot_product_and_ReLU[13].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$1571(.Z({ \dot_product_and_ReLU[13].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$1572(.Z({ \dot_product_and_ReLU[13].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$1573(.Z({ \dot_product_and_ReLU[13].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$1574(.Z({ \dot_product_and_ReLU[13].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$1575(.Z({ \dot_product_and_ReLU[13].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$1576(.Z({ \dot_product_and_ReLU[13].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$1577(.Z({ \dot_product_and_ReLU[13].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$1578(.Z({ \dot_product_and_ReLU[13].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$1579(.Z({ \dot_product_and_ReLU[13].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$1580(.Z({ \dot_product_and_ReLU[13].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$1581(.Z({ \dot_product_and_ReLU[13].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$1582(.Z({ \dot_product_and_ReLU[13].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$1583(.Z({ \dot_product_and_ReLU[13].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$1584(.Z({ \dot_product_and_ReLU[13].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$1585(.Z({ \dot_product_and_ReLU[13].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$1586(.Z({ \dot_product_and_ReLU[13].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$1587(.Z({ \dot_product_and_ReLU[13].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$1588(.Z({ \dot_product_and_ReLU[13].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$1589(.Z({ \dot_product_and_ReLU[13].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$1590(.Z({ \dot_product_and_ReLU[13].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$1591(.Z({ \dot_product_and_ReLU[13].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$1592(.Z({ \dot_product_and_ReLU[13].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$1593(.Z({ \dot_product_and_ReLU[13].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$1594(.Z({ \dot_product_and_ReLU[13].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$1595(.Z({ \dot_product_and_ReLU[13].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$1596(.Z({ \dot_product_and_ReLU[13].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$1597(.Z({ \dot_product_and_ReLU[13].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$1598(.Z({ \dot_product_and_ReLU[13].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$1599(.Z({ \dot_product_and_ReLU[13].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$1600(.Z({ \dot_product_and_ReLU[13].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$1601(.Z({ \dot_product_and_ReLU[13].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$1602(.Z({ \dot_product_and_ReLU[13].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$1603(.Z({ \dot_product_and_ReLU[13].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$1604(.Z({ \dot_product_and_ReLU[13].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$1605(.Z({ \dot_product_and_ReLU[13].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$1606(.Z({ \dot_product_and_ReLU[13].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$1607(.Z({ \dot_product_and_ReLU[13].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$1608(.Z({ \dot_product_and_ReLU[13].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$1609(.Z({ \dot_product_and_ReLU[13].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$1610(.Z({ \dot_product_and_ReLU[13].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$1611(.Z({ \dot_product_and_ReLU[13].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$1612(.Z({ \dot_product_and_ReLU[13].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$1613(.Z({ \dot_product_and_ReLU[13].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$1614(.Z({ \dot_product_and_ReLU[13].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$1615(.Z({ \dot_product_and_ReLU[13].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$1616(.Z({ \dot_product_and_ReLU[13].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$1617(.Z({ \dot_product_and_ReLU[13].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$1618(.Z({ \dot_product_and_ReLU[13].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$1619(.Z({ \dot_product_and_ReLU[13].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$1620(.Z({ \dot_product_and_ReLU[13].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$1621(.Z({ \dot_product_and_ReLU[13].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$1622(.Z({ \dot_product_and_ReLU[13].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$1623(.Z({ \dot_product_and_ReLU[13].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$1624(.Z({ \dot_product_and_ReLU[13].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$1625(.Z({ \dot_product_and_ReLU[13].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$1626(.Z({ \dot_product_and_ReLU[13].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$1627(.Z({ \dot_product_and_ReLU[13].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$1628(.Z({ \dot_product_and_ReLU[13].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$1629(.Z({ \dot_product_and_ReLU[13].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$1630(.Z({ \dot_product_and_ReLU[13].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$1631(.Z({ \dot_product_and_ReLU[13].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$1632(.Z({ \dot_product_and_ReLU[13].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$1633(.Z({ \dot_product_and_ReLU[13].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$1634(.Z({ \dot_product_and_ReLU[13].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$1635(.Z({ \dot_product_and_ReLU[13].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$1636(.Z({ \dot_product_and_ReLU[13].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$1637(.Z({ \dot_product_and_ReLU[13].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$1638(.Z({ \dot_product_and_ReLU[13].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$1639(.Z({ \dot_product_and_ReLU[13].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$1640(.Z({ \dot_product_and_ReLU[13].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$1641(.Z({ \dot_product_and_ReLU[13].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$1642(.Z({ \dot_product_and_ReLU[13].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$1643(.Z({ \dot_product_and_ReLU[13].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$1644(.Z({ \dot_product_and_ReLU[13].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$1645(.Z({ \dot_product_and_ReLU[13].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$1646(.Z({ \dot_product_and_ReLU[13].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$1647(.Z({ \dot_product_and_ReLU[13].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$1648(.Z({ \dot_product_and_ReLU[13].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$1649(.Z({ \dot_product_and_ReLU[13].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$1650(.Z({ \dot_product_and_ReLU[13].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$1651(.Z({ \dot_product_and_ReLU[13].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$1652(.Z({ \dot_product_and_ReLU[13].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$1653(.Z({ \dot_product_and_ReLU[13].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$1654(.Z({ \dot_product_and_ReLU[13].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$1655(.Z({ \dot_product_and_ReLU[13].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$1656(.Z({ \dot_product_and_ReLU[13].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$1657(.Z({ \dot_product_and_ReLU[13].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$1658(.Z({ \dot_product_and_ReLU[13].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$1659(.Z({ \dot_product_and_ReLU[13].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$1660(.Z({ \dot_product_and_ReLU[13].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$1661(.Z({ \dot_product_and_ReLU[13].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$1662(.Z({ \dot_product_and_ReLU[13].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$1663(.Z({ \dot_product_and_ReLU[13].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$1664(.Z({ \dot_product_and_ReLU[13].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$1665(.Z({ \dot_product_and_ReLU[13].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$1666(.Z({ \dot_product_and_ReLU[13].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$1667(.Z({ \dot_product_and_ReLU[13].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$1668(.Z({ \dot_product_and_ReLU[13].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$1669(.Z({ \dot_product_and_ReLU[13].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$1670(.Z({ \dot_product_and_ReLU[13].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$1671(.Z({ \dot_product_and_ReLU[13].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$1672(.Z({ \dot_product_and_ReLU[13].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$1673(.Z({ \dot_product_and_ReLU[13].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$1674(.Z({ \dot_product_and_ReLU[13].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$1675(.Z({ \dot_product_and_ReLU[13].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$1676(.Z({ \dot_product_and_ReLU[13].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$1677(.Z({ \dot_product_and_ReLU[13].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$1678(.Z({ \dot_product_and_ReLU[13].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$1679(.Z({ \dot_product_and_ReLU[13].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$1680(.Z({ \dot_product_and_ReLU[13].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$1681(.Z({ \dot_product_and_ReLU[13].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$1682(.Z({ \dot_product_and_ReLU[13].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$1683(.Z({ \dot_product_and_ReLU[13].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$1684(.Z({ \dot_product_and_ReLU[13].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$1685(.Z({ \dot_product_and_ReLU[13].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$1686(.Z({ \dot_product_and_ReLU[13].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$1687(.Z({ \dot_product_and_ReLU[13].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$1688(.Z({ \dot_product_and_ReLU[13].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$1689(.Z({ \dot_product_and_ReLU[13].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$1690(.Z({ \dot_product_and_ReLU[13].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$1691(.Z({ \dot_product_and_ReLU[13].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$1692(.Z({ \dot_product_and_ReLU[13].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$1693(.Z({ \dot_product_and_ReLU[13].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$1694(.Z({ \dot_product_and_ReLU[13].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$1695(.Z({ \dot_product_and_ReLU[13].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$1696(.Z({ \dot_product_and_ReLU[13].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$1697(.Z({ \dot_product_and_ReLU[13].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$1698(.Z({ \dot_product_and_ReLU[13].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$1699(.Z({ \dot_product_and_ReLU[13].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$1700(.Z({ \dot_product_and_ReLU[13].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$1701(.Z({ \dot_product_and_ReLU[13].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$1702(.Z({ \dot_product_and_ReLU[13].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$1703(.Z({ \dot_product_and_ReLU[13].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$1704(.Z({ \dot_product_and_ReLU[13].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$1705(.Z({ \dot_product_and_ReLU[13].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$1706(.Z({ \dot_product_and_ReLU[13].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$1707(.Z({ \dot_product_and_ReLU[13].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$1708(.Z({ \dot_product_and_ReLU[13].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$1709(.Z({ \dot_product_and_ReLU[13].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$1710(.Z({ \dot_product_and_ReLU[13].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$1711(.Z({ \dot_product_and_ReLU[13].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$1712(.Z({ \dot_product_and_ReLU[13].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$1713(.Z({ \dot_product_and_ReLU[13].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$1714(.Z({ \dot_product_and_ReLU[13].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$1715(.Z({ \dot_product_and_ReLU[13].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$1716(.Z({ \dot_product_and_ReLU[13].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$1717(.Z({ \dot_product_and_ReLU[13].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$1718(.Z({ \dot_product_and_ReLU[13].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$1719(.Z({ \dot_product_and_ReLU[13].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$1720(.Z({ \dot_product_and_ReLU[13].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$1721(.Z({ \dot_product_and_ReLU[13].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$1722(.Z({ \dot_product_and_ReLU[13].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$1723(.Z({ \dot_product_and_ReLU[13].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$1724(.Z({ \dot_product_and_ReLU[13].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$1725(.Z({ \dot_product_and_ReLU[13].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$1726(.Z({ \dot_product_and_ReLU[13].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$1727(.Z({ \dot_product_and_ReLU[13].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$1728(.Z({ \dot_product_and_ReLU[13].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$1729(.Z({ \dot_product_and_ReLU[13].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$1730(.Z({ \dot_product_and_ReLU[13].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$1731(.Z({ \dot_product_and_ReLU[13].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$1732(.Z({ \dot_product_and_ReLU[13].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$1733(.Z({ \dot_product_and_ReLU[13].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$1734(.Z({ \dot_product_and_ReLU[13].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$1735(.Z({ \dot_product_and_ReLU[13].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$1736(.Z({ \dot_product_and_ReLU[13].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$1737(.Z({ \dot_product_and_ReLU[13].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$1738(.Z({ \dot_product_and_ReLU[13].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$1739(.Z({ \dot_product_and_ReLU[13].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$1740(.Z({ \dot_product_and_ReLU[13].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$1741(.Z({ \dot_product_and_ReLU[13].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$1742(.Z({ \dot_product_and_ReLU[13].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$1743(.Z({ \dot_product_and_ReLU[13].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$1744(.Z({ \dot_product_and_ReLU[13].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$1745(.Z({ \dot_product_and_ReLU[13].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$1746(.Z({ \dot_product_and_ReLU[13].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$1747(.Z({ \dot_product_and_ReLU[13].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$1748(.Z({ \dot_product_and_ReLU[13].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$1749(.Z({ \dot_product_and_ReLU[13].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$1750(.Z({ \dot_product_and_ReLU[13].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$1751(.Z({ \dot_product_and_ReLU[13].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$1752(.Z({ \dot_product_and_ReLU[13].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$1753(.Z({ \dot_product_and_ReLU[13].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$1754(.Z({ \dot_product_and_ReLU[13].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$1755(.Z({ \dot_product_and_ReLU[13].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$1756(.Z({ \dot_product_and_ReLU[13].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$1757(.Z({ \dot_product_and_ReLU[13].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$1758(.Z({ \dot_product_and_ReLU[13].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$1759(.Z({ \dot_product_and_ReLU[13].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$1760(.Z({ \dot_product_and_ReLU[13].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$1761(.Z({ \dot_product_and_ReLU[13].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$1762(.Z({ \dot_product_and_ReLU[13].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$1763(.Z({ \dot_product_and_ReLU[13].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$1764(.Z({ \dot_product_and_ReLU[13].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$1765(.Z({ \dot_product_and_ReLU[13].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$1766(.Z({ \dot_product_and_ReLU[13].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$1767(.Z({ \dot_product_and_ReLU[13].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$1768(.Z({ \dot_product_and_ReLU[13].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$1769(.Z({ \dot_product_and_ReLU[13].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$1770(.Z({ \dot_product_and_ReLU[13].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$1771(.Z({ \dot_product_and_ReLU[13].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$1772(.Z({ \dot_product_and_ReLU[13].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$1773(.Z({ \dot_product_and_ReLU[13].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$1774(.Z({ \dot_product_and_ReLU[13].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$1775(.Z({ \dot_product_and_ReLU[13].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$1776(.Z({ \dot_product_and_ReLU[13].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$1777(.Z({ \dot_product_and_ReLU[13].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$1778(.Z({ \dot_product_and_ReLU[13].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$1779(.Z({ \dot_product_and_ReLU[13].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$1780(.Z({ \dot_product_and_ReLU[13].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$1781(.Z({ \dot_product_and_ReLU[13].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$1782(.Z({ \dot_product_and_ReLU[13].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$1783(.Z({ \dot_product_and_ReLU[13].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$1784(.Z({ \dot_product_and_ReLU[13].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$1785(.Z({ \dot_product_and_ReLU[13].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$1786(.Z({ \dot_product_and_ReLU[13].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$1787(.Z({ \dot_product_and_ReLU[13].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$1788(.Z({ \dot_product_and_ReLU[13].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$1789(.Z({ \dot_product_and_ReLU[13].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$1790(.Z({ \dot_product_and_ReLU[13].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$1791(.Z({ \dot_product_and_ReLU[13].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$1792(.Z({ \dot_product_and_ReLU[13].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[13][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$1793(.Z({ \dot_product_and_ReLU[12].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$1794(.Z({ \dot_product_and_ReLU[12].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$1795(.Z({ \dot_product_and_ReLU[12].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$1796(.Z({ \dot_product_and_ReLU[12].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$1797(.Z({ \dot_product_and_ReLU[12].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$1798(.Z({ \dot_product_and_ReLU[12].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$1799(.Z({ \dot_product_and_ReLU[12].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$1800(.Z({ \dot_product_and_ReLU[12].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$1801(.Z({ \dot_product_and_ReLU[12].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$1802(.Z({ \dot_product_and_ReLU[12].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$1803(.Z({ \dot_product_and_ReLU[12].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$1804(.Z({ \dot_product_and_ReLU[12].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$1805(.Z({ \dot_product_and_ReLU[12].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$1806(.Z({ \dot_product_and_ReLU[12].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$1807(.Z({ \dot_product_and_ReLU[12].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$1808(.Z({ \dot_product_and_ReLU[12].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$1809(.Z({ \dot_product_and_ReLU[12].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$1810(.Z({ \dot_product_and_ReLU[12].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$1811(.Z({ \dot_product_and_ReLU[12].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$1812(.Z({ \dot_product_and_ReLU[12].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$1813(.Z({ \dot_product_and_ReLU[12].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$1814(.Z({ \dot_product_and_ReLU[12].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$1815(.Z({ \dot_product_and_ReLU[12].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$1816(.Z({ \dot_product_and_ReLU[12].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$1817(.Z({ \dot_product_and_ReLU[12].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$1818(.Z({ \dot_product_and_ReLU[12].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$1819(.Z({ \dot_product_and_ReLU[12].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$1820(.Z({ \dot_product_and_ReLU[12].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$1821(.Z({ \dot_product_and_ReLU[12].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$1822(.Z({ \dot_product_and_ReLU[12].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$1823(.Z({ \dot_product_and_ReLU[12].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$1824(.Z({ \dot_product_and_ReLU[12].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$1825(.Z({ \dot_product_and_ReLU[12].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$1826(.Z({ \dot_product_and_ReLU[12].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$1827(.Z({ \dot_product_and_ReLU[12].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$1828(.Z({ \dot_product_and_ReLU[12].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$1829(.Z({ \dot_product_and_ReLU[12].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$1830(.Z({ \dot_product_and_ReLU[12].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$1831(.Z({ \dot_product_and_ReLU[12].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$1832(.Z({ \dot_product_and_ReLU[12].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$1833(.Z({ \dot_product_and_ReLU[12].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$1834(.Z({ \dot_product_and_ReLU[12].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$1835(.Z({ \dot_product_and_ReLU[12].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$1836(.Z({ \dot_product_and_ReLU[12].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$1837(.Z({ \dot_product_and_ReLU[12].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$1838(.Z({ \dot_product_and_ReLU[12].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$1839(.Z({ \dot_product_and_ReLU[12].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$1840(.Z({ \dot_product_and_ReLU[12].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$1841(.Z({ \dot_product_and_ReLU[12].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$1842(.Z({ \dot_product_and_ReLU[12].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$1843(.Z({ \dot_product_and_ReLU[12].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$1844(.Z({ \dot_product_and_ReLU[12].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$1845(.Z({ \dot_product_and_ReLU[12].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$1846(.Z({ \dot_product_and_ReLU[12].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$1847(.Z({ \dot_product_and_ReLU[12].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$1848(.Z({ \dot_product_and_ReLU[12].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$1849(.Z({ \dot_product_and_ReLU[12].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$1850(.Z({ \dot_product_and_ReLU[12].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$1851(.Z({ \dot_product_and_ReLU[12].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$1852(.Z({ \dot_product_and_ReLU[12].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$1853(.Z({ \dot_product_and_ReLU[12].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$1854(.Z({ \dot_product_and_ReLU[12].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$1855(.Z({ \dot_product_and_ReLU[12].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$1856(.Z({ \dot_product_and_ReLU[12].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$1857(.Z({ \dot_product_and_ReLU[12].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$1858(.Z({ \dot_product_and_ReLU[12].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$1859(.Z({ \dot_product_and_ReLU[12].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$1860(.Z({ \dot_product_and_ReLU[12].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$1861(.Z({ \dot_product_and_ReLU[12].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$1862(.Z({ \dot_product_and_ReLU[12].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$1863(.Z({ \dot_product_and_ReLU[12].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$1864(.Z({ \dot_product_and_ReLU[12].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$1865(.Z({ \dot_product_and_ReLU[12].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$1866(.Z({ \dot_product_and_ReLU[12].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$1867(.Z({ \dot_product_and_ReLU[12].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$1868(.Z({ \dot_product_and_ReLU[12].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$1869(.Z({ \dot_product_and_ReLU[12].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$1870(.Z({ \dot_product_and_ReLU[12].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$1871(.Z({ \dot_product_and_ReLU[12].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$1872(.Z({ \dot_product_and_ReLU[12].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$1873(.Z({ \dot_product_and_ReLU[12].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$1874(.Z({ \dot_product_and_ReLU[12].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$1875(.Z({ \dot_product_and_ReLU[12].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$1876(.Z({ \dot_product_and_ReLU[12].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$1877(.Z({ \dot_product_and_ReLU[12].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$1878(.Z({ \dot_product_and_ReLU[12].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$1879(.Z({ \dot_product_and_ReLU[12].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$1880(.Z({ \dot_product_and_ReLU[12].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$1881(.Z({ \dot_product_and_ReLU[12].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$1882(.Z({ \dot_product_and_ReLU[12].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$1883(.Z({ \dot_product_and_ReLU[12].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$1884(.Z({ \dot_product_and_ReLU[12].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$1885(.Z({ \dot_product_and_ReLU[12].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$1886(.Z({ \dot_product_and_ReLU[12].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$1887(.Z({ \dot_product_and_ReLU[12].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$1888(.Z({ \dot_product_and_ReLU[12].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$1889(.Z({ \dot_product_and_ReLU[12].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$1890(.Z({ \dot_product_and_ReLU[12].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$1891(.Z({ \dot_product_and_ReLU[12].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$1892(.Z({ \dot_product_and_ReLU[12].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$1893(.Z({ \dot_product_and_ReLU[12].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$1894(.Z({ \dot_product_and_ReLU[12].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$1895(.Z({ \dot_product_and_ReLU[12].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$1896(.Z({ \dot_product_and_ReLU[12].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$1897(.Z({ \dot_product_and_ReLU[12].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$1898(.Z({ \dot_product_and_ReLU[12].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$1899(.Z({ \dot_product_and_ReLU[12].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$1900(.Z({ \dot_product_and_ReLU[12].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$1901(.Z({ \dot_product_and_ReLU[12].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$1902(.Z({ \dot_product_and_ReLU[12].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$1903(.Z({ \dot_product_and_ReLU[12].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$1904(.Z({ \dot_product_and_ReLU[12].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$1905(.Z({ \dot_product_and_ReLU[12].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$1906(.Z({ \dot_product_and_ReLU[12].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$1907(.Z({ \dot_product_and_ReLU[12].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$1908(.Z({ \dot_product_and_ReLU[12].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$1909(.Z({ \dot_product_and_ReLU[12].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$1910(.Z({ \dot_product_and_ReLU[12].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$1911(.Z({ \dot_product_and_ReLU[12].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$1912(.Z({ \dot_product_and_ReLU[12].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$1913(.Z({ \dot_product_and_ReLU[12].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$1914(.Z({ \dot_product_and_ReLU[12].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$1915(.Z({ \dot_product_and_ReLU[12].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$1916(.Z({ \dot_product_and_ReLU[12].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$1917(.Z({ \dot_product_and_ReLU[12].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$1918(.Z({ \dot_product_and_ReLU[12].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$1919(.Z({ \dot_product_and_ReLU[12].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$1920(.Z({ \dot_product_and_ReLU[12].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$1921(.Z({ \dot_product_and_ReLU[12].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$1922(.Z({ \dot_product_and_ReLU[12].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$1923(.Z({ \dot_product_and_ReLU[12].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$1924(.Z({ \dot_product_and_ReLU[12].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$1925(.Z({ \dot_product_and_ReLU[12].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$1926(.Z({ \dot_product_and_ReLU[12].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$1927(.Z({ \dot_product_and_ReLU[12].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$1928(.Z({ \dot_product_and_ReLU[12].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$1929(.Z({ \dot_product_and_ReLU[12].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$1930(.Z({ \dot_product_and_ReLU[12].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$1931(.Z({ \dot_product_and_ReLU[12].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$1932(.Z({ \dot_product_and_ReLU[12].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$1933(.Z({ \dot_product_and_ReLU[12].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$1934(.Z({ \dot_product_and_ReLU[12].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$1935(.Z({ \dot_product_and_ReLU[12].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$1936(.Z({ \dot_product_and_ReLU[12].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$1937(.Z({ \dot_product_and_ReLU[12].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$1938(.Z({ \dot_product_and_ReLU[12].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$1939(.Z({ \dot_product_and_ReLU[12].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$1940(.Z({ \dot_product_and_ReLU[12].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$1941(.Z({ \dot_product_and_ReLU[12].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$1942(.Z({ \dot_product_and_ReLU[12].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$1943(.Z({ \dot_product_and_ReLU[12].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$1944(.Z({ \dot_product_and_ReLU[12].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$1945(.Z({ \dot_product_and_ReLU[12].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$1946(.Z({ \dot_product_and_ReLU[12].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$1947(.Z({ \dot_product_and_ReLU[12].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$1948(.Z({ \dot_product_and_ReLU[12].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$1949(.Z({ \dot_product_and_ReLU[12].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$1950(.Z({ \dot_product_and_ReLU[12].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$1951(.Z({ \dot_product_and_ReLU[12].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$1952(.Z({ \dot_product_and_ReLU[12].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$1953(.Z({ \dot_product_and_ReLU[12].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$1954(.Z({ \dot_product_and_ReLU[12].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$1955(.Z({ \dot_product_and_ReLU[12].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$1956(.Z({ \dot_product_and_ReLU[12].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$1957(.Z({ \dot_product_and_ReLU[12].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$1958(.Z({ \dot_product_and_ReLU[12].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$1959(.Z({ \dot_product_and_ReLU[12].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$1960(.Z({ \dot_product_and_ReLU[12].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$1961(.Z({ \dot_product_and_ReLU[12].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$1962(.Z({ \dot_product_and_ReLU[12].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$1963(.Z({ \dot_product_and_ReLU[12].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$1964(.Z({ \dot_product_and_ReLU[12].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$1965(.Z({ \dot_product_and_ReLU[12].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$1966(.Z({ \dot_product_and_ReLU[12].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$1967(.Z({ \dot_product_and_ReLU[12].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$1968(.Z({ \dot_product_and_ReLU[12].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$1969(.Z({ \dot_product_and_ReLU[12].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$1970(.Z({ \dot_product_and_ReLU[12].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$1971(.Z({ \dot_product_and_ReLU[12].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$1972(.Z({ \dot_product_and_ReLU[12].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$1973(.Z({ \dot_product_and_ReLU[12].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$1974(.Z({ \dot_product_and_ReLU[12].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$1975(.Z({ \dot_product_and_ReLU[12].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$1976(.Z({ \dot_product_and_ReLU[12].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$1977(.Z({ \dot_product_and_ReLU[12].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$1978(.Z({ \dot_product_and_ReLU[12].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$1979(.Z({ \dot_product_and_ReLU[12].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$1980(.Z({ \dot_product_and_ReLU[12].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$1981(.Z({ \dot_product_and_ReLU[12].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$1982(.Z({ \dot_product_and_ReLU[12].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$1983(.Z({ \dot_product_and_ReLU[12].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$1984(.Z({ \dot_product_and_ReLU[12].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$1985(.Z({ \dot_product_and_ReLU[12].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$1986(.Z({ \dot_product_and_ReLU[12].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$1987(.Z({ \dot_product_and_ReLU[12].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$1988(.Z({ \dot_product_and_ReLU[12].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$1989(.Z({ \dot_product_and_ReLU[12].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$1990(.Z({ \dot_product_and_ReLU[12].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$1991(.Z({ \dot_product_and_ReLU[12].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$1992(.Z({ \dot_product_and_ReLU[12].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$1993(.Z({ \dot_product_and_ReLU[12].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$1994(.Z({ \dot_product_and_ReLU[12].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$1995(.Z({ \dot_product_and_ReLU[12].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$1996(.Z({ \dot_product_and_ReLU[12].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$1997(.Z({ \dot_product_and_ReLU[12].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$1998(.Z({ \dot_product_and_ReLU[12].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$1999(.Z({ \dot_product_and_ReLU[12].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$2000(.Z({ \dot_product_and_ReLU[12].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$2001(.Z({ \dot_product_and_ReLU[12].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$2002(.Z({ \dot_product_and_ReLU[12].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$2003(.Z({ \dot_product_and_ReLU[12].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$2004(.Z({ \dot_product_and_ReLU[12].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$2005(.Z({ \dot_product_and_ReLU[12].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$2006(.Z({ \dot_product_and_ReLU[12].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$2007(.Z({ \dot_product_and_ReLU[12].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$2008(.Z({ \dot_product_and_ReLU[12].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$2009(.Z({ \dot_product_and_ReLU[12].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$2010(.Z({ \dot_product_and_ReLU[12].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$2011(.Z({ \dot_product_and_ReLU[12].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$2012(.Z({ \dot_product_and_ReLU[12].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$2013(.Z({ \dot_product_and_ReLU[12].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$2014(.Z({ \dot_product_and_ReLU[12].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$2015(.Z({ \dot_product_and_ReLU[12].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$2016(.Z({ \dot_product_and_ReLU[12].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$2017(.Z({ \dot_product_and_ReLU[12].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$2018(.Z({ \dot_product_and_ReLU[12].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$2019(.Z({ \dot_product_and_ReLU[12].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$2020(.Z({ \dot_product_and_ReLU[12].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$2021(.Z({ \dot_product_and_ReLU[12].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$2022(.Z({ \dot_product_and_ReLU[12].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$2023(.Z({ \dot_product_and_ReLU[12].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$2024(.Z({ \dot_product_and_ReLU[12].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$2025(.Z({ \dot_product_and_ReLU[12].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$2026(.Z({ \dot_product_and_ReLU[12].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$2027(.Z({ \dot_product_and_ReLU[12].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$2028(.Z({ \dot_product_and_ReLU[12].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$2029(.Z({ \dot_product_and_ReLU[12].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$2030(.Z({ \dot_product_and_ReLU[12].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$2031(.Z({ \dot_product_and_ReLU[12].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$2032(.Z({ \dot_product_and_ReLU[12].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$2033(.Z({ \dot_product_and_ReLU[12].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$2034(.Z({ \dot_product_and_ReLU[12].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$2035(.Z({ \dot_product_and_ReLU[12].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$2036(.Z({ \dot_product_and_ReLU[12].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$2037(.Z({ \dot_product_and_ReLU[12].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$2038(.Z({ \dot_product_and_ReLU[12].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$2039(.Z({ \dot_product_and_ReLU[12].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$2040(.Z({ \dot_product_and_ReLU[12].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$2041(.Z({ \dot_product_and_ReLU[12].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$2042(.Z({ \dot_product_and_ReLU[12].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$2043(.Z({ \dot_product_and_ReLU[12].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$2044(.Z({ \dot_product_and_ReLU[12].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$2045(.Z({ \dot_product_and_ReLU[12].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$2046(.Z({ \dot_product_and_ReLU[12].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$2047(.Z({ \dot_product_and_ReLU[12].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$2048(.Z({ \dot_product_and_ReLU[12].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[12][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$2049(.Z({ \dot_product_and_ReLU[11].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$2050(.Z({ \dot_product_and_ReLU[11].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$2051(.Z({ \dot_product_and_ReLU[11].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$2052(.Z({ \dot_product_and_ReLU[11].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$2053(.Z({ \dot_product_and_ReLU[11].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$2054(.Z({ \dot_product_and_ReLU[11].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$2055(.Z({ \dot_product_and_ReLU[11].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$2056(.Z({ \dot_product_and_ReLU[11].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$2057(.Z({ \dot_product_and_ReLU[11].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$2058(.Z({ \dot_product_and_ReLU[11].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$2059(.Z({ \dot_product_and_ReLU[11].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$2060(.Z({ \dot_product_and_ReLU[11].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$2061(.Z({ \dot_product_and_ReLU[11].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$2062(.Z({ \dot_product_and_ReLU[11].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$2063(.Z({ \dot_product_and_ReLU[11].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$2064(.Z({ \dot_product_and_ReLU[11].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$2065(.Z({ \dot_product_and_ReLU[11].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$2066(.Z({ \dot_product_and_ReLU[11].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$2067(.Z({ \dot_product_and_ReLU[11].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$2068(.Z({ \dot_product_and_ReLU[11].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$2069(.Z({ \dot_product_and_ReLU[11].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$2070(.Z({ \dot_product_and_ReLU[11].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$2071(.Z({ \dot_product_and_ReLU[11].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$2072(.Z({ \dot_product_and_ReLU[11].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$2073(.Z({ \dot_product_and_ReLU[11].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$2074(.Z({ \dot_product_and_ReLU[11].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$2075(.Z({ \dot_product_and_ReLU[11].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$2076(.Z({ \dot_product_and_ReLU[11].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$2077(.Z({ \dot_product_and_ReLU[11].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$2078(.Z({ \dot_product_and_ReLU[11].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$2079(.Z({ \dot_product_and_ReLU[11].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$2080(.Z({ \dot_product_and_ReLU[11].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$2081(.Z({ \dot_product_and_ReLU[11].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$2082(.Z({ \dot_product_and_ReLU[11].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$2083(.Z({ \dot_product_and_ReLU[11].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$2084(.Z({ \dot_product_and_ReLU[11].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$2085(.Z({ \dot_product_and_ReLU[11].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$2086(.Z({ \dot_product_and_ReLU[11].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$2087(.Z({ \dot_product_and_ReLU[11].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$2088(.Z({ \dot_product_and_ReLU[11].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$2089(.Z({ \dot_product_and_ReLU[11].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$2090(.Z({ \dot_product_and_ReLU[11].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$2091(.Z({ \dot_product_and_ReLU[11].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$2092(.Z({ \dot_product_and_ReLU[11].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$2093(.Z({ \dot_product_and_ReLU[11].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$2094(.Z({ \dot_product_and_ReLU[11].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$2095(.Z({ \dot_product_and_ReLU[11].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$2096(.Z({ \dot_product_and_ReLU[11].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$2097(.Z({ \dot_product_and_ReLU[11].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$2098(.Z({ \dot_product_and_ReLU[11].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$2099(.Z({ \dot_product_and_ReLU[11].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$2100(.Z({ \dot_product_and_ReLU[11].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$2101(.Z({ \dot_product_and_ReLU[11].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$2102(.Z({ \dot_product_and_ReLU[11].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$2103(.Z({ \dot_product_and_ReLU[11].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$2104(.Z({ \dot_product_and_ReLU[11].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$2105(.Z({ \dot_product_and_ReLU[11].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$2106(.Z({ \dot_product_and_ReLU[11].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$2107(.Z({ \dot_product_and_ReLU[11].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$2108(.Z({ \dot_product_and_ReLU[11].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$2109(.Z({ \dot_product_and_ReLU[11].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$2110(.Z({ \dot_product_and_ReLU[11].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$2111(.Z({ \dot_product_and_ReLU[11].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$2112(.Z({ \dot_product_and_ReLU[11].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$2113(.Z({ \dot_product_and_ReLU[11].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$2114(.Z({ \dot_product_and_ReLU[11].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$2115(.Z({ \dot_product_and_ReLU[11].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$2116(.Z({ \dot_product_and_ReLU[11].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$2117(.Z({ \dot_product_and_ReLU[11].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$2118(.Z({ \dot_product_and_ReLU[11].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$2119(.Z({ \dot_product_and_ReLU[11].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$2120(.Z({ \dot_product_and_ReLU[11].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$2121(.Z({ \dot_product_and_ReLU[11].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$2122(.Z({ \dot_product_and_ReLU[11].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$2123(.Z({ \dot_product_and_ReLU[11].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$2124(.Z({ \dot_product_and_ReLU[11].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$2125(.Z({ \dot_product_and_ReLU[11].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$2126(.Z({ \dot_product_and_ReLU[11].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$2127(.Z({ \dot_product_and_ReLU[11].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$2128(.Z({ \dot_product_and_ReLU[11].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$2129(.Z({ \dot_product_and_ReLU[11].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$2130(.Z({ \dot_product_and_ReLU[11].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$2131(.Z({ \dot_product_and_ReLU[11].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$2132(.Z({ \dot_product_and_ReLU[11].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$2133(.Z({ \dot_product_and_ReLU[11].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$2134(.Z({ \dot_product_and_ReLU[11].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$2135(.Z({ \dot_product_and_ReLU[11].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$2136(.Z({ \dot_product_and_ReLU[11].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$2137(.Z({ \dot_product_and_ReLU[11].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$2138(.Z({ \dot_product_and_ReLU[11].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$2139(.Z({ \dot_product_and_ReLU[11].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$2140(.Z({ \dot_product_and_ReLU[11].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$2141(.Z({ \dot_product_and_ReLU[11].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$2142(.Z({ \dot_product_and_ReLU[11].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$2143(.Z({ \dot_product_and_ReLU[11].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$2144(.Z({ \dot_product_and_ReLU[11].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$2145(.Z({ \dot_product_and_ReLU[11].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$2146(.Z({ \dot_product_and_ReLU[11].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$2147(.Z({ \dot_product_and_ReLU[11].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$2148(.Z({ \dot_product_and_ReLU[11].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$2149(.Z({ \dot_product_and_ReLU[11].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$2150(.Z({ \dot_product_and_ReLU[11].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$2151(.Z({ \dot_product_and_ReLU[11].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$2152(.Z({ \dot_product_and_ReLU[11].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$2153(.Z({ \dot_product_and_ReLU[11].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$2154(.Z({ \dot_product_and_ReLU[11].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$2155(.Z({ \dot_product_and_ReLU[11].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$2156(.Z({ \dot_product_and_ReLU[11].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$2157(.Z({ \dot_product_and_ReLU[11].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$2158(.Z({ \dot_product_and_ReLU[11].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$2159(.Z({ \dot_product_and_ReLU[11].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$2160(.Z({ \dot_product_and_ReLU[11].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$2161(.Z({ \dot_product_and_ReLU[11].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$2162(.Z({ \dot_product_and_ReLU[11].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$2163(.Z({ \dot_product_and_ReLU[11].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$2164(.Z({ \dot_product_and_ReLU[11].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$2165(.Z({ \dot_product_and_ReLU[11].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$2166(.Z({ \dot_product_and_ReLU[11].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$2167(.Z({ \dot_product_and_ReLU[11].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$2168(.Z({ \dot_product_and_ReLU[11].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$2169(.Z({ \dot_product_and_ReLU[11].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$2170(.Z({ \dot_product_and_ReLU[11].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$2171(.Z({ \dot_product_and_ReLU[11].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$2172(.Z({ \dot_product_and_ReLU[11].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$2173(.Z({ \dot_product_and_ReLU[11].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$2174(.Z({ \dot_product_and_ReLU[11].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$2175(.Z({ \dot_product_and_ReLU[11].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$2176(.Z({ \dot_product_and_ReLU[11].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$2177(.Z({ \dot_product_and_ReLU[11].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$2178(.Z({ \dot_product_and_ReLU[11].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$2179(.Z({ \dot_product_and_ReLU[11].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$2180(.Z({ \dot_product_and_ReLU[11].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$2181(.Z({ \dot_product_and_ReLU[11].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$2182(.Z({ \dot_product_and_ReLU[11].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$2183(.Z({ \dot_product_and_ReLU[11].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$2184(.Z({ \dot_product_and_ReLU[11].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$2185(.Z({ \dot_product_and_ReLU[11].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$2186(.Z({ \dot_product_and_ReLU[11].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$2187(.Z({ \dot_product_and_ReLU[11].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$2188(.Z({ \dot_product_and_ReLU[11].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$2189(.Z({ \dot_product_and_ReLU[11].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$2190(.Z({ \dot_product_and_ReLU[11].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$2191(.Z({ \dot_product_and_ReLU[11].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$2192(.Z({ \dot_product_and_ReLU[11].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$2193(.Z({ \dot_product_and_ReLU[11].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$2194(.Z({ \dot_product_and_ReLU[11].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$2195(.Z({ \dot_product_and_ReLU[11].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$2196(.Z({ \dot_product_and_ReLU[11].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$2197(.Z({ \dot_product_and_ReLU[11].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$2198(.Z({ \dot_product_and_ReLU[11].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$2199(.Z({ \dot_product_and_ReLU[11].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$2200(.Z({ \dot_product_and_ReLU[11].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$2201(.Z({ \dot_product_and_ReLU[11].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$2202(.Z({ \dot_product_and_ReLU[11].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$2203(.Z({ \dot_product_and_ReLU[11].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$2204(.Z({ \dot_product_and_ReLU[11].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$2205(.Z({ \dot_product_and_ReLU[11].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$2206(.Z({ \dot_product_and_ReLU[11].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$2207(.Z({ \dot_product_and_ReLU[11].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$2208(.Z({ \dot_product_and_ReLU[11].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$2209(.Z({ \dot_product_and_ReLU[11].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$2210(.Z({ \dot_product_and_ReLU[11].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$2211(.Z({ \dot_product_and_ReLU[11].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$2212(.Z({ \dot_product_and_ReLU[11].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$2213(.Z({ \dot_product_and_ReLU[11].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$2214(.Z({ \dot_product_and_ReLU[11].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$2215(.Z({ \dot_product_and_ReLU[11].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$2216(.Z({ \dot_product_and_ReLU[11].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$2217(.Z({ \dot_product_and_ReLU[11].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$2218(.Z({ \dot_product_and_ReLU[11].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$2219(.Z({ \dot_product_and_ReLU[11].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$2220(.Z({ \dot_product_and_ReLU[11].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$2221(.Z({ \dot_product_and_ReLU[11].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$2222(.Z({ \dot_product_and_ReLU[11].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$2223(.Z({ \dot_product_and_ReLU[11].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$2224(.Z({ \dot_product_and_ReLU[11].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$2225(.Z({ \dot_product_and_ReLU[11].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$2226(.Z({ \dot_product_and_ReLU[11].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$2227(.Z({ \dot_product_and_ReLU[11].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$2228(.Z({ \dot_product_and_ReLU[11].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$2229(.Z({ \dot_product_and_ReLU[11].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$2230(.Z({ \dot_product_and_ReLU[11].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$2231(.Z({ \dot_product_and_ReLU[11].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$2232(.Z({ \dot_product_and_ReLU[11].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$2233(.Z({ \dot_product_and_ReLU[11].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$2234(.Z({ \dot_product_and_ReLU[11].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$2235(.Z({ \dot_product_and_ReLU[11].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$2236(.Z({ \dot_product_and_ReLU[11].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$2237(.Z({ \dot_product_and_ReLU[11].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$2238(.Z({ \dot_product_and_ReLU[11].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$2239(.Z({ \dot_product_and_ReLU[11].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$2240(.Z({ \dot_product_and_ReLU[11].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$2241(.Z({ \dot_product_and_ReLU[11].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$2242(.Z({ \dot_product_and_ReLU[11].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$2243(.Z({ \dot_product_and_ReLU[11].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$2244(.Z({ \dot_product_and_ReLU[11].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$2245(.Z({ \dot_product_and_ReLU[11].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$2246(.Z({ \dot_product_and_ReLU[11].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$2247(.Z({ \dot_product_and_ReLU[11].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$2248(.Z({ \dot_product_and_ReLU[11].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$2249(.Z({ \dot_product_and_ReLU[11].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$2250(.Z({ \dot_product_and_ReLU[11].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$2251(.Z({ \dot_product_and_ReLU[11].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$2252(.Z({ \dot_product_and_ReLU[11].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$2253(.Z({ \dot_product_and_ReLU[11].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$2254(.Z({ \dot_product_and_ReLU[11].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$2255(.Z({ \dot_product_and_ReLU[11].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$2256(.Z({ \dot_product_and_ReLU[11].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$2257(.Z({ \dot_product_and_ReLU[11].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$2258(.Z({ \dot_product_and_ReLU[11].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$2259(.Z({ \dot_product_and_ReLU[11].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$2260(.Z({ \dot_product_and_ReLU[11].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$2261(.Z({ \dot_product_and_ReLU[11].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$2262(.Z({ \dot_product_and_ReLU[11].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$2263(.Z({ \dot_product_and_ReLU[11].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$2264(.Z({ \dot_product_and_ReLU[11].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$2265(.Z({ \dot_product_and_ReLU[11].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$2266(.Z({ \dot_product_and_ReLU[11].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$2267(.Z({ \dot_product_and_ReLU[11].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$2268(.Z({ \dot_product_and_ReLU[11].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$2269(.Z({ \dot_product_and_ReLU[11].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$2270(.Z({ \dot_product_and_ReLU[11].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$2271(.Z({ \dot_product_and_ReLU[11].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$2272(.Z({ \dot_product_and_ReLU[11].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$2273(.Z({ \dot_product_and_ReLU[11].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$2274(.Z({ \dot_product_and_ReLU[11].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$2275(.Z({ \dot_product_and_ReLU[11].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$2276(.Z({ \dot_product_and_ReLU[11].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$2277(.Z({ \dot_product_and_ReLU[11].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$2278(.Z({ \dot_product_and_ReLU[11].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$2279(.Z({ \dot_product_and_ReLU[11].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$2280(.Z({ \dot_product_and_ReLU[11].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$2281(.Z({ \dot_product_and_ReLU[11].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$2282(.Z({ \dot_product_and_ReLU[11].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$2283(.Z({ \dot_product_and_ReLU[11].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$2284(.Z({ \dot_product_and_ReLU[11].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$2285(.Z({ \dot_product_and_ReLU[11].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$2286(.Z({ \dot_product_and_ReLU[11].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$2287(.Z({ \dot_product_and_ReLU[11].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$2288(.Z({ \dot_product_and_ReLU[11].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$2289(.Z({ \dot_product_and_ReLU[11].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$2290(.Z({ \dot_product_and_ReLU[11].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$2291(.Z({ \dot_product_and_ReLU[11].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$2292(.Z({ \dot_product_and_ReLU[11].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$2293(.Z({ \dot_product_and_ReLU[11].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$2294(.Z({ \dot_product_and_ReLU[11].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$2295(.Z({ \dot_product_and_ReLU[11].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$2296(.Z({ \dot_product_and_ReLU[11].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$2297(.Z({ \dot_product_and_ReLU[11].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$2298(.Z({ \dot_product_and_ReLU[11].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$2299(.Z({ \dot_product_and_ReLU[11].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$2300(.Z({ \dot_product_and_ReLU[11].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$2301(.Z({ \dot_product_and_ReLU[11].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$2302(.Z({ \dot_product_and_ReLU[11].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$2303(.Z({ \dot_product_and_ReLU[11].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$2304(.Z({ \dot_product_and_ReLU[11].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[11][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$2305(.Z({ \dot_product_and_ReLU[10].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$2306(.Z({ \dot_product_and_ReLU[10].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$2307(.Z({ \dot_product_and_ReLU[10].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$2308(.Z({ \dot_product_and_ReLU[10].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$2309(.Z({ \dot_product_and_ReLU[10].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$2310(.Z({ \dot_product_and_ReLU[10].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$2311(.Z({ \dot_product_and_ReLU[10].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$2312(.Z({ \dot_product_and_ReLU[10].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$2313(.Z({ \dot_product_and_ReLU[10].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$2314(.Z({ \dot_product_and_ReLU[10].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$2315(.Z({ \dot_product_and_ReLU[10].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$2316(.Z({ \dot_product_and_ReLU[10].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$2317(.Z({ \dot_product_and_ReLU[10].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$2318(.Z({ \dot_product_and_ReLU[10].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$2319(.Z({ \dot_product_and_ReLU[10].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$2320(.Z({ \dot_product_and_ReLU[10].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$2321(.Z({ \dot_product_and_ReLU[10].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$2322(.Z({ \dot_product_and_ReLU[10].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$2323(.Z({ \dot_product_and_ReLU[10].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$2324(.Z({ \dot_product_and_ReLU[10].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$2325(.Z({ \dot_product_and_ReLU[10].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$2326(.Z({ \dot_product_and_ReLU[10].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$2327(.Z({ \dot_product_and_ReLU[10].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$2328(.Z({ \dot_product_and_ReLU[10].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$2329(.Z({ \dot_product_and_ReLU[10].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$2330(.Z({ \dot_product_and_ReLU[10].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$2331(.Z({ \dot_product_and_ReLU[10].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$2332(.Z({ \dot_product_and_ReLU[10].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$2333(.Z({ \dot_product_and_ReLU[10].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$2334(.Z({ \dot_product_and_ReLU[10].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$2335(.Z({ \dot_product_and_ReLU[10].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$2336(.Z({ \dot_product_and_ReLU[10].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$2337(.Z({ \dot_product_and_ReLU[10].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$2338(.Z({ \dot_product_and_ReLU[10].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$2339(.Z({ \dot_product_and_ReLU[10].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$2340(.Z({ \dot_product_and_ReLU[10].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$2341(.Z({ \dot_product_and_ReLU[10].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$2342(.Z({ \dot_product_and_ReLU[10].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$2343(.Z({ \dot_product_and_ReLU[10].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$2344(.Z({ \dot_product_and_ReLU[10].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$2345(.Z({ \dot_product_and_ReLU[10].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$2346(.Z({ \dot_product_and_ReLU[10].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$2347(.Z({ \dot_product_and_ReLU[10].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$2348(.Z({ \dot_product_and_ReLU[10].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$2349(.Z({ \dot_product_and_ReLU[10].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$2350(.Z({ \dot_product_and_ReLU[10].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$2351(.Z({ \dot_product_and_ReLU[10].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$2352(.Z({ \dot_product_and_ReLU[10].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$2353(.Z({ \dot_product_and_ReLU[10].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$2354(.Z({ \dot_product_and_ReLU[10].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$2355(.Z({ \dot_product_and_ReLU[10].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$2356(.Z({ \dot_product_and_ReLU[10].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$2357(.Z({ \dot_product_and_ReLU[10].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$2358(.Z({ \dot_product_and_ReLU[10].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$2359(.Z({ \dot_product_and_ReLU[10].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$2360(.Z({ \dot_product_and_ReLU[10].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$2361(.Z({ \dot_product_and_ReLU[10].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$2362(.Z({ \dot_product_and_ReLU[10].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$2363(.Z({ \dot_product_and_ReLU[10].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$2364(.Z({ \dot_product_and_ReLU[10].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$2365(.Z({ \dot_product_and_ReLU[10].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$2366(.Z({ \dot_product_and_ReLU[10].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$2367(.Z({ \dot_product_and_ReLU[10].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$2368(.Z({ \dot_product_and_ReLU[10].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$2369(.Z({ \dot_product_and_ReLU[10].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$2370(.Z({ \dot_product_and_ReLU[10].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$2371(.Z({ \dot_product_and_ReLU[10].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$2372(.Z({ \dot_product_and_ReLU[10].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$2373(.Z({ \dot_product_and_ReLU[10].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$2374(.Z({ \dot_product_and_ReLU[10].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$2375(.Z({ \dot_product_and_ReLU[10].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$2376(.Z({ \dot_product_and_ReLU[10].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$2377(.Z({ \dot_product_and_ReLU[10].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$2378(.Z({ \dot_product_and_ReLU[10].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$2379(.Z({ \dot_product_and_ReLU[10].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$2380(.Z({ \dot_product_and_ReLU[10].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$2381(.Z({ \dot_product_and_ReLU[10].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$2382(.Z({ \dot_product_and_ReLU[10].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$2383(.Z({ \dot_product_and_ReLU[10].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$2384(.Z({ \dot_product_and_ReLU[10].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$2385(.Z({ \dot_product_and_ReLU[10].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$2386(.Z({ \dot_product_and_ReLU[10].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$2387(.Z({ \dot_product_and_ReLU[10].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$2388(.Z({ \dot_product_and_ReLU[10].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$2389(.Z({ \dot_product_and_ReLU[10].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$2390(.Z({ \dot_product_and_ReLU[10].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$2391(.Z({ \dot_product_and_ReLU[10].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$2392(.Z({ \dot_product_and_ReLU[10].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$2393(.Z({ \dot_product_and_ReLU[10].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$2394(.Z({ \dot_product_and_ReLU[10].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$2395(.Z({ \dot_product_and_ReLU[10].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$2396(.Z({ \dot_product_and_ReLU[10].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$2397(.Z({ \dot_product_and_ReLU[10].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$2398(.Z({ \dot_product_and_ReLU[10].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$2399(.Z({ \dot_product_and_ReLU[10].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$2400(.Z({ \dot_product_and_ReLU[10].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$2401(.Z({ \dot_product_and_ReLU[10].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$2402(.Z({ \dot_product_and_ReLU[10].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$2403(.Z({ \dot_product_and_ReLU[10].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$2404(.Z({ \dot_product_and_ReLU[10].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$2405(.Z({ \dot_product_and_ReLU[10].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$2406(.Z({ \dot_product_and_ReLU[10].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$2407(.Z({ \dot_product_and_ReLU[10].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$2408(.Z({ \dot_product_and_ReLU[10].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$2409(.Z({ \dot_product_and_ReLU[10].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$2410(.Z({ \dot_product_and_ReLU[10].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$2411(.Z({ \dot_product_and_ReLU[10].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$2412(.Z({ \dot_product_and_ReLU[10].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$2413(.Z({ \dot_product_and_ReLU[10].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$2414(.Z({ \dot_product_and_ReLU[10].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$2415(.Z({ \dot_product_and_ReLU[10].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$2416(.Z({ \dot_product_and_ReLU[10].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$2417(.Z({ \dot_product_and_ReLU[10].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$2418(.Z({ \dot_product_and_ReLU[10].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$2419(.Z({ \dot_product_and_ReLU[10].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$2420(.Z({ \dot_product_and_ReLU[10].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$2421(.Z({ \dot_product_and_ReLU[10].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$2422(.Z({ \dot_product_and_ReLU[10].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$2423(.Z({ \dot_product_and_ReLU[10].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$2424(.Z({ \dot_product_and_ReLU[10].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$2425(.Z({ \dot_product_and_ReLU[10].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$2426(.Z({ \dot_product_and_ReLU[10].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$2427(.Z({ \dot_product_and_ReLU[10].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$2428(.Z({ \dot_product_and_ReLU[10].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$2429(.Z({ \dot_product_and_ReLU[10].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$2430(.Z({ \dot_product_and_ReLU[10].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$2431(.Z({ \dot_product_and_ReLU[10].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$2432(.Z({ \dot_product_and_ReLU[10].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$2433(.Z({ \dot_product_and_ReLU[10].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$2434(.Z({ \dot_product_and_ReLU[10].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$2435(.Z({ \dot_product_and_ReLU[10].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$2436(.Z({ \dot_product_and_ReLU[10].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$2437(.Z({ \dot_product_and_ReLU[10].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$2438(.Z({ \dot_product_and_ReLU[10].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$2439(.Z({ \dot_product_and_ReLU[10].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$2440(.Z({ \dot_product_and_ReLU[10].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$2441(.Z({ \dot_product_and_ReLU[10].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$2442(.Z({ \dot_product_and_ReLU[10].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$2443(.Z({ \dot_product_and_ReLU[10].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$2444(.Z({ \dot_product_and_ReLU[10].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$2445(.Z({ \dot_product_and_ReLU[10].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$2446(.Z({ \dot_product_and_ReLU[10].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$2447(.Z({ \dot_product_and_ReLU[10].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$2448(.Z({ \dot_product_and_ReLU[10].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$2449(.Z({ \dot_product_and_ReLU[10].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$2450(.Z({ \dot_product_and_ReLU[10].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$2451(.Z({ \dot_product_and_ReLU[10].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$2452(.Z({ \dot_product_and_ReLU[10].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$2453(.Z({ \dot_product_and_ReLU[10].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$2454(.Z({ \dot_product_and_ReLU[10].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$2455(.Z({ \dot_product_and_ReLU[10].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$2456(.Z({ \dot_product_and_ReLU[10].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$2457(.Z({ \dot_product_and_ReLU[10].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$2458(.Z({ \dot_product_and_ReLU[10].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$2459(.Z({ \dot_product_and_ReLU[10].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$2460(.Z({ \dot_product_and_ReLU[10].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$2461(.Z({ \dot_product_and_ReLU[10].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$2462(.Z({ \dot_product_and_ReLU[10].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$2463(.Z({ \dot_product_and_ReLU[10].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$2464(.Z({ \dot_product_and_ReLU[10].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$2465(.Z({ \dot_product_and_ReLU[10].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$2466(.Z({ \dot_product_and_ReLU[10].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$2467(.Z({ \dot_product_and_ReLU[10].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$2468(.Z({ \dot_product_and_ReLU[10].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$2469(.Z({ \dot_product_and_ReLU[10].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$2470(.Z({ \dot_product_and_ReLU[10].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$2471(.Z({ \dot_product_and_ReLU[10].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$2472(.Z({ \dot_product_and_ReLU[10].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$2473(.Z({ \dot_product_and_ReLU[10].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$2474(.Z({ \dot_product_and_ReLU[10].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$2475(.Z({ \dot_product_and_ReLU[10].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$2476(.Z({ \dot_product_and_ReLU[10].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$2477(.Z({ \dot_product_and_ReLU[10].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$2478(.Z({ \dot_product_and_ReLU[10].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$2479(.Z({ \dot_product_and_ReLU[10].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$2480(.Z({ \dot_product_and_ReLU[10].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$2481(.Z({ \dot_product_and_ReLU[10].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$2482(.Z({ \dot_product_and_ReLU[10].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$2483(.Z({ \dot_product_and_ReLU[10].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$2484(.Z({ \dot_product_and_ReLU[10].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$2485(.Z({ \dot_product_and_ReLU[10].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$2486(.Z({ \dot_product_and_ReLU[10].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$2487(.Z({ \dot_product_and_ReLU[10].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$2488(.Z({ \dot_product_and_ReLU[10].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$2489(.Z({ \dot_product_and_ReLU[10].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$2490(.Z({ \dot_product_and_ReLU[10].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$2491(.Z({ \dot_product_and_ReLU[10].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$2492(.Z({ \dot_product_and_ReLU[10].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$2493(.Z({ \dot_product_and_ReLU[10].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$2494(.Z({ \dot_product_and_ReLU[10].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$2495(.Z({ \dot_product_and_ReLU[10].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$2496(.Z({ \dot_product_and_ReLU[10].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$2497(.Z({ \dot_product_and_ReLU[10].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$2498(.Z({ \dot_product_and_ReLU[10].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$2499(.Z({ \dot_product_and_ReLU[10].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$2500(.Z({ \dot_product_and_ReLU[10].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$2501(.Z({ \dot_product_and_ReLU[10].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$2502(.Z({ \dot_product_and_ReLU[10].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$2503(.Z({ \dot_product_and_ReLU[10].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$2504(.Z({ \dot_product_and_ReLU[10].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$2505(.Z({ \dot_product_and_ReLU[10].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$2506(.Z({ \dot_product_and_ReLU[10].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$2507(.Z({ \dot_product_and_ReLU[10].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$2508(.Z({ \dot_product_and_ReLU[10].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$2509(.Z({ \dot_product_and_ReLU[10].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$2510(.Z({ \dot_product_and_ReLU[10].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$2511(.Z({ \dot_product_and_ReLU[10].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$2512(.Z({ \dot_product_and_ReLU[10].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$2513(.Z({ \dot_product_and_ReLU[10].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$2514(.Z({ \dot_product_and_ReLU[10].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$2515(.Z({ \dot_product_and_ReLU[10].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$2516(.Z({ \dot_product_and_ReLU[10].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$2517(.Z({ \dot_product_and_ReLU[10].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$2518(.Z({ \dot_product_and_ReLU[10].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$2519(.Z({ \dot_product_and_ReLU[10].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$2520(.Z({ \dot_product_and_ReLU[10].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$2521(.Z({ \dot_product_and_ReLU[10].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$2522(.Z({ \dot_product_and_ReLU[10].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$2523(.Z({ \dot_product_and_ReLU[10].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$2524(.Z({ \dot_product_and_ReLU[10].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$2525(.Z({ \dot_product_and_ReLU[10].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$2526(.Z({ \dot_product_and_ReLU[10].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$2527(.Z({ \dot_product_and_ReLU[10].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$2528(.Z({ \dot_product_and_ReLU[10].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$2529(.Z({ \dot_product_and_ReLU[10].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$2530(.Z({ \dot_product_and_ReLU[10].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$2531(.Z({ \dot_product_and_ReLU[10].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$2532(.Z({ \dot_product_and_ReLU[10].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$2533(.Z({ \dot_product_and_ReLU[10].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$2534(.Z({ \dot_product_and_ReLU[10].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$2535(.Z({ \dot_product_and_ReLU[10].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$2536(.Z({ \dot_product_and_ReLU[10].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$2537(.Z({ \dot_product_and_ReLU[10].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$2538(.Z({ \dot_product_and_ReLU[10].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$2539(.Z({ \dot_product_and_ReLU[10].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$2540(.Z({ \dot_product_and_ReLU[10].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$2541(.Z({ \dot_product_and_ReLU[10].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$2542(.Z({ \dot_product_and_ReLU[10].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$2543(.Z({ \dot_product_and_ReLU[10].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$2544(.Z({ \dot_product_and_ReLU[10].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$2545(.Z({ \dot_product_and_ReLU[10].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$2546(.Z({ \dot_product_and_ReLU[10].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$2547(.Z({ \dot_product_and_ReLU[10].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$2548(.Z({ \dot_product_and_ReLU[10].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$2549(.Z({ \dot_product_and_ReLU[10].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$2550(.Z({ \dot_product_and_ReLU[10].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$2551(.Z({ \dot_product_and_ReLU[10].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$2552(.Z({ \dot_product_and_ReLU[10].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$2553(.Z({ \dot_product_and_ReLU[10].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$2554(.Z({ \dot_product_and_ReLU[10].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$2555(.Z({ \dot_product_and_ReLU[10].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$2556(.Z({ \dot_product_and_ReLU[10].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$2557(.Z({ \dot_product_and_ReLU[10].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$2558(.Z({ \dot_product_and_ReLU[10].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$2559(.Z({ \dot_product_and_ReLU[10].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$2560(.Z({ \dot_product_and_ReLU[10].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[10][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$2561(.Z({ \dot_product_and_ReLU[9].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$2562(.Z({ \dot_product_and_ReLU[9].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$2563(.Z({ \dot_product_and_ReLU[9].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$2564(.Z({ \dot_product_and_ReLU[9].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$2565(.Z({ \dot_product_and_ReLU[9].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$2566(.Z({ \dot_product_and_ReLU[9].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$2567(.Z({ \dot_product_and_ReLU[9].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$2568(.Z({ \dot_product_and_ReLU[9].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$2569(.Z({ \dot_product_and_ReLU[9].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$2570(.Z({ \dot_product_and_ReLU[9].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$2571(.Z({ \dot_product_and_ReLU[9].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$2572(.Z({ \dot_product_and_ReLU[9].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$2573(.Z({ \dot_product_and_ReLU[9].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$2574(.Z({ \dot_product_and_ReLU[9].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$2575(.Z({ \dot_product_and_ReLU[9].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$2576(.Z({ \dot_product_and_ReLU[9].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$2577(.Z({ \dot_product_and_ReLU[9].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$2578(.Z({ \dot_product_and_ReLU[9].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$2579(.Z({ \dot_product_and_ReLU[9].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$2580(.Z({ \dot_product_and_ReLU[9].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$2581(.Z({ \dot_product_and_ReLU[9].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$2582(.Z({ \dot_product_and_ReLU[9].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$2583(.Z({ \dot_product_and_ReLU[9].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$2584(.Z({ \dot_product_and_ReLU[9].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$2585(.Z({ \dot_product_and_ReLU[9].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$2586(.Z({ \dot_product_and_ReLU[9].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$2587(.Z({ \dot_product_and_ReLU[9].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$2588(.Z({ \dot_product_and_ReLU[9].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$2589(.Z({ \dot_product_and_ReLU[9].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$2590(.Z({ \dot_product_and_ReLU[9].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$2591(.Z({ \dot_product_and_ReLU[9].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$2592(.Z({ \dot_product_and_ReLU[9].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$2593(.Z({ \dot_product_and_ReLU[9].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$2594(.Z({ \dot_product_and_ReLU[9].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$2595(.Z({ \dot_product_and_ReLU[9].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$2596(.Z({ \dot_product_and_ReLU[9].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$2597(.Z({ \dot_product_and_ReLU[9].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$2598(.Z({ \dot_product_and_ReLU[9].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$2599(.Z({ \dot_product_and_ReLU[9].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$2600(.Z({ \dot_product_and_ReLU[9].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$2601(.Z({ \dot_product_and_ReLU[9].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$2602(.Z({ \dot_product_and_ReLU[9].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$2603(.Z({ \dot_product_and_ReLU[9].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$2604(.Z({ \dot_product_and_ReLU[9].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$2605(.Z({ \dot_product_and_ReLU[9].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$2606(.Z({ \dot_product_and_ReLU[9].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$2607(.Z({ \dot_product_and_ReLU[9].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$2608(.Z({ \dot_product_and_ReLU[9].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$2609(.Z({ \dot_product_and_ReLU[9].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$2610(.Z({ \dot_product_and_ReLU[9].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$2611(.Z({ \dot_product_and_ReLU[9].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$2612(.Z({ \dot_product_and_ReLU[9].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$2613(.Z({ \dot_product_and_ReLU[9].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$2614(.Z({ \dot_product_and_ReLU[9].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$2615(.Z({ \dot_product_and_ReLU[9].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$2616(.Z({ \dot_product_and_ReLU[9].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$2617(.Z({ \dot_product_and_ReLU[9].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$2618(.Z({ \dot_product_and_ReLU[9].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$2619(.Z({ \dot_product_and_ReLU[9].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$2620(.Z({ \dot_product_and_ReLU[9].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$2621(.Z({ \dot_product_and_ReLU[9].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$2622(.Z({ \dot_product_and_ReLU[9].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$2623(.Z({ \dot_product_and_ReLU[9].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$2624(.Z({ \dot_product_and_ReLU[9].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$2625(.Z({ \dot_product_and_ReLU[9].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$2626(.Z({ \dot_product_and_ReLU[9].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$2627(.Z({ \dot_product_and_ReLU[9].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$2628(.Z({ \dot_product_and_ReLU[9].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$2629(.Z({ \dot_product_and_ReLU[9].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$2630(.Z({ \dot_product_and_ReLU[9].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$2631(.Z({ \dot_product_and_ReLU[9].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$2632(.Z({ \dot_product_and_ReLU[9].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$2633(.Z({ \dot_product_and_ReLU[9].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$2634(.Z({ \dot_product_and_ReLU[9].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$2635(.Z({ \dot_product_and_ReLU[9].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$2636(.Z({ \dot_product_and_ReLU[9].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$2637(.Z({ \dot_product_and_ReLU[9].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$2638(.Z({ \dot_product_and_ReLU[9].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$2639(.Z({ \dot_product_and_ReLU[9].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$2640(.Z({ \dot_product_and_ReLU[9].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$2641(.Z({ \dot_product_and_ReLU[9].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$2642(.Z({ \dot_product_and_ReLU[9].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$2643(.Z({ \dot_product_and_ReLU[9].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$2644(.Z({ \dot_product_and_ReLU[9].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$2645(.Z({ \dot_product_and_ReLU[9].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$2646(.Z({ \dot_product_and_ReLU[9].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$2647(.Z({ \dot_product_and_ReLU[9].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$2648(.Z({ \dot_product_and_ReLU[9].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$2649(.Z({ \dot_product_and_ReLU[9].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$2650(.Z({ \dot_product_and_ReLU[9].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$2651(.Z({ \dot_product_and_ReLU[9].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$2652(.Z({ \dot_product_and_ReLU[9].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$2653(.Z({ \dot_product_and_ReLU[9].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$2654(.Z({ \dot_product_and_ReLU[9].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$2655(.Z({ \dot_product_and_ReLU[9].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$2656(.Z({ \dot_product_and_ReLU[9].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$2657(.Z({ \dot_product_and_ReLU[9].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$2658(.Z({ \dot_product_and_ReLU[9].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$2659(.Z({ \dot_product_and_ReLU[9].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$2660(.Z({ \dot_product_and_ReLU[9].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$2661(.Z({ \dot_product_and_ReLU[9].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$2662(.Z({ \dot_product_and_ReLU[9].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$2663(.Z({ \dot_product_and_ReLU[9].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$2664(.Z({ \dot_product_and_ReLU[9].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$2665(.Z({ \dot_product_and_ReLU[9].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$2666(.Z({ \dot_product_and_ReLU[9].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$2667(.Z({ \dot_product_and_ReLU[9].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$2668(.Z({ \dot_product_and_ReLU[9].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$2669(.Z({ \dot_product_and_ReLU[9].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$2670(.Z({ \dot_product_and_ReLU[9].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$2671(.Z({ \dot_product_and_ReLU[9].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$2672(.Z({ \dot_product_and_ReLU[9].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$2673(.Z({ \dot_product_and_ReLU[9].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$2674(.Z({ \dot_product_and_ReLU[9].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$2675(.Z({ \dot_product_and_ReLU[9].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$2676(.Z({ \dot_product_and_ReLU[9].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$2677(.Z({ \dot_product_and_ReLU[9].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$2678(.Z({ \dot_product_and_ReLU[9].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$2679(.Z({ \dot_product_and_ReLU[9].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$2680(.Z({ \dot_product_and_ReLU[9].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$2681(.Z({ \dot_product_and_ReLU[9].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$2682(.Z({ \dot_product_and_ReLU[9].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$2683(.Z({ \dot_product_and_ReLU[9].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$2684(.Z({ \dot_product_and_ReLU[9].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$2685(.Z({ \dot_product_and_ReLU[9].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$2686(.Z({ \dot_product_and_ReLU[9].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$2687(.Z({ \dot_product_and_ReLU[9].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$2688(.Z({ \dot_product_and_ReLU[9].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$2689(.Z({ \dot_product_and_ReLU[9].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$2690(.Z({ \dot_product_and_ReLU[9].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$2691(.Z({ \dot_product_and_ReLU[9].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$2692(.Z({ \dot_product_and_ReLU[9].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$2693(.Z({ \dot_product_and_ReLU[9].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$2694(.Z({ \dot_product_and_ReLU[9].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$2695(.Z({ \dot_product_and_ReLU[9].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$2696(.Z({ \dot_product_and_ReLU[9].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$2697(.Z({ \dot_product_and_ReLU[9].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$2698(.Z({ \dot_product_and_ReLU[9].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$2699(.Z({ \dot_product_and_ReLU[9].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$2700(.Z({ \dot_product_and_ReLU[9].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$2701(.Z({ \dot_product_and_ReLU[9].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$2702(.Z({ \dot_product_and_ReLU[9].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$2703(.Z({ \dot_product_and_ReLU[9].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$2704(.Z({ \dot_product_and_ReLU[9].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$2705(.Z({ \dot_product_and_ReLU[9].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$2706(.Z({ \dot_product_and_ReLU[9].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$2707(.Z({ \dot_product_and_ReLU[9].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$2708(.Z({ \dot_product_and_ReLU[9].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$2709(.Z({ \dot_product_and_ReLU[9].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$2710(.Z({ \dot_product_and_ReLU[9].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$2711(.Z({ \dot_product_and_ReLU[9].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$2712(.Z({ \dot_product_and_ReLU[9].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$2713(.Z({ \dot_product_and_ReLU[9].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$2714(.Z({ \dot_product_and_ReLU[9].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$2715(.Z({ \dot_product_and_ReLU[9].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$2716(.Z({ \dot_product_and_ReLU[9].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$2717(.Z({ \dot_product_and_ReLU[9].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$2718(.Z({ \dot_product_and_ReLU[9].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$2719(.Z({ \dot_product_and_ReLU[9].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$2720(.Z({ \dot_product_and_ReLU[9].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$2721(.Z({ \dot_product_and_ReLU[9].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$2722(.Z({ \dot_product_and_ReLU[9].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$2723(.Z({ \dot_product_and_ReLU[9].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$2724(.Z({ \dot_product_and_ReLU[9].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$2725(.Z({ \dot_product_and_ReLU[9].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$2726(.Z({ \dot_product_and_ReLU[9].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$2727(.Z({ \dot_product_and_ReLU[9].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$2728(.Z({ \dot_product_and_ReLU[9].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$2729(.Z({ \dot_product_and_ReLU[9].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$2730(.Z({ \dot_product_and_ReLU[9].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$2731(.Z({ \dot_product_and_ReLU[9].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$2732(.Z({ \dot_product_and_ReLU[9].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$2733(.Z({ \dot_product_and_ReLU[9].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$2734(.Z({ \dot_product_and_ReLU[9].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$2735(.Z({ \dot_product_and_ReLU[9].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$2736(.Z({ \dot_product_and_ReLU[9].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$2737(.Z({ \dot_product_and_ReLU[9].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$2738(.Z({ \dot_product_and_ReLU[9].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$2739(.Z({ \dot_product_and_ReLU[9].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$2740(.Z({ \dot_product_and_ReLU[9].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$2741(.Z({ \dot_product_and_ReLU[9].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$2742(.Z({ \dot_product_and_ReLU[9].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$2743(.Z({ \dot_product_and_ReLU[9].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$2744(.Z({ \dot_product_and_ReLU[9].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$2745(.Z({ \dot_product_and_ReLU[9].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$2746(.Z({ \dot_product_and_ReLU[9].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$2747(.Z({ \dot_product_and_ReLU[9].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$2748(.Z({ \dot_product_and_ReLU[9].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$2749(.Z({ \dot_product_and_ReLU[9].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$2750(.Z({ \dot_product_and_ReLU[9].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$2751(.Z({ \dot_product_and_ReLU[9].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$2752(.Z({ \dot_product_and_ReLU[9].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$2753(.Z({ \dot_product_and_ReLU[9].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$2754(.Z({ \dot_product_and_ReLU[9].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$2755(.Z({ \dot_product_and_ReLU[9].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$2756(.Z({ \dot_product_and_ReLU[9].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$2757(.Z({ \dot_product_and_ReLU[9].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$2758(.Z({ \dot_product_and_ReLU[9].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$2759(.Z({ \dot_product_and_ReLU[9].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$2760(.Z({ \dot_product_and_ReLU[9].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$2761(.Z({ \dot_product_and_ReLU[9].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$2762(.Z({ \dot_product_and_ReLU[9].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$2763(.Z({ \dot_product_and_ReLU[9].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$2764(.Z({ \dot_product_and_ReLU[9].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$2765(.Z({ \dot_product_and_ReLU[9].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$2766(.Z({ \dot_product_and_ReLU[9].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$2767(.Z({ \dot_product_and_ReLU[9].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$2768(.Z({ \dot_product_and_ReLU[9].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$2769(.Z({ \dot_product_and_ReLU[9].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$2770(.Z({ \dot_product_and_ReLU[9].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$2771(.Z({ \dot_product_and_ReLU[9].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$2772(.Z({ \dot_product_and_ReLU[9].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$2773(.Z({ \dot_product_and_ReLU[9].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$2774(.Z({ \dot_product_and_ReLU[9].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$2775(.Z({ \dot_product_and_ReLU[9].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$2776(.Z({ \dot_product_and_ReLU[9].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$2777(.Z({ \dot_product_and_ReLU[9].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$2778(.Z({ \dot_product_and_ReLU[9].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$2779(.Z({ \dot_product_and_ReLU[9].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$2780(.Z({ \dot_product_and_ReLU[9].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$2781(.Z({ \dot_product_and_ReLU[9].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$2782(.Z({ \dot_product_and_ReLU[9].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$2783(.Z({ \dot_product_and_ReLU[9].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$2784(.Z({ \dot_product_and_ReLU[9].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$2785(.Z({ \dot_product_and_ReLU[9].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$2786(.Z({ \dot_product_and_ReLU[9].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$2787(.Z({ \dot_product_and_ReLU[9].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$2788(.Z({ \dot_product_and_ReLU[9].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$2789(.Z({ \dot_product_and_ReLU[9].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$2790(.Z({ \dot_product_and_ReLU[9].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$2791(.Z({ \dot_product_and_ReLU[9].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$2792(.Z({ \dot_product_and_ReLU[9].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$2793(.Z({ \dot_product_and_ReLU[9].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$2794(.Z({ \dot_product_and_ReLU[9].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$2795(.Z({ \dot_product_and_ReLU[9].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$2796(.Z({ \dot_product_and_ReLU[9].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$2797(.Z({ \dot_product_and_ReLU[9].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$2798(.Z({ \dot_product_and_ReLU[9].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$2799(.Z({ \dot_product_and_ReLU[9].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$2800(.Z({ \dot_product_and_ReLU[9].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$2801(.Z({ \dot_product_and_ReLU[9].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$2802(.Z({ \dot_product_and_ReLU[9].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$2803(.Z({ \dot_product_and_ReLU[9].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$2804(.Z({ \dot_product_and_ReLU[9].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$2805(.Z({ \dot_product_and_ReLU[9].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$2806(.Z({ \dot_product_and_ReLU[9].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$2807(.Z({ \dot_product_and_ReLU[9].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$2808(.Z({ \dot_product_and_ReLU[9].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$2809(.Z({ \dot_product_and_ReLU[9].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$2810(.Z({ \dot_product_and_ReLU[9].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$2811(.Z({ \dot_product_and_ReLU[9].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$2812(.Z({ \dot_product_and_ReLU[9].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$2813(.Z({ \dot_product_and_ReLU[9].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$2814(.Z({ \dot_product_and_ReLU[9].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$2815(.Z({ \dot_product_and_ReLU[9].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$2816(.Z({ \dot_product_and_ReLU[9].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[9][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$2817(.Z({ \dot_product_and_ReLU[8].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$2818(.Z({ \dot_product_and_ReLU[8].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$2819(.Z({ \dot_product_and_ReLU[8].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$2820(.Z({ \dot_product_and_ReLU[8].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$2821(.Z({ \dot_product_and_ReLU[8].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$2822(.Z({ \dot_product_and_ReLU[8].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$2823(.Z({ \dot_product_and_ReLU[8].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$2824(.Z({ \dot_product_and_ReLU[8].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$2825(.Z({ \dot_product_and_ReLU[8].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$2826(.Z({ \dot_product_and_ReLU[8].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$2827(.Z({ \dot_product_and_ReLU[8].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$2828(.Z({ \dot_product_and_ReLU[8].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$2829(.Z({ \dot_product_and_ReLU[8].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$2830(.Z({ \dot_product_and_ReLU[8].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$2831(.Z({ \dot_product_and_ReLU[8].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$2832(.Z({ \dot_product_and_ReLU[8].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$2833(.Z({ \dot_product_and_ReLU[8].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$2834(.Z({ \dot_product_and_ReLU[8].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$2835(.Z({ \dot_product_and_ReLU[8].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$2836(.Z({ \dot_product_and_ReLU[8].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$2837(.Z({ \dot_product_and_ReLU[8].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$2838(.Z({ \dot_product_and_ReLU[8].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$2839(.Z({ \dot_product_and_ReLU[8].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$2840(.Z({ \dot_product_and_ReLU[8].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$2841(.Z({ \dot_product_and_ReLU[8].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$2842(.Z({ \dot_product_and_ReLU[8].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$2843(.Z({ \dot_product_and_ReLU[8].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$2844(.Z({ \dot_product_and_ReLU[8].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$2845(.Z({ \dot_product_and_ReLU[8].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$2846(.Z({ \dot_product_and_ReLU[8].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$2847(.Z({ \dot_product_and_ReLU[8].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$2848(.Z({ \dot_product_and_ReLU[8].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$2849(.Z({ \dot_product_and_ReLU[8].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$2850(.Z({ \dot_product_and_ReLU[8].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$2851(.Z({ \dot_product_and_ReLU[8].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$2852(.Z({ \dot_product_and_ReLU[8].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$2853(.Z({ \dot_product_and_ReLU[8].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$2854(.Z({ \dot_product_and_ReLU[8].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$2855(.Z({ \dot_product_and_ReLU[8].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$2856(.Z({ \dot_product_and_ReLU[8].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$2857(.Z({ \dot_product_and_ReLU[8].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$2858(.Z({ \dot_product_and_ReLU[8].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$2859(.Z({ \dot_product_and_ReLU[8].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$2860(.Z({ \dot_product_and_ReLU[8].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$2861(.Z({ \dot_product_and_ReLU[8].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$2862(.Z({ \dot_product_and_ReLU[8].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$2863(.Z({ \dot_product_and_ReLU[8].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$2864(.Z({ \dot_product_and_ReLU[8].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$2865(.Z({ \dot_product_and_ReLU[8].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$2866(.Z({ \dot_product_and_ReLU[8].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$2867(.Z({ \dot_product_and_ReLU[8].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$2868(.Z({ \dot_product_and_ReLU[8].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$2869(.Z({ \dot_product_and_ReLU[8].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$2870(.Z({ \dot_product_and_ReLU[8].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$2871(.Z({ \dot_product_and_ReLU[8].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$2872(.Z({ \dot_product_and_ReLU[8].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$2873(.Z({ \dot_product_and_ReLU[8].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$2874(.Z({ \dot_product_and_ReLU[8].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$2875(.Z({ \dot_product_and_ReLU[8].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$2876(.Z({ \dot_product_and_ReLU[8].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$2877(.Z({ \dot_product_and_ReLU[8].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$2878(.Z({ \dot_product_and_ReLU[8].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$2879(.Z({ \dot_product_and_ReLU[8].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$2880(.Z({ \dot_product_and_ReLU[8].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$2881(.Z({ \dot_product_and_ReLU[8].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$2882(.Z({ \dot_product_and_ReLU[8].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$2883(.Z({ \dot_product_and_ReLU[8].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$2884(.Z({ \dot_product_and_ReLU[8].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$2885(.Z({ \dot_product_and_ReLU[8].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$2886(.Z({ \dot_product_and_ReLU[8].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$2887(.Z({ \dot_product_and_ReLU[8].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$2888(.Z({ \dot_product_and_ReLU[8].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$2889(.Z({ \dot_product_and_ReLU[8].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$2890(.Z({ \dot_product_and_ReLU[8].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$2891(.Z({ \dot_product_and_ReLU[8].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$2892(.Z({ \dot_product_and_ReLU[8].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$2893(.Z({ \dot_product_and_ReLU[8].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$2894(.Z({ \dot_product_and_ReLU[8].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$2895(.Z({ \dot_product_and_ReLU[8].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$2896(.Z({ \dot_product_and_ReLU[8].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$2897(.Z({ \dot_product_and_ReLU[8].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$2898(.Z({ \dot_product_and_ReLU[8].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$2899(.Z({ \dot_product_and_ReLU[8].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$2900(.Z({ \dot_product_and_ReLU[8].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$2901(.Z({ \dot_product_and_ReLU[8].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$2902(.Z({ \dot_product_and_ReLU[8].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$2903(.Z({ \dot_product_and_ReLU[8].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$2904(.Z({ \dot_product_and_ReLU[8].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$2905(.Z({ \dot_product_and_ReLU[8].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$2906(.Z({ \dot_product_and_ReLU[8].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$2907(.Z({ \dot_product_and_ReLU[8].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$2908(.Z({ \dot_product_and_ReLU[8].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$2909(.Z({ \dot_product_and_ReLU[8].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$2910(.Z({ \dot_product_and_ReLU[8].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$2911(.Z({ \dot_product_and_ReLU[8].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$2912(.Z({ \dot_product_and_ReLU[8].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$2913(.Z({ \dot_product_and_ReLU[8].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$2914(.Z({ \dot_product_and_ReLU[8].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$2915(.Z({ \dot_product_and_ReLU[8].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$2916(.Z({ \dot_product_and_ReLU[8].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$2917(.Z({ \dot_product_and_ReLU[8].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$2918(.Z({ \dot_product_and_ReLU[8].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$2919(.Z({ \dot_product_and_ReLU[8].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$2920(.Z({ \dot_product_and_ReLU[8].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$2921(.Z({ \dot_product_and_ReLU[8].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$2922(.Z({ \dot_product_and_ReLU[8].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$2923(.Z({ \dot_product_and_ReLU[8].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$2924(.Z({ \dot_product_and_ReLU[8].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$2925(.Z({ \dot_product_and_ReLU[8].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$2926(.Z({ \dot_product_and_ReLU[8].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$2927(.Z({ \dot_product_and_ReLU[8].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$2928(.Z({ \dot_product_and_ReLU[8].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$2929(.Z({ \dot_product_and_ReLU[8].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$2930(.Z({ \dot_product_and_ReLU[8].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$2931(.Z({ \dot_product_and_ReLU[8].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$2932(.Z({ \dot_product_and_ReLU[8].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$2933(.Z({ \dot_product_and_ReLU[8].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$2934(.Z({ \dot_product_and_ReLU[8].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$2935(.Z({ \dot_product_and_ReLU[8].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$2936(.Z({ \dot_product_and_ReLU[8].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$2937(.Z({ \dot_product_and_ReLU[8].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$2938(.Z({ \dot_product_and_ReLU[8].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$2939(.Z({ \dot_product_and_ReLU[8].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$2940(.Z({ \dot_product_and_ReLU[8].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$2941(.Z({ \dot_product_and_ReLU[8].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$2942(.Z({ \dot_product_and_ReLU[8].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$2943(.Z({ \dot_product_and_ReLU[8].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$2944(.Z({ \dot_product_and_ReLU[8].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$2945(.Z({ \dot_product_and_ReLU[8].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$2946(.Z({ \dot_product_and_ReLU[8].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$2947(.Z({ \dot_product_and_ReLU[8].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$2948(.Z({ \dot_product_and_ReLU[8].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$2949(.Z({ \dot_product_and_ReLU[8].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$2950(.Z({ \dot_product_and_ReLU[8].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$2951(.Z({ \dot_product_and_ReLU[8].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$2952(.Z({ \dot_product_and_ReLU[8].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$2953(.Z({ \dot_product_and_ReLU[8].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$2954(.Z({ \dot_product_and_ReLU[8].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$2955(.Z({ \dot_product_and_ReLU[8].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$2956(.Z({ \dot_product_and_ReLU[8].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$2957(.Z({ \dot_product_and_ReLU[8].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$2958(.Z({ \dot_product_and_ReLU[8].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$2959(.Z({ \dot_product_and_ReLU[8].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$2960(.Z({ \dot_product_and_ReLU[8].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$2961(.Z({ \dot_product_and_ReLU[8].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$2962(.Z({ \dot_product_and_ReLU[8].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$2963(.Z({ \dot_product_and_ReLU[8].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$2964(.Z({ \dot_product_and_ReLU[8].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$2965(.Z({ \dot_product_and_ReLU[8].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$2966(.Z({ \dot_product_and_ReLU[8].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$2967(.Z({ \dot_product_and_ReLU[8].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$2968(.Z({ \dot_product_and_ReLU[8].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$2969(.Z({ \dot_product_and_ReLU[8].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$2970(.Z({ \dot_product_and_ReLU[8].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$2971(.Z({ \dot_product_and_ReLU[8].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$2972(.Z({ \dot_product_and_ReLU[8].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$2973(.Z({ \dot_product_and_ReLU[8].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$2974(.Z({ \dot_product_and_ReLU[8].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$2975(.Z({ \dot_product_and_ReLU[8].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$2976(.Z({ \dot_product_and_ReLU[8].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$2977(.Z({ \dot_product_and_ReLU[8].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$2978(.Z({ \dot_product_and_ReLU[8].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$2979(.Z({ \dot_product_and_ReLU[8].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$2980(.Z({ \dot_product_and_ReLU[8].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$2981(.Z({ \dot_product_and_ReLU[8].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$2982(.Z({ \dot_product_and_ReLU[8].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$2983(.Z({ \dot_product_and_ReLU[8].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$2984(.Z({ \dot_product_and_ReLU[8].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$2985(.Z({ \dot_product_and_ReLU[8].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$2986(.Z({ \dot_product_and_ReLU[8].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$2987(.Z({ \dot_product_and_ReLU[8].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$2988(.Z({ \dot_product_and_ReLU[8].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$2989(.Z({ \dot_product_and_ReLU[8].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$2990(.Z({ \dot_product_and_ReLU[8].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$2991(.Z({ \dot_product_and_ReLU[8].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$2992(.Z({ \dot_product_and_ReLU[8].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$2993(.Z({ \dot_product_and_ReLU[8].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$2994(.Z({ \dot_product_and_ReLU[8].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$2995(.Z({ \dot_product_and_ReLU[8].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$2996(.Z({ \dot_product_and_ReLU[8].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$2997(.Z({ \dot_product_and_ReLU[8].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$2998(.Z({ \dot_product_and_ReLU[8].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$2999(.Z({ \dot_product_and_ReLU[8].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$3000(.Z({ \dot_product_and_ReLU[8].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$3001(.Z({ \dot_product_and_ReLU[8].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$3002(.Z({ \dot_product_and_ReLU[8].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$3003(.Z({ \dot_product_and_ReLU[8].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$3004(.Z({ \dot_product_and_ReLU[8].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$3005(.Z({ \dot_product_and_ReLU[8].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$3006(.Z({ \dot_product_and_ReLU[8].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$3007(.Z({ \dot_product_and_ReLU[8].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$3008(.Z({ \dot_product_and_ReLU[8].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$3009(.Z({ \dot_product_and_ReLU[8].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$3010(.Z({ \dot_product_and_ReLU[8].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$3011(.Z({ \dot_product_and_ReLU[8].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$3012(.Z({ \dot_product_and_ReLU[8].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$3013(.Z({ \dot_product_and_ReLU[8].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$3014(.Z({ \dot_product_and_ReLU[8].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$3015(.Z({ \dot_product_and_ReLU[8].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$3016(.Z({ \dot_product_and_ReLU[8].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$3017(.Z({ \dot_product_and_ReLU[8].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$3018(.Z({ \dot_product_and_ReLU[8].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$3019(.Z({ \dot_product_and_ReLU[8].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$3020(.Z({ \dot_product_and_ReLU[8].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$3021(.Z({ \dot_product_and_ReLU[8].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$3022(.Z({ \dot_product_and_ReLU[8].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$3023(.Z({ \dot_product_and_ReLU[8].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$3024(.Z({ \dot_product_and_ReLU[8].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$3025(.Z({ \dot_product_and_ReLU[8].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$3026(.Z({ \dot_product_and_ReLU[8].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$3027(.Z({ \dot_product_and_ReLU[8].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$3028(.Z({ \dot_product_and_ReLU[8].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$3029(.Z({ \dot_product_and_ReLU[8].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$3030(.Z({ \dot_product_and_ReLU[8].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$3031(.Z({ \dot_product_and_ReLU[8].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$3032(.Z({ \dot_product_and_ReLU[8].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$3033(.Z({ \dot_product_and_ReLU[8].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$3034(.Z({ \dot_product_and_ReLU[8].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$3035(.Z({ \dot_product_and_ReLU[8].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$3036(.Z({ \dot_product_and_ReLU[8].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$3037(.Z({ \dot_product_and_ReLU[8].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$3038(.Z({ \dot_product_and_ReLU[8].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$3039(.Z({ \dot_product_and_ReLU[8].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$3040(.Z({ \dot_product_and_ReLU[8].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$3041(.Z({ \dot_product_and_ReLU[8].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$3042(.Z({ \dot_product_and_ReLU[8].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$3043(.Z({ \dot_product_and_ReLU[8].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$3044(.Z({ \dot_product_and_ReLU[8].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$3045(.Z({ \dot_product_and_ReLU[8].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$3046(.Z({ \dot_product_and_ReLU[8].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$3047(.Z({ \dot_product_and_ReLU[8].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$3048(.Z({ \dot_product_and_ReLU[8].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$3049(.Z({ \dot_product_and_ReLU[8].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$3050(.Z({ \dot_product_and_ReLU[8].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$3051(.Z({ \dot_product_and_ReLU[8].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$3052(.Z({ \dot_product_and_ReLU[8].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$3053(.Z({ \dot_product_and_ReLU[8].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$3054(.Z({ \dot_product_and_ReLU[8].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$3055(.Z({ \dot_product_and_ReLU[8].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$3056(.Z({ \dot_product_and_ReLU[8].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$3057(.Z({ \dot_product_and_ReLU[8].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$3058(.Z({ \dot_product_and_ReLU[8].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$3059(.Z({ \dot_product_and_ReLU[8].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$3060(.Z({ \dot_product_and_ReLU[8].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$3061(.Z({ \dot_product_and_ReLU[8].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$3062(.Z({ \dot_product_and_ReLU[8].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$3063(.Z({ \dot_product_and_ReLU[8].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$3064(.Z({ \dot_product_and_ReLU[8].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$3065(.Z({ \dot_product_and_ReLU[8].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$3066(.Z({ \dot_product_and_ReLU[8].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$3067(.Z({ \dot_product_and_ReLU[8].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$3068(.Z({ \dot_product_and_ReLU[8].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$3069(.Z({ \dot_product_and_ReLU[8].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$3070(.Z({ \dot_product_and_ReLU[8].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$3071(.Z({ \dot_product_and_ReLU[8].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$3072(.Z({ \dot_product_and_ReLU[8].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[8][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$3073(.Z({ \dot_product_and_ReLU[7].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$3074(.Z({ \dot_product_and_ReLU[7].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$3075(.Z({ \dot_product_and_ReLU[7].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$3076(.Z({ \dot_product_and_ReLU[7].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$3077(.Z({ \dot_product_and_ReLU[7].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$3078(.Z({ \dot_product_and_ReLU[7].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$3079(.Z({ \dot_product_and_ReLU[7].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$3080(.Z({ \dot_product_and_ReLU[7].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$3081(.Z({ \dot_product_and_ReLU[7].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$3082(.Z({ \dot_product_and_ReLU[7].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$3083(.Z({ \dot_product_and_ReLU[7].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$3084(.Z({ \dot_product_and_ReLU[7].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$3085(.Z({ \dot_product_and_ReLU[7].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$3086(.Z({ \dot_product_and_ReLU[7].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$3087(.Z({ \dot_product_and_ReLU[7].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$3088(.Z({ \dot_product_and_ReLU[7].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$3089(.Z({ \dot_product_and_ReLU[7].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$3090(.Z({ \dot_product_and_ReLU[7].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$3091(.Z({ \dot_product_and_ReLU[7].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$3092(.Z({ \dot_product_and_ReLU[7].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$3093(.Z({ \dot_product_and_ReLU[7].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$3094(.Z({ \dot_product_and_ReLU[7].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$3095(.Z({ \dot_product_and_ReLU[7].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$3096(.Z({ \dot_product_and_ReLU[7].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$3097(.Z({ \dot_product_and_ReLU[7].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$3098(.Z({ \dot_product_and_ReLU[7].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$3099(.Z({ \dot_product_and_ReLU[7].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$3100(.Z({ \dot_product_and_ReLU[7].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$3101(.Z({ \dot_product_and_ReLU[7].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$3102(.Z({ \dot_product_and_ReLU[7].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$3103(.Z({ \dot_product_and_ReLU[7].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$3104(.Z({ \dot_product_and_ReLU[7].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$3105(.Z({ \dot_product_and_ReLU[7].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$3106(.Z({ \dot_product_and_ReLU[7].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$3107(.Z({ \dot_product_and_ReLU[7].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$3108(.Z({ \dot_product_and_ReLU[7].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$3109(.Z({ \dot_product_and_ReLU[7].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$3110(.Z({ \dot_product_and_ReLU[7].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$3111(.Z({ \dot_product_and_ReLU[7].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$3112(.Z({ \dot_product_and_ReLU[7].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$3113(.Z({ \dot_product_and_ReLU[7].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$3114(.Z({ \dot_product_and_ReLU[7].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$3115(.Z({ \dot_product_and_ReLU[7].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$3116(.Z({ \dot_product_and_ReLU[7].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$3117(.Z({ \dot_product_and_ReLU[7].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$3118(.Z({ \dot_product_and_ReLU[7].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$3119(.Z({ \dot_product_and_ReLU[7].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$3120(.Z({ \dot_product_and_ReLU[7].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$3121(.Z({ \dot_product_and_ReLU[7].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$3122(.Z({ \dot_product_and_ReLU[7].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$3123(.Z({ \dot_product_and_ReLU[7].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$3124(.Z({ \dot_product_and_ReLU[7].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$3125(.Z({ \dot_product_and_ReLU[7].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$3126(.Z({ \dot_product_and_ReLU[7].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$3127(.Z({ \dot_product_and_ReLU[7].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$3128(.Z({ \dot_product_and_ReLU[7].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$3129(.Z({ \dot_product_and_ReLU[7].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$3130(.Z({ \dot_product_and_ReLU[7].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$3131(.Z({ \dot_product_and_ReLU[7].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$3132(.Z({ \dot_product_and_ReLU[7].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$3133(.Z({ \dot_product_and_ReLU[7].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$3134(.Z({ \dot_product_and_ReLU[7].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$3135(.Z({ \dot_product_and_ReLU[7].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$3136(.Z({ \dot_product_and_ReLU[7].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$3137(.Z({ \dot_product_and_ReLU[7].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$3138(.Z({ \dot_product_and_ReLU[7].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$3139(.Z({ \dot_product_and_ReLU[7].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$3140(.Z({ \dot_product_and_ReLU[7].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$3141(.Z({ \dot_product_and_ReLU[7].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$3142(.Z({ \dot_product_and_ReLU[7].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$3143(.Z({ \dot_product_and_ReLU[7].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$3144(.Z({ \dot_product_and_ReLU[7].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$3145(.Z({ \dot_product_and_ReLU[7].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$3146(.Z({ \dot_product_and_ReLU[7].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$3147(.Z({ \dot_product_and_ReLU[7].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$3148(.Z({ \dot_product_and_ReLU[7].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$3149(.Z({ \dot_product_and_ReLU[7].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$3150(.Z({ \dot_product_and_ReLU[7].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$3151(.Z({ \dot_product_and_ReLU[7].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$3152(.Z({ \dot_product_and_ReLU[7].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$3153(.Z({ \dot_product_and_ReLU[7].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$3154(.Z({ \dot_product_and_ReLU[7].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$3155(.Z({ \dot_product_and_ReLU[7].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$3156(.Z({ \dot_product_and_ReLU[7].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$3157(.Z({ \dot_product_and_ReLU[7].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$3158(.Z({ \dot_product_and_ReLU[7].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$3159(.Z({ \dot_product_and_ReLU[7].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$3160(.Z({ \dot_product_and_ReLU[7].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$3161(.Z({ \dot_product_and_ReLU[7].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$3162(.Z({ \dot_product_and_ReLU[7].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$3163(.Z({ \dot_product_and_ReLU[7].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$3164(.Z({ \dot_product_and_ReLU[7].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$3165(.Z({ \dot_product_and_ReLU[7].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$3166(.Z({ \dot_product_and_ReLU[7].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$3167(.Z({ \dot_product_and_ReLU[7].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$3168(.Z({ \dot_product_and_ReLU[7].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$3169(.Z({ \dot_product_and_ReLU[7].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$3170(.Z({ \dot_product_and_ReLU[7].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$3171(.Z({ \dot_product_and_ReLU[7].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$3172(.Z({ \dot_product_and_ReLU[7].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$3173(.Z({ \dot_product_and_ReLU[7].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$3174(.Z({ \dot_product_and_ReLU[7].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$3175(.Z({ \dot_product_and_ReLU[7].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$3176(.Z({ \dot_product_and_ReLU[7].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$3177(.Z({ \dot_product_and_ReLU[7].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$3178(.Z({ \dot_product_and_ReLU[7].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$3179(.Z({ \dot_product_and_ReLU[7].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$3180(.Z({ \dot_product_and_ReLU[7].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$3181(.Z({ \dot_product_and_ReLU[7].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$3182(.Z({ \dot_product_and_ReLU[7].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$3183(.Z({ \dot_product_and_ReLU[7].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$3184(.Z({ \dot_product_and_ReLU[7].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$3185(.Z({ \dot_product_and_ReLU[7].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$3186(.Z({ \dot_product_and_ReLU[7].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$3187(.Z({ \dot_product_and_ReLU[7].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$3188(.Z({ \dot_product_and_ReLU[7].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$3189(.Z({ \dot_product_and_ReLU[7].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$3190(.Z({ \dot_product_and_ReLU[7].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$3191(.Z({ \dot_product_and_ReLU[7].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$3192(.Z({ \dot_product_and_ReLU[7].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$3193(.Z({ \dot_product_and_ReLU[7].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$3194(.Z({ \dot_product_and_ReLU[7].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$3195(.Z({ \dot_product_and_ReLU[7].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$3196(.Z({ \dot_product_and_ReLU[7].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$3197(.Z({ \dot_product_and_ReLU[7].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$3198(.Z({ \dot_product_and_ReLU[7].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$3199(.Z({ \dot_product_and_ReLU[7].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$3200(.Z({ \dot_product_and_ReLU[7].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$3201(.Z({ \dot_product_and_ReLU[7].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$3202(.Z({ \dot_product_and_ReLU[7].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$3203(.Z({ \dot_product_and_ReLU[7].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$3204(.Z({ \dot_product_and_ReLU[7].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$3205(.Z({ \dot_product_and_ReLU[7].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$3206(.Z({ \dot_product_and_ReLU[7].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$3207(.Z({ \dot_product_and_ReLU[7].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$3208(.Z({ \dot_product_and_ReLU[7].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$3209(.Z({ \dot_product_and_ReLU[7].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$3210(.Z({ \dot_product_and_ReLU[7].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$3211(.Z({ \dot_product_and_ReLU[7].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$3212(.Z({ \dot_product_and_ReLU[7].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$3213(.Z({ \dot_product_and_ReLU[7].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$3214(.Z({ \dot_product_and_ReLU[7].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$3215(.Z({ \dot_product_and_ReLU[7].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$3216(.Z({ \dot_product_and_ReLU[7].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$3217(.Z({ \dot_product_and_ReLU[7].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$3218(.Z({ \dot_product_and_ReLU[7].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$3219(.Z({ \dot_product_and_ReLU[7].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$3220(.Z({ \dot_product_and_ReLU[7].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$3221(.Z({ \dot_product_and_ReLU[7].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$3222(.Z({ \dot_product_and_ReLU[7].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$3223(.Z({ \dot_product_and_ReLU[7].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$3224(.Z({ \dot_product_and_ReLU[7].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$3225(.Z({ \dot_product_and_ReLU[7].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$3226(.Z({ \dot_product_and_ReLU[7].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$3227(.Z({ \dot_product_and_ReLU[7].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$3228(.Z({ \dot_product_and_ReLU[7].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$3229(.Z({ \dot_product_and_ReLU[7].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$3230(.Z({ \dot_product_and_ReLU[7].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$3231(.Z({ \dot_product_and_ReLU[7].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$3232(.Z({ \dot_product_and_ReLU[7].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$3233(.Z({ \dot_product_and_ReLU[7].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$3234(.Z({ \dot_product_and_ReLU[7].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$3235(.Z({ \dot_product_and_ReLU[7].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$3236(.Z({ \dot_product_and_ReLU[7].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$3237(.Z({ \dot_product_and_ReLU[7].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$3238(.Z({ \dot_product_and_ReLU[7].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$3239(.Z({ \dot_product_and_ReLU[7].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$3240(.Z({ \dot_product_and_ReLU[7].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$3241(.Z({ \dot_product_and_ReLU[7].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$3242(.Z({ \dot_product_and_ReLU[7].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$3243(.Z({ \dot_product_and_ReLU[7].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$3244(.Z({ \dot_product_and_ReLU[7].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$3245(.Z({ \dot_product_and_ReLU[7].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$3246(.Z({ \dot_product_and_ReLU[7].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$3247(.Z({ \dot_product_and_ReLU[7].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$3248(.Z({ \dot_product_and_ReLU[7].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$3249(.Z({ \dot_product_and_ReLU[7].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$3250(.Z({ \dot_product_and_ReLU[7].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$3251(.Z({ \dot_product_and_ReLU[7].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$3252(.Z({ \dot_product_and_ReLU[7].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$3253(.Z({ \dot_product_and_ReLU[7].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$3254(.Z({ \dot_product_and_ReLU[7].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$3255(.Z({ \dot_product_and_ReLU[7].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$3256(.Z({ \dot_product_and_ReLU[7].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$3257(.Z({ \dot_product_and_ReLU[7].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$3258(.Z({ \dot_product_and_ReLU[7].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$3259(.Z({ \dot_product_and_ReLU[7].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$3260(.Z({ \dot_product_and_ReLU[7].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$3261(.Z({ \dot_product_and_ReLU[7].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$3262(.Z({ \dot_product_and_ReLU[7].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$3263(.Z({ \dot_product_and_ReLU[7].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$3264(.Z({ \dot_product_and_ReLU[7].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$3265(.Z({ \dot_product_and_ReLU[7].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$3266(.Z({ \dot_product_and_ReLU[7].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$3267(.Z({ \dot_product_and_ReLU[7].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$3268(.Z({ \dot_product_and_ReLU[7].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$3269(.Z({ \dot_product_and_ReLU[7].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$3270(.Z({ \dot_product_and_ReLU[7].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$3271(.Z({ \dot_product_and_ReLU[7].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$3272(.Z({ \dot_product_and_ReLU[7].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$3273(.Z({ \dot_product_and_ReLU[7].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$3274(.Z({ \dot_product_and_ReLU[7].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$3275(.Z({ \dot_product_and_ReLU[7].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$3276(.Z({ \dot_product_and_ReLU[7].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$3277(.Z({ \dot_product_and_ReLU[7].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$3278(.Z({ \dot_product_and_ReLU[7].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$3279(.Z({ \dot_product_and_ReLU[7].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$3280(.Z({ \dot_product_and_ReLU[7].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$3281(.Z({ \dot_product_and_ReLU[7].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$3282(.Z({ \dot_product_and_ReLU[7].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$3283(.Z({ \dot_product_and_ReLU[7].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$3284(.Z({ \dot_product_and_ReLU[7].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$3285(.Z({ \dot_product_and_ReLU[7].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$3286(.Z({ \dot_product_and_ReLU[7].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$3287(.Z({ \dot_product_and_ReLU[7].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$3288(.Z({ \dot_product_and_ReLU[7].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$3289(.Z({ \dot_product_and_ReLU[7].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$3290(.Z({ \dot_product_and_ReLU[7].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$3291(.Z({ \dot_product_and_ReLU[7].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$3292(.Z({ \dot_product_and_ReLU[7].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$3293(.Z({ \dot_product_and_ReLU[7].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$3294(.Z({ \dot_product_and_ReLU[7].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$3295(.Z({ \dot_product_and_ReLU[7].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$3296(.Z({ \dot_product_and_ReLU[7].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$3297(.Z({ \dot_product_and_ReLU[7].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$3298(.Z({ \dot_product_and_ReLU[7].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$3299(.Z({ \dot_product_and_ReLU[7].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$3300(.Z({ \dot_product_and_ReLU[7].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$3301(.Z({ \dot_product_and_ReLU[7].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$3302(.Z({ \dot_product_and_ReLU[7].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$3303(.Z({ \dot_product_and_ReLU[7].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$3304(.Z({ \dot_product_and_ReLU[7].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$3305(.Z({ \dot_product_and_ReLU[7].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$3306(.Z({ \dot_product_and_ReLU[7].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$3307(.Z({ \dot_product_and_ReLU[7].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$3308(.Z({ \dot_product_and_ReLU[7].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$3309(.Z({ \dot_product_and_ReLU[7].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$3310(.Z({ \dot_product_and_ReLU[7].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$3311(.Z({ \dot_product_and_ReLU[7].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$3312(.Z({ \dot_product_and_ReLU[7].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$3313(.Z({ \dot_product_and_ReLU[7].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$3314(.Z({ \dot_product_and_ReLU[7].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$3315(.Z({ \dot_product_and_ReLU[7].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$3316(.Z({ \dot_product_and_ReLU[7].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$3317(.Z({ \dot_product_and_ReLU[7].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$3318(.Z({ \dot_product_and_ReLU[7].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$3319(.Z({ \dot_product_and_ReLU[7].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$3320(.Z({ \dot_product_and_ReLU[7].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$3321(.Z({ \dot_product_and_ReLU[7].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$3322(.Z({ \dot_product_and_ReLU[7].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$3323(.Z({ \dot_product_and_ReLU[7].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$3324(.Z({ \dot_product_and_ReLU[7].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$3325(.Z({ \dot_product_and_ReLU[7].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$3326(.Z({ \dot_product_and_ReLU[7].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$3327(.Z({ \dot_product_and_ReLU[7].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$3328(.Z({ \dot_product_and_ReLU[7].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[7][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$3329(.Z({ \dot_product_and_ReLU[6].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$3330(.Z({ \dot_product_and_ReLU[6].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$3331(.Z({ \dot_product_and_ReLU[6].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$3332(.Z({ \dot_product_and_ReLU[6].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$3333(.Z({ \dot_product_and_ReLU[6].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$3334(.Z({ \dot_product_and_ReLU[6].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$3335(.Z({ \dot_product_and_ReLU[6].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$3336(.Z({ \dot_product_and_ReLU[6].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$3337(.Z({ \dot_product_and_ReLU[6].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$3338(.Z({ \dot_product_and_ReLU[6].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$3339(.Z({ \dot_product_and_ReLU[6].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$3340(.Z({ \dot_product_and_ReLU[6].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$3341(.Z({ \dot_product_and_ReLU[6].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$3342(.Z({ \dot_product_and_ReLU[6].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$3343(.Z({ \dot_product_and_ReLU[6].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$3344(.Z({ \dot_product_and_ReLU[6].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$3345(.Z({ \dot_product_and_ReLU[6].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$3346(.Z({ \dot_product_and_ReLU[6].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$3347(.Z({ \dot_product_and_ReLU[6].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$3348(.Z({ \dot_product_and_ReLU[6].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$3349(.Z({ \dot_product_and_ReLU[6].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$3350(.Z({ \dot_product_and_ReLU[6].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$3351(.Z({ \dot_product_and_ReLU[6].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$3352(.Z({ \dot_product_and_ReLU[6].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$3353(.Z({ \dot_product_and_ReLU[6].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$3354(.Z({ \dot_product_and_ReLU[6].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$3355(.Z({ \dot_product_and_ReLU[6].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$3356(.Z({ \dot_product_and_ReLU[6].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$3357(.Z({ \dot_product_and_ReLU[6].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$3358(.Z({ \dot_product_and_ReLU[6].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$3359(.Z({ \dot_product_and_ReLU[6].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$3360(.Z({ \dot_product_and_ReLU[6].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$3361(.Z({ \dot_product_and_ReLU[6].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$3362(.Z({ \dot_product_and_ReLU[6].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$3363(.Z({ \dot_product_and_ReLU[6].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$3364(.Z({ \dot_product_and_ReLU[6].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$3365(.Z({ \dot_product_and_ReLU[6].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$3366(.Z({ \dot_product_and_ReLU[6].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$3367(.Z({ \dot_product_and_ReLU[6].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$3368(.Z({ \dot_product_and_ReLU[6].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$3369(.Z({ \dot_product_and_ReLU[6].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$3370(.Z({ \dot_product_and_ReLU[6].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$3371(.Z({ \dot_product_and_ReLU[6].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$3372(.Z({ \dot_product_and_ReLU[6].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$3373(.Z({ \dot_product_and_ReLU[6].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$3374(.Z({ \dot_product_and_ReLU[6].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$3375(.Z({ \dot_product_and_ReLU[6].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$3376(.Z({ \dot_product_and_ReLU[6].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$3377(.Z({ \dot_product_and_ReLU[6].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$3378(.Z({ \dot_product_and_ReLU[6].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$3379(.Z({ \dot_product_and_ReLU[6].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$3380(.Z({ \dot_product_and_ReLU[6].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$3381(.Z({ \dot_product_and_ReLU[6].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$3382(.Z({ \dot_product_and_ReLU[6].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$3383(.Z({ \dot_product_and_ReLU[6].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$3384(.Z({ \dot_product_and_ReLU[6].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$3385(.Z({ \dot_product_and_ReLU[6].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$3386(.Z({ \dot_product_and_ReLU[6].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$3387(.Z({ \dot_product_and_ReLU[6].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$3388(.Z({ \dot_product_and_ReLU[6].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$3389(.Z({ \dot_product_and_ReLU[6].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$3390(.Z({ \dot_product_and_ReLU[6].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$3391(.Z({ \dot_product_and_ReLU[6].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$3392(.Z({ \dot_product_and_ReLU[6].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$3393(.Z({ \dot_product_and_ReLU[6].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$3394(.Z({ \dot_product_and_ReLU[6].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$3395(.Z({ \dot_product_and_ReLU[6].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$3396(.Z({ \dot_product_and_ReLU[6].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$3397(.Z({ \dot_product_and_ReLU[6].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$3398(.Z({ \dot_product_and_ReLU[6].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$3399(.Z({ \dot_product_and_ReLU[6].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$3400(.Z({ \dot_product_and_ReLU[6].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$3401(.Z({ \dot_product_and_ReLU[6].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$3402(.Z({ \dot_product_and_ReLU[6].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$3403(.Z({ \dot_product_and_ReLU[6].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$3404(.Z({ \dot_product_and_ReLU[6].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$3405(.Z({ \dot_product_and_ReLU[6].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$3406(.Z({ \dot_product_and_ReLU[6].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$3407(.Z({ \dot_product_and_ReLU[6].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$3408(.Z({ \dot_product_and_ReLU[6].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$3409(.Z({ \dot_product_and_ReLU[6].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$3410(.Z({ \dot_product_and_ReLU[6].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$3411(.Z({ \dot_product_and_ReLU[6].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$3412(.Z({ \dot_product_and_ReLU[6].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$3413(.Z({ \dot_product_and_ReLU[6].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$3414(.Z({ \dot_product_and_ReLU[6].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$3415(.Z({ \dot_product_and_ReLU[6].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$3416(.Z({ \dot_product_and_ReLU[6].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$3417(.Z({ \dot_product_and_ReLU[6].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$3418(.Z({ \dot_product_and_ReLU[6].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$3419(.Z({ \dot_product_and_ReLU[6].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$3420(.Z({ \dot_product_and_ReLU[6].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$3421(.Z({ \dot_product_and_ReLU[6].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$3422(.Z({ \dot_product_and_ReLU[6].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$3423(.Z({ \dot_product_and_ReLU[6].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$3424(.Z({ \dot_product_and_ReLU[6].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$3425(.Z({ \dot_product_and_ReLU[6].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$3426(.Z({ \dot_product_and_ReLU[6].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$3427(.Z({ \dot_product_and_ReLU[6].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$3428(.Z({ \dot_product_and_ReLU[6].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$3429(.Z({ \dot_product_and_ReLU[6].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$3430(.Z({ \dot_product_and_ReLU[6].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$3431(.Z({ \dot_product_and_ReLU[6].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$3432(.Z({ \dot_product_and_ReLU[6].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$3433(.Z({ \dot_product_and_ReLU[6].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$3434(.Z({ \dot_product_and_ReLU[6].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$3435(.Z({ \dot_product_and_ReLU[6].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$3436(.Z({ \dot_product_and_ReLU[6].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$3437(.Z({ \dot_product_and_ReLU[6].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$3438(.Z({ \dot_product_and_ReLU[6].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$3439(.Z({ \dot_product_and_ReLU[6].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$3440(.Z({ \dot_product_and_ReLU[6].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$3441(.Z({ \dot_product_and_ReLU[6].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$3442(.Z({ \dot_product_and_ReLU[6].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$3443(.Z({ \dot_product_and_ReLU[6].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$3444(.Z({ \dot_product_and_ReLU[6].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$3445(.Z({ \dot_product_and_ReLU[6].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$3446(.Z({ \dot_product_and_ReLU[6].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$3447(.Z({ \dot_product_and_ReLU[6].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$3448(.Z({ \dot_product_and_ReLU[6].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$3449(.Z({ \dot_product_and_ReLU[6].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$3450(.Z({ \dot_product_and_ReLU[6].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$3451(.Z({ \dot_product_and_ReLU[6].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$3452(.Z({ \dot_product_and_ReLU[6].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$3453(.Z({ \dot_product_and_ReLU[6].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$3454(.Z({ \dot_product_and_ReLU[6].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$3455(.Z({ \dot_product_and_ReLU[6].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$3456(.Z({ \dot_product_and_ReLU[6].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$3457(.Z({ \dot_product_and_ReLU[6].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$3458(.Z({ \dot_product_and_ReLU[6].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$3459(.Z({ \dot_product_and_ReLU[6].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$3460(.Z({ \dot_product_and_ReLU[6].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$3461(.Z({ \dot_product_and_ReLU[6].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$3462(.Z({ \dot_product_and_ReLU[6].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$3463(.Z({ \dot_product_and_ReLU[6].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$3464(.Z({ \dot_product_and_ReLU[6].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$3465(.Z({ \dot_product_and_ReLU[6].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$3466(.Z({ \dot_product_and_ReLU[6].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$3467(.Z({ \dot_product_and_ReLU[6].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$3468(.Z({ \dot_product_and_ReLU[6].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$3469(.Z({ \dot_product_and_ReLU[6].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$3470(.Z({ \dot_product_and_ReLU[6].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$3471(.Z({ \dot_product_and_ReLU[6].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$3472(.Z({ \dot_product_and_ReLU[6].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$3473(.Z({ \dot_product_and_ReLU[6].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$3474(.Z({ \dot_product_and_ReLU[6].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$3475(.Z({ \dot_product_and_ReLU[6].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$3476(.Z({ \dot_product_and_ReLU[6].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$3477(.Z({ \dot_product_and_ReLU[6].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$3478(.Z({ \dot_product_and_ReLU[6].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$3479(.Z({ \dot_product_and_ReLU[6].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$3480(.Z({ \dot_product_and_ReLU[6].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$3481(.Z({ \dot_product_and_ReLU[6].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$3482(.Z({ \dot_product_and_ReLU[6].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$3483(.Z({ \dot_product_and_ReLU[6].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$3484(.Z({ \dot_product_and_ReLU[6].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$3485(.Z({ \dot_product_and_ReLU[6].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$3486(.Z({ \dot_product_and_ReLU[6].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$3487(.Z({ \dot_product_and_ReLU[6].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$3488(.Z({ \dot_product_and_ReLU[6].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$3489(.Z({ \dot_product_and_ReLU[6].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$3490(.Z({ \dot_product_and_ReLU[6].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$3491(.Z({ \dot_product_and_ReLU[6].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$3492(.Z({ \dot_product_and_ReLU[6].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$3493(.Z({ \dot_product_and_ReLU[6].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$3494(.Z({ \dot_product_and_ReLU[6].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$3495(.Z({ \dot_product_and_ReLU[6].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$3496(.Z({ \dot_product_and_ReLU[6].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$3497(.Z({ \dot_product_and_ReLU[6].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$3498(.Z({ \dot_product_and_ReLU[6].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$3499(.Z({ \dot_product_and_ReLU[6].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$3500(.Z({ \dot_product_and_ReLU[6].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$3501(.Z({ \dot_product_and_ReLU[6].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$3502(.Z({ \dot_product_and_ReLU[6].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$3503(.Z({ \dot_product_and_ReLU[6].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$3504(.Z({ \dot_product_and_ReLU[6].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$3505(.Z({ \dot_product_and_ReLU[6].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$3506(.Z({ \dot_product_and_ReLU[6].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$3507(.Z({ \dot_product_and_ReLU[6].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$3508(.Z({ \dot_product_and_ReLU[6].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$3509(.Z({ \dot_product_and_ReLU[6].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$3510(.Z({ \dot_product_and_ReLU[6].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$3511(.Z({ \dot_product_and_ReLU[6].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$3512(.Z({ \dot_product_and_ReLU[6].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$3513(.Z({ \dot_product_and_ReLU[6].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$3514(.Z({ \dot_product_and_ReLU[6].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$3515(.Z({ \dot_product_and_ReLU[6].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$3516(.Z({ \dot_product_and_ReLU[6].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$3517(.Z({ \dot_product_and_ReLU[6].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$3518(.Z({ \dot_product_and_ReLU[6].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$3519(.Z({ \dot_product_and_ReLU[6].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$3520(.Z({ \dot_product_and_ReLU[6].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$3521(.Z({ \dot_product_and_ReLU[6].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$3522(.Z({ \dot_product_and_ReLU[6].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$3523(.Z({ \dot_product_and_ReLU[6].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$3524(.Z({ \dot_product_and_ReLU[6].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$3525(.Z({ \dot_product_and_ReLU[6].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$3526(.Z({ \dot_product_and_ReLU[6].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$3527(.Z({ \dot_product_and_ReLU[6].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$3528(.Z({ \dot_product_and_ReLU[6].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$3529(.Z({ \dot_product_and_ReLU[6].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$3530(.Z({ \dot_product_and_ReLU[6].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$3531(.Z({ \dot_product_and_ReLU[6].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$3532(.Z({ \dot_product_and_ReLU[6].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$3533(.Z({ \dot_product_and_ReLU[6].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$3534(.Z({ \dot_product_and_ReLU[6].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$3535(.Z({ \dot_product_and_ReLU[6].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$3536(.Z({ \dot_product_and_ReLU[6].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$3537(.Z({ \dot_product_and_ReLU[6].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$3538(.Z({ \dot_product_and_ReLU[6].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$3539(.Z({ \dot_product_and_ReLU[6].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$3540(.Z({ \dot_product_and_ReLU[6].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$3541(.Z({ \dot_product_and_ReLU[6].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$3542(.Z({ \dot_product_and_ReLU[6].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$3543(.Z({ \dot_product_and_ReLU[6].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$3544(.Z({ \dot_product_and_ReLU[6].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$3545(.Z({ \dot_product_and_ReLU[6].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$3546(.Z({ \dot_product_and_ReLU[6].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$3547(.Z({ \dot_product_and_ReLU[6].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$3548(.Z({ \dot_product_and_ReLU[6].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$3549(.Z({ \dot_product_and_ReLU[6].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$3550(.Z({ \dot_product_and_ReLU[6].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$3551(.Z({ \dot_product_and_ReLU[6].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$3552(.Z({ \dot_product_and_ReLU[6].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$3553(.Z({ \dot_product_and_ReLU[6].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$3554(.Z({ \dot_product_and_ReLU[6].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$3555(.Z({ \dot_product_and_ReLU[6].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$3556(.Z({ \dot_product_and_ReLU[6].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$3557(.Z({ \dot_product_and_ReLU[6].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$3558(.Z({ \dot_product_and_ReLU[6].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$3559(.Z({ \dot_product_and_ReLU[6].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$3560(.Z({ \dot_product_and_ReLU[6].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$3561(.Z({ \dot_product_and_ReLU[6].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$3562(.Z({ \dot_product_and_ReLU[6].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$3563(.Z({ \dot_product_and_ReLU[6].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$3564(.Z({ \dot_product_and_ReLU[6].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$3565(.Z({ \dot_product_and_ReLU[6].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$3566(.Z({ \dot_product_and_ReLU[6].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$3567(.Z({ \dot_product_and_ReLU[6].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$3568(.Z({ \dot_product_and_ReLU[6].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$3569(.Z({ \dot_product_and_ReLU[6].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$3570(.Z({ \dot_product_and_ReLU[6].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$3571(.Z({ \dot_product_and_ReLU[6].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$3572(.Z({ \dot_product_and_ReLU[6].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$3573(.Z({ \dot_product_and_ReLU[6].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$3574(.Z({ \dot_product_and_ReLU[6].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$3575(.Z({ \dot_product_and_ReLU[6].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$3576(.Z({ \dot_product_and_ReLU[6].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$3577(.Z({ \dot_product_and_ReLU[6].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$3578(.Z({ \dot_product_and_ReLU[6].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$3579(.Z({ \dot_product_and_ReLU[6].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$3580(.Z({ \dot_product_and_ReLU[6].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$3581(.Z({ \dot_product_and_ReLU[6].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$3582(.Z({ \dot_product_and_ReLU[6].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$3583(.Z({ \dot_product_and_ReLU[6].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$3584(.Z({ \dot_product_and_ReLU[6].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[6][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$3585(.Z({ \dot_product_and_ReLU[5].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$3586(.Z({ \dot_product_and_ReLU[5].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$3587(.Z({ \dot_product_and_ReLU[5].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$3588(.Z({ \dot_product_and_ReLU[5].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$3589(.Z({ \dot_product_and_ReLU[5].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$3590(.Z({ \dot_product_and_ReLU[5].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$3591(.Z({ \dot_product_and_ReLU[5].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$3592(.Z({ \dot_product_and_ReLU[5].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$3593(.Z({ \dot_product_and_ReLU[5].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$3594(.Z({ \dot_product_and_ReLU[5].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$3595(.Z({ \dot_product_and_ReLU[5].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$3596(.Z({ \dot_product_and_ReLU[5].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$3597(.Z({ \dot_product_and_ReLU[5].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$3598(.Z({ \dot_product_and_ReLU[5].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$3599(.Z({ \dot_product_and_ReLU[5].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$3600(.Z({ \dot_product_and_ReLU[5].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$3601(.Z({ \dot_product_and_ReLU[5].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$3602(.Z({ \dot_product_and_ReLU[5].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$3603(.Z({ \dot_product_and_ReLU[5].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$3604(.Z({ \dot_product_and_ReLU[5].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$3605(.Z({ \dot_product_and_ReLU[5].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$3606(.Z({ \dot_product_and_ReLU[5].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$3607(.Z({ \dot_product_and_ReLU[5].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$3608(.Z({ \dot_product_and_ReLU[5].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$3609(.Z({ \dot_product_and_ReLU[5].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$3610(.Z({ \dot_product_and_ReLU[5].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$3611(.Z({ \dot_product_and_ReLU[5].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$3612(.Z({ \dot_product_and_ReLU[5].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$3613(.Z({ \dot_product_and_ReLU[5].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$3614(.Z({ \dot_product_and_ReLU[5].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$3615(.Z({ \dot_product_and_ReLU[5].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$3616(.Z({ \dot_product_and_ReLU[5].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$3617(.Z({ \dot_product_and_ReLU[5].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$3618(.Z({ \dot_product_and_ReLU[5].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$3619(.Z({ \dot_product_and_ReLU[5].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$3620(.Z({ \dot_product_and_ReLU[5].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$3621(.Z({ \dot_product_and_ReLU[5].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$3622(.Z({ \dot_product_and_ReLU[5].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$3623(.Z({ \dot_product_and_ReLU[5].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$3624(.Z({ \dot_product_and_ReLU[5].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$3625(.Z({ \dot_product_and_ReLU[5].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$3626(.Z({ \dot_product_and_ReLU[5].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$3627(.Z({ \dot_product_and_ReLU[5].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$3628(.Z({ \dot_product_and_ReLU[5].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$3629(.Z({ \dot_product_and_ReLU[5].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$3630(.Z({ \dot_product_and_ReLU[5].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$3631(.Z({ \dot_product_and_ReLU[5].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$3632(.Z({ \dot_product_and_ReLU[5].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$3633(.Z({ \dot_product_and_ReLU[5].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$3634(.Z({ \dot_product_and_ReLU[5].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$3635(.Z({ \dot_product_and_ReLU[5].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$3636(.Z({ \dot_product_and_ReLU[5].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$3637(.Z({ \dot_product_and_ReLU[5].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$3638(.Z({ \dot_product_and_ReLU[5].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$3639(.Z({ \dot_product_and_ReLU[5].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$3640(.Z({ \dot_product_and_ReLU[5].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$3641(.Z({ \dot_product_and_ReLU[5].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$3642(.Z({ \dot_product_and_ReLU[5].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$3643(.Z({ \dot_product_and_ReLU[5].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$3644(.Z({ \dot_product_and_ReLU[5].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$3645(.Z({ \dot_product_and_ReLU[5].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$3646(.Z({ \dot_product_and_ReLU[5].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$3647(.Z({ \dot_product_and_ReLU[5].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$3648(.Z({ \dot_product_and_ReLU[5].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$3649(.Z({ \dot_product_and_ReLU[5].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$3650(.Z({ \dot_product_and_ReLU[5].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$3651(.Z({ \dot_product_and_ReLU[5].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$3652(.Z({ \dot_product_and_ReLU[5].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$3653(.Z({ \dot_product_and_ReLU[5].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$3654(.Z({ \dot_product_and_ReLU[5].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$3655(.Z({ \dot_product_and_ReLU[5].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$3656(.Z({ \dot_product_and_ReLU[5].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$3657(.Z({ \dot_product_and_ReLU[5].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$3658(.Z({ \dot_product_and_ReLU[5].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$3659(.Z({ \dot_product_and_ReLU[5].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$3660(.Z({ \dot_product_and_ReLU[5].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$3661(.Z({ \dot_product_and_ReLU[5].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$3662(.Z({ \dot_product_and_ReLU[5].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$3663(.Z({ \dot_product_and_ReLU[5].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$3664(.Z({ \dot_product_and_ReLU[5].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$3665(.Z({ \dot_product_and_ReLU[5].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$3666(.Z({ \dot_product_and_ReLU[5].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$3667(.Z({ \dot_product_and_ReLU[5].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$3668(.Z({ \dot_product_and_ReLU[5].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$3669(.Z({ \dot_product_and_ReLU[5].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$3670(.Z({ \dot_product_and_ReLU[5].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$3671(.Z({ \dot_product_and_ReLU[5].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$3672(.Z({ \dot_product_and_ReLU[5].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$3673(.Z({ \dot_product_and_ReLU[5].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$3674(.Z({ \dot_product_and_ReLU[5].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$3675(.Z({ \dot_product_and_ReLU[5].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$3676(.Z({ \dot_product_and_ReLU[5].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$3677(.Z({ \dot_product_and_ReLU[5].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$3678(.Z({ \dot_product_and_ReLU[5].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$3679(.Z({ \dot_product_and_ReLU[5].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$3680(.Z({ \dot_product_and_ReLU[5].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$3681(.Z({ \dot_product_and_ReLU[5].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$3682(.Z({ \dot_product_and_ReLU[5].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$3683(.Z({ \dot_product_and_ReLU[5].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$3684(.Z({ \dot_product_and_ReLU[5].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$3685(.Z({ \dot_product_and_ReLU[5].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$3686(.Z({ \dot_product_and_ReLU[5].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$3687(.Z({ \dot_product_and_ReLU[5].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$3688(.Z({ \dot_product_and_ReLU[5].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$3689(.Z({ \dot_product_and_ReLU[5].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$3690(.Z({ \dot_product_and_ReLU[5].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$3691(.Z({ \dot_product_and_ReLU[5].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$3692(.Z({ \dot_product_and_ReLU[5].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$3693(.Z({ \dot_product_and_ReLU[5].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$3694(.Z({ \dot_product_and_ReLU[5].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$3695(.Z({ \dot_product_and_ReLU[5].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$3696(.Z({ \dot_product_and_ReLU[5].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$3697(.Z({ \dot_product_and_ReLU[5].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$3698(.Z({ \dot_product_and_ReLU[5].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$3699(.Z({ \dot_product_and_ReLU[5].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$3700(.Z({ \dot_product_and_ReLU[5].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$3701(.Z({ \dot_product_and_ReLU[5].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$3702(.Z({ \dot_product_and_ReLU[5].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$3703(.Z({ \dot_product_and_ReLU[5].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$3704(.Z({ \dot_product_and_ReLU[5].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$3705(.Z({ \dot_product_and_ReLU[5].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$3706(.Z({ \dot_product_and_ReLU[5].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$3707(.Z({ \dot_product_and_ReLU[5].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$3708(.Z({ \dot_product_and_ReLU[5].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$3709(.Z({ \dot_product_and_ReLU[5].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$3710(.Z({ \dot_product_and_ReLU[5].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$3711(.Z({ \dot_product_and_ReLU[5].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$3712(.Z({ \dot_product_and_ReLU[5].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$3713(.Z({ \dot_product_and_ReLU[5].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$3714(.Z({ \dot_product_and_ReLU[5].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$3715(.Z({ \dot_product_and_ReLU[5].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$3716(.Z({ \dot_product_and_ReLU[5].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$3717(.Z({ \dot_product_and_ReLU[5].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$3718(.Z({ \dot_product_and_ReLU[5].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$3719(.Z({ \dot_product_and_ReLU[5].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$3720(.Z({ \dot_product_and_ReLU[5].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$3721(.Z({ \dot_product_and_ReLU[5].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$3722(.Z({ \dot_product_and_ReLU[5].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$3723(.Z({ \dot_product_and_ReLU[5].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$3724(.Z({ \dot_product_and_ReLU[5].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$3725(.Z({ \dot_product_and_ReLU[5].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$3726(.Z({ \dot_product_and_ReLU[5].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$3727(.Z({ \dot_product_and_ReLU[5].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$3728(.Z({ \dot_product_and_ReLU[5].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$3729(.Z({ \dot_product_and_ReLU[5].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$3730(.Z({ \dot_product_and_ReLU[5].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$3731(.Z({ \dot_product_and_ReLU[5].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$3732(.Z({ \dot_product_and_ReLU[5].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$3733(.Z({ \dot_product_and_ReLU[5].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$3734(.Z({ \dot_product_and_ReLU[5].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$3735(.Z({ \dot_product_and_ReLU[5].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$3736(.Z({ \dot_product_and_ReLU[5].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$3737(.Z({ \dot_product_and_ReLU[5].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$3738(.Z({ \dot_product_and_ReLU[5].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$3739(.Z({ \dot_product_and_ReLU[5].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$3740(.Z({ \dot_product_and_ReLU[5].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$3741(.Z({ \dot_product_and_ReLU[5].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$3742(.Z({ \dot_product_and_ReLU[5].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$3743(.Z({ \dot_product_and_ReLU[5].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$3744(.Z({ \dot_product_and_ReLU[5].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$3745(.Z({ \dot_product_and_ReLU[5].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$3746(.Z({ \dot_product_and_ReLU[5].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$3747(.Z({ \dot_product_and_ReLU[5].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$3748(.Z({ \dot_product_and_ReLU[5].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$3749(.Z({ \dot_product_and_ReLU[5].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$3750(.Z({ \dot_product_and_ReLU[5].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$3751(.Z({ \dot_product_and_ReLU[5].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$3752(.Z({ \dot_product_and_ReLU[5].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$3753(.Z({ \dot_product_and_ReLU[5].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$3754(.Z({ \dot_product_and_ReLU[5].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$3755(.Z({ \dot_product_and_ReLU[5].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$3756(.Z({ \dot_product_and_ReLU[5].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$3757(.Z({ \dot_product_and_ReLU[5].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$3758(.Z({ \dot_product_and_ReLU[5].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$3759(.Z({ \dot_product_and_ReLU[5].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$3760(.Z({ \dot_product_and_ReLU[5].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$3761(.Z({ \dot_product_and_ReLU[5].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$3762(.Z({ \dot_product_and_ReLU[5].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$3763(.Z({ \dot_product_and_ReLU[5].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$3764(.Z({ \dot_product_and_ReLU[5].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$3765(.Z({ \dot_product_and_ReLU[5].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$3766(.Z({ \dot_product_and_ReLU[5].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$3767(.Z({ \dot_product_and_ReLU[5].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$3768(.Z({ \dot_product_and_ReLU[5].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$3769(.Z({ \dot_product_and_ReLU[5].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$3770(.Z({ \dot_product_and_ReLU[5].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$3771(.Z({ \dot_product_and_ReLU[5].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$3772(.Z({ \dot_product_and_ReLU[5].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$3773(.Z({ \dot_product_and_ReLU[5].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$3774(.Z({ \dot_product_and_ReLU[5].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$3775(.Z({ \dot_product_and_ReLU[5].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$3776(.Z({ \dot_product_and_ReLU[5].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$3777(.Z({ \dot_product_and_ReLU[5].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$3778(.Z({ \dot_product_and_ReLU[5].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$3779(.Z({ \dot_product_and_ReLU[5].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$3780(.Z({ \dot_product_and_ReLU[5].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$3781(.Z({ \dot_product_and_ReLU[5].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$3782(.Z({ \dot_product_and_ReLU[5].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$3783(.Z({ \dot_product_and_ReLU[5].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$3784(.Z({ \dot_product_and_ReLU[5].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$3785(.Z({ \dot_product_and_ReLU[5].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$3786(.Z({ \dot_product_and_ReLU[5].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$3787(.Z({ \dot_product_and_ReLU[5].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$3788(.Z({ \dot_product_and_ReLU[5].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$3789(.Z({ \dot_product_and_ReLU[5].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$3790(.Z({ \dot_product_and_ReLU[5].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$3791(.Z({ \dot_product_and_ReLU[5].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$3792(.Z({ \dot_product_and_ReLU[5].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$3793(.Z({ \dot_product_and_ReLU[5].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$3794(.Z({ \dot_product_and_ReLU[5].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$3795(.Z({ \dot_product_and_ReLU[5].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$3796(.Z({ \dot_product_and_ReLU[5].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$3797(.Z({ \dot_product_and_ReLU[5].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$3798(.Z({ \dot_product_and_ReLU[5].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$3799(.Z({ \dot_product_and_ReLU[5].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$3800(.Z({ \dot_product_and_ReLU[5].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$3801(.Z({ \dot_product_and_ReLU[5].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$3802(.Z({ \dot_product_and_ReLU[5].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$3803(.Z({ \dot_product_and_ReLU[5].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$3804(.Z({ \dot_product_and_ReLU[5].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$3805(.Z({ \dot_product_and_ReLU[5].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$3806(.Z({ \dot_product_and_ReLU[5].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$3807(.Z({ \dot_product_and_ReLU[5].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$3808(.Z({ \dot_product_and_ReLU[5].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$3809(.Z({ \dot_product_and_ReLU[5].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$3810(.Z({ \dot_product_and_ReLU[5].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$3811(.Z({ \dot_product_and_ReLU[5].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$3812(.Z({ \dot_product_and_ReLU[5].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$3813(.Z({ \dot_product_and_ReLU[5].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$3814(.Z({ \dot_product_and_ReLU[5].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$3815(.Z({ \dot_product_and_ReLU[5].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$3816(.Z({ \dot_product_and_ReLU[5].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$3817(.Z({ \dot_product_and_ReLU[5].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$3818(.Z({ \dot_product_and_ReLU[5].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$3819(.Z({ \dot_product_and_ReLU[5].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$3820(.Z({ \dot_product_and_ReLU[5].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$3821(.Z({ \dot_product_and_ReLU[5].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$3822(.Z({ \dot_product_and_ReLU[5].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$3823(.Z({ \dot_product_and_ReLU[5].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$3824(.Z({ \dot_product_and_ReLU[5].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$3825(.Z({ \dot_product_and_ReLU[5].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$3826(.Z({ \dot_product_and_ReLU[5].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$3827(.Z({ \dot_product_and_ReLU[5].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$3828(.Z({ \dot_product_and_ReLU[5].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$3829(.Z({ \dot_product_and_ReLU[5].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$3830(.Z({ \dot_product_and_ReLU[5].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$3831(.Z({ \dot_product_and_ReLU[5].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$3832(.Z({ \dot_product_and_ReLU[5].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$3833(.Z({ \dot_product_and_ReLU[5].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$3834(.Z({ \dot_product_and_ReLU[5].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$3835(.Z({ \dot_product_and_ReLU[5].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$3836(.Z({ \dot_product_and_ReLU[5].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$3837(.Z({ \dot_product_and_ReLU[5].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$3838(.Z({ \dot_product_and_ReLU[5].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$3839(.Z({ \dot_product_and_ReLU[5].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$3840(.Z({ \dot_product_and_ReLU[5].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[5][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$3841(.Z({ \dot_product_and_ReLU[4].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$3842(.Z({ \dot_product_and_ReLU[4].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$3843(.Z({ \dot_product_and_ReLU[4].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$3844(.Z({ \dot_product_and_ReLU[4].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$3845(.Z({ \dot_product_and_ReLU[4].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$3846(.Z({ \dot_product_and_ReLU[4].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$3847(.Z({ \dot_product_and_ReLU[4].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$3848(.Z({ \dot_product_and_ReLU[4].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$3849(.Z({ \dot_product_and_ReLU[4].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$3850(.Z({ \dot_product_and_ReLU[4].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$3851(.Z({ \dot_product_and_ReLU[4].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$3852(.Z({ \dot_product_and_ReLU[4].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$3853(.Z({ \dot_product_and_ReLU[4].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$3854(.Z({ \dot_product_and_ReLU[4].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$3855(.Z({ \dot_product_and_ReLU[4].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$3856(.Z({ \dot_product_and_ReLU[4].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$3857(.Z({ \dot_product_and_ReLU[4].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$3858(.Z({ \dot_product_and_ReLU[4].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$3859(.Z({ \dot_product_and_ReLU[4].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$3860(.Z({ \dot_product_and_ReLU[4].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$3861(.Z({ \dot_product_and_ReLU[4].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$3862(.Z({ \dot_product_and_ReLU[4].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$3863(.Z({ \dot_product_and_ReLU[4].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$3864(.Z({ \dot_product_and_ReLU[4].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$3865(.Z({ \dot_product_and_ReLU[4].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$3866(.Z({ \dot_product_and_ReLU[4].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$3867(.Z({ \dot_product_and_ReLU[4].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$3868(.Z({ \dot_product_and_ReLU[4].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$3869(.Z({ \dot_product_and_ReLU[4].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$3870(.Z({ \dot_product_and_ReLU[4].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$3871(.Z({ \dot_product_and_ReLU[4].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$3872(.Z({ \dot_product_and_ReLU[4].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$3873(.Z({ \dot_product_and_ReLU[4].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$3874(.Z({ \dot_product_and_ReLU[4].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$3875(.Z({ \dot_product_and_ReLU[4].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$3876(.Z({ \dot_product_and_ReLU[4].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$3877(.Z({ \dot_product_and_ReLU[4].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$3878(.Z({ \dot_product_and_ReLU[4].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$3879(.Z({ \dot_product_and_ReLU[4].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$3880(.Z({ \dot_product_and_ReLU[4].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$3881(.Z({ \dot_product_and_ReLU[4].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$3882(.Z({ \dot_product_and_ReLU[4].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$3883(.Z({ \dot_product_and_ReLU[4].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$3884(.Z({ \dot_product_and_ReLU[4].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$3885(.Z({ \dot_product_and_ReLU[4].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$3886(.Z({ \dot_product_and_ReLU[4].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$3887(.Z({ \dot_product_and_ReLU[4].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$3888(.Z({ \dot_product_and_ReLU[4].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$3889(.Z({ \dot_product_and_ReLU[4].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$3890(.Z({ \dot_product_and_ReLU[4].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$3891(.Z({ \dot_product_and_ReLU[4].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$3892(.Z({ \dot_product_and_ReLU[4].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$3893(.Z({ \dot_product_and_ReLU[4].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$3894(.Z({ \dot_product_and_ReLU[4].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$3895(.Z({ \dot_product_and_ReLU[4].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$3896(.Z({ \dot_product_and_ReLU[4].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$3897(.Z({ \dot_product_and_ReLU[4].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$3898(.Z({ \dot_product_and_ReLU[4].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$3899(.Z({ \dot_product_and_ReLU[4].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$3900(.Z({ \dot_product_and_ReLU[4].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$3901(.Z({ \dot_product_and_ReLU[4].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$3902(.Z({ \dot_product_and_ReLU[4].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$3903(.Z({ \dot_product_and_ReLU[4].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$3904(.Z({ \dot_product_and_ReLU[4].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$3905(.Z({ \dot_product_and_ReLU[4].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$3906(.Z({ \dot_product_and_ReLU[4].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$3907(.Z({ \dot_product_and_ReLU[4].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$3908(.Z({ \dot_product_and_ReLU[4].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$3909(.Z({ \dot_product_and_ReLU[4].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$3910(.Z({ \dot_product_and_ReLU[4].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$3911(.Z({ \dot_product_and_ReLU[4].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$3912(.Z({ \dot_product_and_ReLU[4].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$3913(.Z({ \dot_product_and_ReLU[4].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$3914(.Z({ \dot_product_and_ReLU[4].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$3915(.Z({ \dot_product_and_ReLU[4].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$3916(.Z({ \dot_product_and_ReLU[4].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$3917(.Z({ \dot_product_and_ReLU[4].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$3918(.Z({ \dot_product_and_ReLU[4].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$3919(.Z({ \dot_product_and_ReLU[4].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$3920(.Z({ \dot_product_and_ReLU[4].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$3921(.Z({ \dot_product_and_ReLU[4].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$3922(.Z({ \dot_product_and_ReLU[4].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$3923(.Z({ \dot_product_and_ReLU[4].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$3924(.Z({ \dot_product_and_ReLU[4].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$3925(.Z({ \dot_product_and_ReLU[4].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$3926(.Z({ \dot_product_and_ReLU[4].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$3927(.Z({ \dot_product_and_ReLU[4].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$3928(.Z({ \dot_product_and_ReLU[4].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$3929(.Z({ \dot_product_and_ReLU[4].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$3930(.Z({ \dot_product_and_ReLU[4].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$3931(.Z({ \dot_product_and_ReLU[4].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$3932(.Z({ \dot_product_and_ReLU[4].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$3933(.Z({ \dot_product_and_ReLU[4].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$3934(.Z({ \dot_product_and_ReLU[4].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$3935(.Z({ \dot_product_and_ReLU[4].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$3936(.Z({ \dot_product_and_ReLU[4].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$3937(.Z({ \dot_product_and_ReLU[4].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$3938(.Z({ \dot_product_and_ReLU[4].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$3939(.Z({ \dot_product_and_ReLU[4].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$3940(.Z({ \dot_product_and_ReLU[4].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$3941(.Z({ \dot_product_and_ReLU[4].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$3942(.Z({ \dot_product_and_ReLU[4].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$3943(.Z({ \dot_product_and_ReLU[4].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$3944(.Z({ \dot_product_and_ReLU[4].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$3945(.Z({ \dot_product_and_ReLU[4].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$3946(.Z({ \dot_product_and_ReLU[4].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$3947(.Z({ \dot_product_and_ReLU[4].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$3948(.Z({ \dot_product_and_ReLU[4].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$3949(.Z({ \dot_product_and_ReLU[4].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$3950(.Z({ \dot_product_and_ReLU[4].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$3951(.Z({ \dot_product_and_ReLU[4].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$3952(.Z({ \dot_product_and_ReLU[4].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$3953(.Z({ \dot_product_and_ReLU[4].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$3954(.Z({ \dot_product_and_ReLU[4].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$3955(.Z({ \dot_product_and_ReLU[4].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$3956(.Z({ \dot_product_and_ReLU[4].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$3957(.Z({ \dot_product_and_ReLU[4].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$3958(.Z({ \dot_product_and_ReLU[4].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$3959(.Z({ \dot_product_and_ReLU[4].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$3960(.Z({ \dot_product_and_ReLU[4].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$3961(.Z({ \dot_product_and_ReLU[4].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$3962(.Z({ \dot_product_and_ReLU[4].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$3963(.Z({ \dot_product_and_ReLU[4].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$3964(.Z({ \dot_product_and_ReLU[4].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$3965(.Z({ \dot_product_and_ReLU[4].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$3966(.Z({ \dot_product_and_ReLU[4].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$3967(.Z({ \dot_product_and_ReLU[4].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$3968(.Z({ \dot_product_and_ReLU[4].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$3969(.Z({ \dot_product_and_ReLU[4].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$3970(.Z({ \dot_product_and_ReLU[4].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$3971(.Z({ \dot_product_and_ReLU[4].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$3972(.Z({ \dot_product_and_ReLU[4].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$3973(.Z({ \dot_product_and_ReLU[4].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$3974(.Z({ \dot_product_and_ReLU[4].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$3975(.Z({ \dot_product_and_ReLU[4].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$3976(.Z({ \dot_product_and_ReLU[4].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$3977(.Z({ \dot_product_and_ReLU[4].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$3978(.Z({ \dot_product_and_ReLU[4].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$3979(.Z({ \dot_product_and_ReLU[4].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$3980(.Z({ \dot_product_and_ReLU[4].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$3981(.Z({ \dot_product_and_ReLU[4].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$3982(.Z({ \dot_product_and_ReLU[4].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$3983(.Z({ \dot_product_and_ReLU[4].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$3984(.Z({ \dot_product_and_ReLU[4].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$3985(.Z({ \dot_product_and_ReLU[4].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$3986(.Z({ \dot_product_and_ReLU[4].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$3987(.Z({ \dot_product_and_ReLU[4].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$3988(.Z({ \dot_product_and_ReLU[4].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$3989(.Z({ \dot_product_and_ReLU[4].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$3990(.Z({ \dot_product_and_ReLU[4].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$3991(.Z({ \dot_product_and_ReLU[4].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$3992(.Z({ \dot_product_and_ReLU[4].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$3993(.Z({ \dot_product_and_ReLU[4].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$3994(.Z({ \dot_product_and_ReLU[4].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$3995(.Z({ \dot_product_and_ReLU[4].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$3996(.Z({ \dot_product_and_ReLU[4].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$3997(.Z({ \dot_product_and_ReLU[4].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$3998(.Z({ \dot_product_and_ReLU[4].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$3999(.Z({ \dot_product_and_ReLU[4].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$4000(.Z({ \dot_product_and_ReLU[4].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$4001(.Z({ \dot_product_and_ReLU[4].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$4002(.Z({ \dot_product_and_ReLU[4].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$4003(.Z({ \dot_product_and_ReLU[4].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$4004(.Z({ \dot_product_and_ReLU[4].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$4005(.Z({ \dot_product_and_ReLU[4].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$4006(.Z({ \dot_product_and_ReLU[4].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$4007(.Z({ \dot_product_and_ReLU[4].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$4008(.Z({ \dot_product_and_ReLU[4].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$4009(.Z({ \dot_product_and_ReLU[4].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$4010(.Z({ \dot_product_and_ReLU[4].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$4011(.Z({ \dot_product_and_ReLU[4].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$4012(.Z({ \dot_product_and_ReLU[4].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$4013(.Z({ \dot_product_and_ReLU[4].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$4014(.Z({ \dot_product_and_ReLU[4].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$4015(.Z({ \dot_product_and_ReLU[4].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$4016(.Z({ \dot_product_and_ReLU[4].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$4017(.Z({ \dot_product_and_ReLU[4].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$4018(.Z({ \dot_product_and_ReLU[4].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$4019(.Z({ \dot_product_and_ReLU[4].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$4020(.Z({ \dot_product_and_ReLU[4].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$4021(.Z({ \dot_product_and_ReLU[4].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$4022(.Z({ \dot_product_and_ReLU[4].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$4023(.Z({ \dot_product_and_ReLU[4].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$4024(.Z({ \dot_product_and_ReLU[4].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$4025(.Z({ \dot_product_and_ReLU[4].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$4026(.Z({ \dot_product_and_ReLU[4].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$4027(.Z({ \dot_product_and_ReLU[4].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$4028(.Z({ \dot_product_and_ReLU[4].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$4029(.Z({ \dot_product_and_ReLU[4].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$4030(.Z({ \dot_product_and_ReLU[4].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$4031(.Z({ \dot_product_and_ReLU[4].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$4032(.Z({ \dot_product_and_ReLU[4].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$4033(.Z({ \dot_product_and_ReLU[4].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$4034(.Z({ \dot_product_and_ReLU[4].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$4035(.Z({ \dot_product_and_ReLU[4].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$4036(.Z({ \dot_product_and_ReLU[4].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$4037(.Z({ \dot_product_and_ReLU[4].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$4038(.Z({ \dot_product_and_ReLU[4].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$4039(.Z({ \dot_product_and_ReLU[4].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$4040(.Z({ \dot_product_and_ReLU[4].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$4041(.Z({ \dot_product_and_ReLU[4].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$4042(.Z({ \dot_product_and_ReLU[4].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$4043(.Z({ \dot_product_and_ReLU[4].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$4044(.Z({ \dot_product_and_ReLU[4].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$4045(.Z({ \dot_product_and_ReLU[4].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$4046(.Z({ \dot_product_and_ReLU[4].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$4047(.Z({ \dot_product_and_ReLU[4].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$4048(.Z({ \dot_product_and_ReLU[4].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$4049(.Z({ \dot_product_and_ReLU[4].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$4050(.Z({ \dot_product_and_ReLU[4].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$4051(.Z({ \dot_product_and_ReLU[4].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$4052(.Z({ \dot_product_and_ReLU[4].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$4053(.Z({ \dot_product_and_ReLU[4].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$4054(.Z({ \dot_product_and_ReLU[4].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$4055(.Z({ \dot_product_and_ReLU[4].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$4056(.Z({ \dot_product_and_ReLU[4].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$4057(.Z({ \dot_product_and_ReLU[4].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$4058(.Z({ \dot_product_and_ReLU[4].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$4059(.Z({ \dot_product_and_ReLU[4].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$4060(.Z({ \dot_product_and_ReLU[4].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$4061(.Z({ \dot_product_and_ReLU[4].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$4062(.Z({ \dot_product_and_ReLU[4].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$4063(.Z({ \dot_product_and_ReLU[4].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$4064(.Z({ \dot_product_and_ReLU[4].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$4065(.Z({ \dot_product_and_ReLU[4].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$4066(.Z({ \dot_product_and_ReLU[4].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$4067(.Z({ \dot_product_and_ReLU[4].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$4068(.Z({ \dot_product_and_ReLU[4].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$4069(.Z({ \dot_product_and_ReLU[4].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$4070(.Z({ \dot_product_and_ReLU[4].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$4071(.Z({ \dot_product_and_ReLU[4].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$4072(.Z({ \dot_product_and_ReLU[4].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$4073(.Z({ \dot_product_and_ReLU[4].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$4074(.Z({ \dot_product_and_ReLU[4].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$4075(.Z({ \dot_product_and_ReLU[4].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$4076(.Z({ \dot_product_and_ReLU[4].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$4077(.Z({ \dot_product_and_ReLU[4].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$4078(.Z({ \dot_product_and_ReLU[4].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$4079(.Z({ \dot_product_and_ReLU[4].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$4080(.Z({ \dot_product_and_ReLU[4].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$4081(.Z({ \dot_product_and_ReLU[4].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$4082(.Z({ \dot_product_and_ReLU[4].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$4083(.Z({ \dot_product_and_ReLU[4].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$4084(.Z({ \dot_product_and_ReLU[4].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$4085(.Z({ \dot_product_and_ReLU[4].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$4086(.Z({ \dot_product_and_ReLU[4].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$4087(.Z({ \dot_product_and_ReLU[4].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$4088(.Z({ \dot_product_and_ReLU[4].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$4089(.Z({ \dot_product_and_ReLU[4].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$4090(.Z({ \dot_product_and_ReLU[4].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$4091(.Z({ \dot_product_and_ReLU[4].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$4092(.Z({ \dot_product_and_ReLU[4].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$4093(.Z({ \dot_product_and_ReLU[4].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$4094(.Z({ \dot_product_and_ReLU[4].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$4095(.Z({ \dot_product_and_ReLU[4].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$4096(.Z({ \dot_product_and_ReLU[4].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[4][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$4097(.Z({ \dot_product_and_ReLU[3].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$4098(.Z({ \dot_product_and_ReLU[3].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$4099(.Z({ \dot_product_and_ReLU[3].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$4100(.Z({ \dot_product_and_ReLU[3].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$4101(.Z({ \dot_product_and_ReLU[3].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$4102(.Z({ \dot_product_and_ReLU[3].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$4103(.Z({ \dot_product_and_ReLU[3].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$4104(.Z({ \dot_product_and_ReLU[3].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$4105(.Z({ \dot_product_and_ReLU[3].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$4106(.Z({ \dot_product_and_ReLU[3].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$4107(.Z({ \dot_product_and_ReLU[3].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$4108(.Z({ \dot_product_and_ReLU[3].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$4109(.Z({ \dot_product_and_ReLU[3].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$4110(.Z({ \dot_product_and_ReLU[3].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$4111(.Z({ \dot_product_and_ReLU[3].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$4112(.Z({ \dot_product_and_ReLU[3].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$4113(.Z({ \dot_product_and_ReLU[3].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$4114(.Z({ \dot_product_and_ReLU[3].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$4115(.Z({ \dot_product_and_ReLU[3].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$4116(.Z({ \dot_product_and_ReLU[3].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$4117(.Z({ \dot_product_and_ReLU[3].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$4118(.Z({ \dot_product_and_ReLU[3].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$4119(.Z({ \dot_product_and_ReLU[3].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$4120(.Z({ \dot_product_and_ReLU[3].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$4121(.Z({ \dot_product_and_ReLU[3].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$4122(.Z({ \dot_product_and_ReLU[3].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$4123(.Z({ \dot_product_and_ReLU[3].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$4124(.Z({ \dot_product_and_ReLU[3].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$4125(.Z({ \dot_product_and_ReLU[3].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$4126(.Z({ \dot_product_and_ReLU[3].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$4127(.Z({ \dot_product_and_ReLU[3].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$4128(.Z({ \dot_product_and_ReLU[3].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$4129(.Z({ \dot_product_and_ReLU[3].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$4130(.Z({ \dot_product_and_ReLU[3].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$4131(.Z({ \dot_product_and_ReLU[3].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$4132(.Z({ \dot_product_and_ReLU[3].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$4133(.Z({ \dot_product_and_ReLU[3].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$4134(.Z({ \dot_product_and_ReLU[3].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$4135(.Z({ \dot_product_and_ReLU[3].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$4136(.Z({ \dot_product_and_ReLU[3].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$4137(.Z({ \dot_product_and_ReLU[3].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$4138(.Z({ \dot_product_and_ReLU[3].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$4139(.Z({ \dot_product_and_ReLU[3].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$4140(.Z({ \dot_product_and_ReLU[3].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$4141(.Z({ \dot_product_and_ReLU[3].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$4142(.Z({ \dot_product_and_ReLU[3].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$4143(.Z({ \dot_product_and_ReLU[3].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$4144(.Z({ \dot_product_and_ReLU[3].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$4145(.Z({ \dot_product_and_ReLU[3].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$4146(.Z({ \dot_product_and_ReLU[3].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$4147(.Z({ \dot_product_and_ReLU[3].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$4148(.Z({ \dot_product_and_ReLU[3].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$4149(.Z({ \dot_product_and_ReLU[3].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$4150(.Z({ \dot_product_and_ReLU[3].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$4151(.Z({ \dot_product_and_ReLU[3].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$4152(.Z({ \dot_product_and_ReLU[3].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$4153(.Z({ \dot_product_and_ReLU[3].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$4154(.Z({ \dot_product_and_ReLU[3].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$4155(.Z({ \dot_product_and_ReLU[3].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$4156(.Z({ \dot_product_and_ReLU[3].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$4157(.Z({ \dot_product_and_ReLU[3].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$4158(.Z({ \dot_product_and_ReLU[3].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$4159(.Z({ \dot_product_and_ReLU[3].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$4160(.Z({ \dot_product_and_ReLU[3].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$4161(.Z({ \dot_product_and_ReLU[3].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$4162(.Z({ \dot_product_and_ReLU[3].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$4163(.Z({ \dot_product_and_ReLU[3].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$4164(.Z({ \dot_product_and_ReLU[3].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$4165(.Z({ \dot_product_and_ReLU[3].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$4166(.Z({ \dot_product_and_ReLU[3].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$4167(.Z({ \dot_product_and_ReLU[3].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$4168(.Z({ \dot_product_and_ReLU[3].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$4169(.Z({ \dot_product_and_ReLU[3].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$4170(.Z({ \dot_product_and_ReLU[3].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$4171(.Z({ \dot_product_and_ReLU[3].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$4172(.Z({ \dot_product_and_ReLU[3].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$4173(.Z({ \dot_product_and_ReLU[3].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$4174(.Z({ \dot_product_and_ReLU[3].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$4175(.Z({ \dot_product_and_ReLU[3].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$4176(.Z({ \dot_product_and_ReLU[3].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$4177(.Z({ \dot_product_and_ReLU[3].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$4178(.Z({ \dot_product_and_ReLU[3].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$4179(.Z({ \dot_product_and_ReLU[3].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$4180(.Z({ \dot_product_and_ReLU[3].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$4181(.Z({ \dot_product_and_ReLU[3].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$4182(.Z({ \dot_product_and_ReLU[3].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$4183(.Z({ \dot_product_and_ReLU[3].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$4184(.Z({ \dot_product_and_ReLU[3].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$4185(.Z({ \dot_product_and_ReLU[3].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$4186(.Z({ \dot_product_and_ReLU[3].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$4187(.Z({ \dot_product_and_ReLU[3].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$4188(.Z({ \dot_product_and_ReLU[3].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$4189(.Z({ \dot_product_and_ReLU[3].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$4190(.Z({ \dot_product_and_ReLU[3].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$4191(.Z({ \dot_product_and_ReLU[3].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$4192(.Z({ \dot_product_and_ReLU[3].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$4193(.Z({ \dot_product_and_ReLU[3].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$4194(.Z({ \dot_product_and_ReLU[3].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$4195(.Z({ \dot_product_and_ReLU[3].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$4196(.Z({ \dot_product_and_ReLU[3].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$4197(.Z({ \dot_product_and_ReLU[3].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$4198(.Z({ \dot_product_and_ReLU[3].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$4199(.Z({ \dot_product_and_ReLU[3].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$4200(.Z({ \dot_product_and_ReLU[3].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$4201(.Z({ \dot_product_and_ReLU[3].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$4202(.Z({ \dot_product_and_ReLU[3].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$4203(.Z({ \dot_product_and_ReLU[3].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$4204(.Z({ \dot_product_and_ReLU[3].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$4205(.Z({ \dot_product_and_ReLU[3].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$4206(.Z({ \dot_product_and_ReLU[3].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$4207(.Z({ \dot_product_and_ReLU[3].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$4208(.Z({ \dot_product_and_ReLU[3].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$4209(.Z({ \dot_product_and_ReLU[3].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$4210(.Z({ \dot_product_and_ReLU[3].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$4211(.Z({ \dot_product_and_ReLU[3].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$4212(.Z({ \dot_product_and_ReLU[3].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$4213(.Z({ \dot_product_and_ReLU[3].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$4214(.Z({ \dot_product_and_ReLU[3].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$4215(.Z({ \dot_product_and_ReLU[3].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$4216(.Z({ \dot_product_and_ReLU[3].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$4217(.Z({ \dot_product_and_ReLU[3].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$4218(.Z({ \dot_product_and_ReLU[3].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$4219(.Z({ \dot_product_and_ReLU[3].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$4220(.Z({ \dot_product_and_ReLU[3].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$4221(.Z({ \dot_product_and_ReLU[3].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$4222(.Z({ \dot_product_and_ReLU[3].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$4223(.Z({ \dot_product_and_ReLU[3].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$4224(.Z({ \dot_product_and_ReLU[3].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$4225(.Z({ \dot_product_and_ReLU[3].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$4226(.Z({ \dot_product_and_ReLU[3].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$4227(.Z({ \dot_product_and_ReLU[3].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$4228(.Z({ \dot_product_and_ReLU[3].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$4229(.Z({ \dot_product_and_ReLU[3].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$4230(.Z({ \dot_product_and_ReLU[3].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$4231(.Z({ \dot_product_and_ReLU[3].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$4232(.Z({ \dot_product_and_ReLU[3].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$4233(.Z({ \dot_product_and_ReLU[3].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$4234(.Z({ \dot_product_and_ReLU[3].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$4235(.Z({ \dot_product_and_ReLU[3].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$4236(.Z({ \dot_product_and_ReLU[3].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$4237(.Z({ \dot_product_and_ReLU[3].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$4238(.Z({ \dot_product_and_ReLU[3].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$4239(.Z({ \dot_product_and_ReLU[3].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$4240(.Z({ \dot_product_and_ReLU[3].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$4241(.Z({ \dot_product_and_ReLU[3].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$4242(.Z({ \dot_product_and_ReLU[3].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$4243(.Z({ \dot_product_and_ReLU[3].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$4244(.Z({ \dot_product_and_ReLU[3].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$4245(.Z({ \dot_product_and_ReLU[3].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$4246(.Z({ \dot_product_and_ReLU[3].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$4247(.Z({ \dot_product_and_ReLU[3].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$4248(.Z({ \dot_product_and_ReLU[3].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$4249(.Z({ \dot_product_and_ReLU[3].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$4250(.Z({ \dot_product_and_ReLU[3].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$4251(.Z({ \dot_product_and_ReLU[3].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$4252(.Z({ \dot_product_and_ReLU[3].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$4253(.Z({ \dot_product_and_ReLU[3].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$4254(.Z({ \dot_product_and_ReLU[3].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$4255(.Z({ \dot_product_and_ReLU[3].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$4256(.Z({ \dot_product_and_ReLU[3].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$4257(.Z({ \dot_product_and_ReLU[3].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$4258(.Z({ \dot_product_and_ReLU[3].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$4259(.Z({ \dot_product_and_ReLU[3].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$4260(.Z({ \dot_product_and_ReLU[3].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$4261(.Z({ \dot_product_and_ReLU[3].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$4262(.Z({ \dot_product_and_ReLU[3].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$4263(.Z({ \dot_product_and_ReLU[3].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$4264(.Z({ \dot_product_and_ReLU[3].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$4265(.Z({ \dot_product_and_ReLU[3].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$4266(.Z({ \dot_product_and_ReLU[3].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$4267(.Z({ \dot_product_and_ReLU[3].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$4268(.Z({ \dot_product_and_ReLU[3].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$4269(.Z({ \dot_product_and_ReLU[3].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$4270(.Z({ \dot_product_and_ReLU[3].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$4271(.Z({ \dot_product_and_ReLU[3].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$4272(.Z({ \dot_product_and_ReLU[3].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$4273(.Z({ \dot_product_and_ReLU[3].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$4274(.Z({ \dot_product_and_ReLU[3].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$4275(.Z({ \dot_product_and_ReLU[3].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$4276(.Z({ \dot_product_and_ReLU[3].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$4277(.Z({ \dot_product_and_ReLU[3].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$4278(.Z({ \dot_product_and_ReLU[3].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$4279(.Z({ \dot_product_and_ReLU[3].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$4280(.Z({ \dot_product_and_ReLU[3].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$4281(.Z({ \dot_product_and_ReLU[3].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$4282(.Z({ \dot_product_and_ReLU[3].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$4283(.Z({ \dot_product_and_ReLU[3].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$4284(.Z({ \dot_product_and_ReLU[3].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$4285(.Z({ \dot_product_and_ReLU[3].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$4286(.Z({ \dot_product_and_ReLU[3].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$4287(.Z({ \dot_product_and_ReLU[3].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$4288(.Z({ \dot_product_and_ReLU[3].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$4289(.Z({ \dot_product_and_ReLU[3].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$4290(.Z({ \dot_product_and_ReLU[3].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$4291(.Z({ \dot_product_and_ReLU[3].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$4292(.Z({ \dot_product_and_ReLU[3].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$4293(.Z({ \dot_product_and_ReLU[3].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$4294(.Z({ \dot_product_and_ReLU[3].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$4295(.Z({ \dot_product_and_ReLU[3].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$4296(.Z({ \dot_product_and_ReLU[3].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$4297(.Z({ \dot_product_and_ReLU[3].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$4298(.Z({ \dot_product_and_ReLU[3].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$4299(.Z({ \dot_product_and_ReLU[3].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$4300(.Z({ \dot_product_and_ReLU[3].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$4301(.Z({ \dot_product_and_ReLU[3].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$4302(.Z({ \dot_product_and_ReLU[3].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$4303(.Z({ \dot_product_and_ReLU[3].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$4304(.Z({ \dot_product_and_ReLU[3].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$4305(.Z({ \dot_product_and_ReLU[3].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$4306(.Z({ \dot_product_and_ReLU[3].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$4307(.Z({ \dot_product_and_ReLU[3].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$4308(.Z({ \dot_product_and_ReLU[3].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$4309(.Z({ \dot_product_and_ReLU[3].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$4310(.Z({ \dot_product_and_ReLU[3].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$4311(.Z({ \dot_product_and_ReLU[3].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$4312(.Z({ \dot_product_and_ReLU[3].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$4313(.Z({ \dot_product_and_ReLU[3].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$4314(.Z({ \dot_product_and_ReLU[3].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$4315(.Z({ \dot_product_and_ReLU[3].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$4316(.Z({ \dot_product_and_ReLU[3].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$4317(.Z({ \dot_product_and_ReLU[3].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$4318(.Z({ \dot_product_and_ReLU[3].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$4319(.Z({ \dot_product_and_ReLU[3].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$4320(.Z({ \dot_product_and_ReLU[3].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$4321(.Z({ \dot_product_and_ReLU[3].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$4322(.Z({ \dot_product_and_ReLU[3].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$4323(.Z({ \dot_product_and_ReLU[3].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$4324(.Z({ \dot_product_and_ReLU[3].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$4325(.Z({ \dot_product_and_ReLU[3].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$4326(.Z({ \dot_product_and_ReLU[3].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$4327(.Z({ \dot_product_and_ReLU[3].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$4328(.Z({ \dot_product_and_ReLU[3].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$4329(.Z({ \dot_product_and_ReLU[3].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$4330(.Z({ \dot_product_and_ReLU[3].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$4331(.Z({ \dot_product_and_ReLU[3].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$4332(.Z({ \dot_product_and_ReLU[3].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$4333(.Z({ \dot_product_and_ReLU[3].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$4334(.Z({ \dot_product_and_ReLU[3].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$4335(.Z({ \dot_product_and_ReLU[3].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$4336(.Z({ \dot_product_and_ReLU[3].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$4337(.Z({ \dot_product_and_ReLU[3].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$4338(.Z({ \dot_product_and_ReLU[3].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$4339(.Z({ \dot_product_and_ReLU[3].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$4340(.Z({ \dot_product_and_ReLU[3].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$4341(.Z({ \dot_product_and_ReLU[3].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$4342(.Z({ \dot_product_and_ReLU[3].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$4343(.Z({ \dot_product_and_ReLU[3].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$4344(.Z({ \dot_product_and_ReLU[3].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$4345(.Z({ \dot_product_and_ReLU[3].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$4346(.Z({ \dot_product_and_ReLU[3].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$4347(.Z({ \dot_product_and_ReLU[3].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$4348(.Z({ \dot_product_and_ReLU[3].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$4349(.Z({ \dot_product_and_ReLU[3].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$4350(.Z({ \dot_product_and_ReLU[3].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$4351(.Z({ \dot_product_and_ReLU[3].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$4352(.Z({ \dot_product_and_ReLU[3].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[3][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$4353(.Z({ \dot_product_and_ReLU[2].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$4354(.Z({ \dot_product_and_ReLU[2].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$4355(.Z({ \dot_product_and_ReLU[2].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$4356(.Z({ \dot_product_and_ReLU[2].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$4357(.Z({ \dot_product_and_ReLU[2].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$4358(.Z({ \dot_product_and_ReLU[2].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$4359(.Z({ \dot_product_and_ReLU[2].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$4360(.Z({ \dot_product_and_ReLU[2].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$4361(.Z({ \dot_product_and_ReLU[2].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$4362(.Z({ \dot_product_and_ReLU[2].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$4363(.Z({ \dot_product_and_ReLU[2].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$4364(.Z({ \dot_product_and_ReLU[2].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$4365(.Z({ \dot_product_and_ReLU[2].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$4366(.Z({ \dot_product_and_ReLU[2].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$4367(.Z({ \dot_product_and_ReLU[2].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$4368(.Z({ \dot_product_and_ReLU[2].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$4369(.Z({ \dot_product_and_ReLU[2].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$4370(.Z({ \dot_product_and_ReLU[2].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$4371(.Z({ \dot_product_and_ReLU[2].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$4372(.Z({ \dot_product_and_ReLU[2].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$4373(.Z({ \dot_product_and_ReLU[2].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$4374(.Z({ \dot_product_and_ReLU[2].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$4375(.Z({ \dot_product_and_ReLU[2].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$4376(.Z({ \dot_product_and_ReLU[2].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$4377(.Z({ \dot_product_and_ReLU[2].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$4378(.Z({ \dot_product_and_ReLU[2].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$4379(.Z({ \dot_product_and_ReLU[2].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$4380(.Z({ \dot_product_and_ReLU[2].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$4381(.Z({ \dot_product_and_ReLU[2].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$4382(.Z({ \dot_product_and_ReLU[2].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$4383(.Z({ \dot_product_and_ReLU[2].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$4384(.Z({ \dot_product_and_ReLU[2].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$4385(.Z({ \dot_product_and_ReLU[2].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$4386(.Z({ \dot_product_and_ReLU[2].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$4387(.Z({ \dot_product_and_ReLU[2].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$4388(.Z({ \dot_product_and_ReLU[2].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$4389(.Z({ \dot_product_and_ReLU[2].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$4390(.Z({ \dot_product_and_ReLU[2].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$4391(.Z({ \dot_product_and_ReLU[2].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$4392(.Z({ \dot_product_and_ReLU[2].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$4393(.Z({ \dot_product_and_ReLU[2].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$4394(.Z({ \dot_product_and_ReLU[2].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$4395(.Z({ \dot_product_and_ReLU[2].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$4396(.Z({ \dot_product_and_ReLU[2].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$4397(.Z({ \dot_product_and_ReLU[2].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$4398(.Z({ \dot_product_and_ReLU[2].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$4399(.Z({ \dot_product_and_ReLU[2].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$4400(.Z({ \dot_product_and_ReLU[2].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$4401(.Z({ \dot_product_and_ReLU[2].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$4402(.Z({ \dot_product_and_ReLU[2].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$4403(.Z({ \dot_product_and_ReLU[2].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$4404(.Z({ \dot_product_and_ReLU[2].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$4405(.Z({ \dot_product_and_ReLU[2].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$4406(.Z({ \dot_product_and_ReLU[2].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$4407(.Z({ \dot_product_and_ReLU[2].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$4408(.Z({ \dot_product_and_ReLU[2].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$4409(.Z({ \dot_product_and_ReLU[2].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$4410(.Z({ \dot_product_and_ReLU[2].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$4411(.Z({ \dot_product_and_ReLU[2].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$4412(.Z({ \dot_product_and_ReLU[2].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$4413(.Z({ \dot_product_and_ReLU[2].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$4414(.Z({ \dot_product_and_ReLU[2].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$4415(.Z({ \dot_product_and_ReLU[2].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$4416(.Z({ \dot_product_and_ReLU[2].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$4417(.Z({ \dot_product_and_ReLU[2].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$4418(.Z({ \dot_product_and_ReLU[2].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$4419(.Z({ \dot_product_and_ReLU[2].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$4420(.Z({ \dot_product_and_ReLU[2].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$4421(.Z({ \dot_product_and_ReLU[2].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$4422(.Z({ \dot_product_and_ReLU[2].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$4423(.Z({ \dot_product_and_ReLU[2].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$4424(.Z({ \dot_product_and_ReLU[2].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$4425(.Z({ \dot_product_and_ReLU[2].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$4426(.Z({ \dot_product_and_ReLU[2].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$4427(.Z({ \dot_product_and_ReLU[2].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$4428(.Z({ \dot_product_and_ReLU[2].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$4429(.Z({ \dot_product_and_ReLU[2].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$4430(.Z({ \dot_product_and_ReLU[2].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$4431(.Z({ \dot_product_and_ReLU[2].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$4432(.Z({ \dot_product_and_ReLU[2].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$4433(.Z({ \dot_product_and_ReLU[2].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$4434(.Z({ \dot_product_and_ReLU[2].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$4435(.Z({ \dot_product_and_ReLU[2].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$4436(.Z({ \dot_product_and_ReLU[2].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$4437(.Z({ \dot_product_and_ReLU[2].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$4438(.Z({ \dot_product_and_ReLU[2].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$4439(.Z({ \dot_product_and_ReLU[2].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$4440(.Z({ \dot_product_and_ReLU[2].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$4441(.Z({ \dot_product_and_ReLU[2].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$4442(.Z({ \dot_product_and_ReLU[2].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$4443(.Z({ \dot_product_and_ReLU[2].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$4444(.Z({ \dot_product_and_ReLU[2].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$4445(.Z({ \dot_product_and_ReLU[2].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$4446(.Z({ \dot_product_and_ReLU[2].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$4447(.Z({ \dot_product_and_ReLU[2].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$4448(.Z({ \dot_product_and_ReLU[2].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$4449(.Z({ \dot_product_and_ReLU[2].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$4450(.Z({ \dot_product_and_ReLU[2].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$4451(.Z({ \dot_product_and_ReLU[2].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$4452(.Z({ \dot_product_and_ReLU[2].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$4453(.Z({ \dot_product_and_ReLU[2].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$4454(.Z({ \dot_product_and_ReLU[2].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$4455(.Z({ \dot_product_and_ReLU[2].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$4456(.Z({ \dot_product_and_ReLU[2].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$4457(.Z({ \dot_product_and_ReLU[2].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$4458(.Z({ \dot_product_and_ReLU[2].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$4459(.Z({ \dot_product_and_ReLU[2].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$4460(.Z({ \dot_product_and_ReLU[2].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$4461(.Z({ \dot_product_and_ReLU[2].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$4462(.Z({ \dot_product_and_ReLU[2].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$4463(.Z({ \dot_product_and_ReLU[2].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$4464(.Z({ \dot_product_and_ReLU[2].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$4465(.Z({ \dot_product_and_ReLU[2].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$4466(.Z({ \dot_product_and_ReLU[2].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$4467(.Z({ \dot_product_and_ReLU[2].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$4468(.Z({ \dot_product_and_ReLU[2].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$4469(.Z({ \dot_product_and_ReLU[2].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$4470(.Z({ \dot_product_and_ReLU[2].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$4471(.Z({ \dot_product_and_ReLU[2].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$4472(.Z({ \dot_product_and_ReLU[2].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$4473(.Z({ \dot_product_and_ReLU[2].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$4474(.Z({ \dot_product_and_ReLU[2].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$4475(.Z({ \dot_product_and_ReLU[2].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$4476(.Z({ \dot_product_and_ReLU[2].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$4477(.Z({ \dot_product_and_ReLU[2].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$4478(.Z({ \dot_product_and_ReLU[2].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$4479(.Z({ \dot_product_and_ReLU[2].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$4480(.Z({ \dot_product_and_ReLU[2].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$4481(.Z({ \dot_product_and_ReLU[2].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$4482(.Z({ \dot_product_and_ReLU[2].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$4483(.Z({ \dot_product_and_ReLU[2].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$4484(.Z({ \dot_product_and_ReLU[2].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$4485(.Z({ \dot_product_and_ReLU[2].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$4486(.Z({ \dot_product_and_ReLU[2].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$4487(.Z({ \dot_product_and_ReLU[2].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$4488(.Z({ \dot_product_and_ReLU[2].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$4489(.Z({ \dot_product_and_ReLU[2].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$4490(.Z({ \dot_product_and_ReLU[2].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$4491(.Z({ \dot_product_and_ReLU[2].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$4492(.Z({ \dot_product_and_ReLU[2].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$4493(.Z({ \dot_product_and_ReLU[2].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$4494(.Z({ \dot_product_and_ReLU[2].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$4495(.Z({ \dot_product_and_ReLU[2].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$4496(.Z({ \dot_product_and_ReLU[2].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$4497(.Z({ \dot_product_and_ReLU[2].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$4498(.Z({ \dot_product_and_ReLU[2].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$4499(.Z({ \dot_product_and_ReLU[2].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$4500(.Z({ \dot_product_and_ReLU[2].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$4501(.Z({ \dot_product_and_ReLU[2].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$4502(.Z({ \dot_product_and_ReLU[2].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$4503(.Z({ \dot_product_and_ReLU[2].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$4504(.Z({ \dot_product_and_ReLU[2].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$4505(.Z({ \dot_product_and_ReLU[2].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$4506(.Z({ \dot_product_and_ReLU[2].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$4507(.Z({ \dot_product_and_ReLU[2].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$4508(.Z({ \dot_product_and_ReLU[2].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$4509(.Z({ \dot_product_and_ReLU[2].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$4510(.Z({ \dot_product_and_ReLU[2].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$4511(.Z({ \dot_product_and_ReLU[2].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$4512(.Z({ \dot_product_and_ReLU[2].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$4513(.Z({ \dot_product_and_ReLU[2].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$4514(.Z({ \dot_product_and_ReLU[2].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$4515(.Z({ \dot_product_and_ReLU[2].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$4516(.Z({ \dot_product_and_ReLU[2].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$4517(.Z({ \dot_product_and_ReLU[2].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$4518(.Z({ \dot_product_and_ReLU[2].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$4519(.Z({ \dot_product_and_ReLU[2].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$4520(.Z({ \dot_product_and_ReLU[2].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$4521(.Z({ \dot_product_and_ReLU[2].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$4522(.Z({ \dot_product_and_ReLU[2].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$4523(.Z({ \dot_product_and_ReLU[2].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$4524(.Z({ \dot_product_and_ReLU[2].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$4525(.Z({ \dot_product_and_ReLU[2].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$4526(.Z({ \dot_product_and_ReLU[2].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$4527(.Z({ \dot_product_and_ReLU[2].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$4528(.Z({ \dot_product_and_ReLU[2].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$4529(.Z({ \dot_product_and_ReLU[2].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$4530(.Z({ \dot_product_and_ReLU[2].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$4531(.Z({ \dot_product_and_ReLU[2].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$4532(.Z({ \dot_product_and_ReLU[2].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$4533(.Z({ \dot_product_and_ReLU[2].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$4534(.Z({ \dot_product_and_ReLU[2].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$4535(.Z({ \dot_product_and_ReLU[2].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$4536(.Z({ \dot_product_and_ReLU[2].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$4537(.Z({ \dot_product_and_ReLU[2].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$4538(.Z({ \dot_product_and_ReLU[2].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$4539(.Z({ \dot_product_and_ReLU[2].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$4540(.Z({ \dot_product_and_ReLU[2].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$4541(.Z({ \dot_product_and_ReLU[2].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$4542(.Z({ \dot_product_and_ReLU[2].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$4543(.Z({ \dot_product_and_ReLU[2].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$4544(.Z({ \dot_product_and_ReLU[2].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$4545(.Z({ \dot_product_and_ReLU[2].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$4546(.Z({ \dot_product_and_ReLU[2].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$4547(.Z({ \dot_product_and_ReLU[2].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$4548(.Z({ \dot_product_and_ReLU[2].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$4549(.Z({ \dot_product_and_ReLU[2].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$4550(.Z({ \dot_product_and_ReLU[2].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$4551(.Z({ \dot_product_and_ReLU[2].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$4552(.Z({ \dot_product_and_ReLU[2].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$4553(.Z({ \dot_product_and_ReLU[2].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$4554(.Z({ \dot_product_and_ReLU[2].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$4555(.Z({ \dot_product_and_ReLU[2].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$4556(.Z({ \dot_product_and_ReLU[2].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$4557(.Z({ \dot_product_and_ReLU[2].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$4558(.Z({ \dot_product_and_ReLU[2].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$4559(.Z({ \dot_product_and_ReLU[2].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$4560(.Z({ \dot_product_and_ReLU[2].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$4561(.Z({ \dot_product_and_ReLU[2].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$4562(.Z({ \dot_product_and_ReLU[2].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$4563(.Z({ \dot_product_and_ReLU[2].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$4564(.Z({ \dot_product_and_ReLU[2].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$4565(.Z({ \dot_product_and_ReLU[2].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$4566(.Z({ \dot_product_and_ReLU[2].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$4567(.Z({ \dot_product_and_ReLU[2].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$4568(.Z({ \dot_product_and_ReLU[2].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$4569(.Z({ \dot_product_and_ReLU[2].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$4570(.Z({ \dot_product_and_ReLU[2].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$4571(.Z({ \dot_product_and_ReLU[2].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$4572(.Z({ \dot_product_and_ReLU[2].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$4573(.Z({ \dot_product_and_ReLU[2].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$4574(.Z({ \dot_product_and_ReLU[2].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$4575(.Z({ \dot_product_and_ReLU[2].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$4576(.Z({ \dot_product_and_ReLU[2].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$4577(.Z({ \dot_product_and_ReLU[2].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$4578(.Z({ \dot_product_and_ReLU[2].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$4579(.Z({ \dot_product_and_ReLU[2].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$4580(.Z({ \dot_product_and_ReLU[2].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$4581(.Z({ \dot_product_and_ReLU[2].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$4582(.Z({ \dot_product_and_ReLU[2].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$4583(.Z({ \dot_product_and_ReLU[2].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$4584(.Z({ \dot_product_and_ReLU[2].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$4585(.Z({ \dot_product_and_ReLU[2].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$4586(.Z({ \dot_product_and_ReLU[2].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$4587(.Z({ \dot_product_and_ReLU[2].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$4588(.Z({ \dot_product_and_ReLU[2].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$4589(.Z({ \dot_product_and_ReLU[2].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$4590(.Z({ \dot_product_and_ReLU[2].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$4591(.Z({ \dot_product_and_ReLU[2].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$4592(.Z({ \dot_product_and_ReLU[2].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$4593(.Z({ \dot_product_and_ReLU[2].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$4594(.Z({ \dot_product_and_ReLU[2].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$4595(.Z({ \dot_product_and_ReLU[2].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$4596(.Z({ \dot_product_and_ReLU[2].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$4597(.Z({ \dot_product_and_ReLU[2].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$4598(.Z({ \dot_product_and_ReLU[2].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$4599(.Z({ \dot_product_and_ReLU[2].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$4600(.Z({ \dot_product_and_ReLU[2].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$4601(.Z({ \dot_product_and_ReLU[2].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$4602(.Z({ \dot_product_and_ReLU[2].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$4603(.Z({ \dot_product_and_ReLU[2].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$4604(.Z({ \dot_product_and_ReLU[2].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$4605(.Z({ \dot_product_and_ReLU[2].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$4606(.Z({ \dot_product_and_ReLU[2].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$4607(.Z({ \dot_product_and_ReLU[2].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$4608(.Z({ \dot_product_and_ReLU[2].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[2][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$4609(.Z({ \dot_product_and_ReLU[1].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$4610(.Z({ \dot_product_and_ReLU[1].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$4611(.Z({ \dot_product_and_ReLU[1].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$4612(.Z({ \dot_product_and_ReLU[1].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$4613(.Z({ \dot_product_and_ReLU[1].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$4614(.Z({ \dot_product_and_ReLU[1].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$4615(.Z({ \dot_product_and_ReLU[1].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$4616(.Z({ \dot_product_and_ReLU[1].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$4617(.Z({ \dot_product_and_ReLU[1].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$4618(.Z({ \dot_product_and_ReLU[1].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$4619(.Z({ \dot_product_and_ReLU[1].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$4620(.Z({ \dot_product_and_ReLU[1].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$4621(.Z({ \dot_product_and_ReLU[1].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$4622(.Z({ \dot_product_and_ReLU[1].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$4623(.Z({ \dot_product_and_ReLU[1].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$4624(.Z({ \dot_product_and_ReLU[1].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$4625(.Z({ \dot_product_and_ReLU[1].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$4626(.Z({ \dot_product_and_ReLU[1].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$4627(.Z({ \dot_product_and_ReLU[1].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$4628(.Z({ \dot_product_and_ReLU[1].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$4629(.Z({ \dot_product_and_ReLU[1].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$4630(.Z({ \dot_product_and_ReLU[1].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$4631(.Z({ \dot_product_and_ReLU[1].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$4632(.Z({ \dot_product_and_ReLU[1].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$4633(.Z({ \dot_product_and_ReLU[1].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$4634(.Z({ \dot_product_and_ReLU[1].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$4635(.Z({ \dot_product_and_ReLU[1].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$4636(.Z({ \dot_product_and_ReLU[1].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$4637(.Z({ \dot_product_and_ReLU[1].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$4638(.Z({ \dot_product_and_ReLU[1].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$4639(.Z({ \dot_product_and_ReLU[1].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$4640(.Z({ \dot_product_and_ReLU[1].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$4641(.Z({ \dot_product_and_ReLU[1].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$4642(.Z({ \dot_product_and_ReLU[1].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$4643(.Z({ \dot_product_and_ReLU[1].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$4644(.Z({ \dot_product_and_ReLU[1].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$4645(.Z({ \dot_product_and_ReLU[1].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$4646(.Z({ \dot_product_and_ReLU[1].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$4647(.Z({ \dot_product_and_ReLU[1].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$4648(.Z({ \dot_product_and_ReLU[1].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$4649(.Z({ \dot_product_and_ReLU[1].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$4650(.Z({ \dot_product_and_ReLU[1].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$4651(.Z({ \dot_product_and_ReLU[1].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$4652(.Z({ \dot_product_and_ReLU[1].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$4653(.Z({ \dot_product_and_ReLU[1].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$4654(.Z({ \dot_product_and_ReLU[1].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$4655(.Z({ \dot_product_and_ReLU[1].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$4656(.Z({ \dot_product_and_ReLU[1].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$4657(.Z({ \dot_product_and_ReLU[1].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$4658(.Z({ \dot_product_and_ReLU[1].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$4659(.Z({ \dot_product_and_ReLU[1].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$4660(.Z({ \dot_product_and_ReLU[1].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$4661(.Z({ \dot_product_and_ReLU[1].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$4662(.Z({ \dot_product_and_ReLU[1].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$4663(.Z({ \dot_product_and_ReLU[1].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$4664(.Z({ \dot_product_and_ReLU[1].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$4665(.Z({ \dot_product_and_ReLU[1].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$4666(.Z({ \dot_product_and_ReLU[1].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$4667(.Z({ \dot_product_and_ReLU[1].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$4668(.Z({ \dot_product_and_ReLU[1].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$4669(.Z({ \dot_product_and_ReLU[1].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$4670(.Z({ \dot_product_and_ReLU[1].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$4671(.Z({ \dot_product_and_ReLU[1].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$4672(.Z({ \dot_product_and_ReLU[1].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$4673(.Z({ \dot_product_and_ReLU[1].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$4674(.Z({ \dot_product_and_ReLU[1].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$4675(.Z({ \dot_product_and_ReLU[1].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$4676(.Z({ \dot_product_and_ReLU[1].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$4677(.Z({ \dot_product_and_ReLU[1].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$4678(.Z({ \dot_product_and_ReLU[1].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$4679(.Z({ \dot_product_and_ReLU[1].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$4680(.Z({ \dot_product_and_ReLU[1].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$4681(.Z({ \dot_product_and_ReLU[1].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$4682(.Z({ \dot_product_and_ReLU[1].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$4683(.Z({ \dot_product_and_ReLU[1].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$4684(.Z({ \dot_product_and_ReLU[1].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$4685(.Z({ \dot_product_and_ReLU[1].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$4686(.Z({ \dot_product_and_ReLU[1].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$4687(.Z({ \dot_product_and_ReLU[1].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$4688(.Z({ \dot_product_and_ReLU[1].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$4689(.Z({ \dot_product_and_ReLU[1].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$4690(.Z({ \dot_product_and_ReLU[1].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$4691(.Z({ \dot_product_and_ReLU[1].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$4692(.Z({ \dot_product_and_ReLU[1].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$4693(.Z({ \dot_product_and_ReLU[1].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$4694(.Z({ \dot_product_and_ReLU[1].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$4695(.Z({ \dot_product_and_ReLU[1].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$4696(.Z({ \dot_product_and_ReLU[1].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$4697(.Z({ \dot_product_and_ReLU[1].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$4698(.Z({ \dot_product_and_ReLU[1].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$4699(.Z({ \dot_product_and_ReLU[1].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$4700(.Z({ \dot_product_and_ReLU[1].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$4701(.Z({ \dot_product_and_ReLU[1].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$4702(.Z({ \dot_product_and_ReLU[1].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$4703(.Z({ \dot_product_and_ReLU[1].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$4704(.Z({ \dot_product_and_ReLU[1].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$4705(.Z({ \dot_product_and_ReLU[1].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$4706(.Z({ \dot_product_and_ReLU[1].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$4707(.Z({ \dot_product_and_ReLU[1].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$4708(.Z({ \dot_product_and_ReLU[1].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$4709(.Z({ \dot_product_and_ReLU[1].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$4710(.Z({ \dot_product_and_ReLU[1].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$4711(.Z({ \dot_product_and_ReLU[1].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$4712(.Z({ \dot_product_and_ReLU[1].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$4713(.Z({ \dot_product_and_ReLU[1].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$4714(.Z({ \dot_product_and_ReLU[1].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$4715(.Z({ \dot_product_and_ReLU[1].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$4716(.Z({ \dot_product_and_ReLU[1].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$4717(.Z({ \dot_product_and_ReLU[1].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$4718(.Z({ \dot_product_and_ReLU[1].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$4719(.Z({ \dot_product_and_ReLU[1].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$4720(.Z({ \dot_product_and_ReLU[1].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$4721(.Z({ \dot_product_and_ReLU[1].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$4722(.Z({ \dot_product_and_ReLU[1].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$4723(.Z({ \dot_product_and_ReLU[1].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$4724(.Z({ \dot_product_and_ReLU[1].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$4725(.Z({ \dot_product_and_ReLU[1].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$4726(.Z({ \dot_product_and_ReLU[1].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$4727(.Z({ \dot_product_and_ReLU[1].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$4728(.Z({ \dot_product_and_ReLU[1].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$4729(.Z({ \dot_product_and_ReLU[1].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$4730(.Z({ \dot_product_and_ReLU[1].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$4731(.Z({ \dot_product_and_ReLU[1].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$4732(.Z({ \dot_product_and_ReLU[1].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$4733(.Z({ \dot_product_and_ReLU[1].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$4734(.Z({ \dot_product_and_ReLU[1].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$4735(.Z({ \dot_product_and_ReLU[1].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$4736(.Z({ \dot_product_and_ReLU[1].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$4737(.Z({ \dot_product_and_ReLU[1].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$4738(.Z({ \dot_product_and_ReLU[1].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$4739(.Z({ \dot_product_and_ReLU[1].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$4740(.Z({ \dot_product_and_ReLU[1].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$4741(.Z({ \dot_product_and_ReLU[1].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$4742(.Z({ \dot_product_and_ReLU[1].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$4743(.Z({ \dot_product_and_ReLU[1].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$4744(.Z({ \dot_product_and_ReLU[1].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$4745(.Z({ \dot_product_and_ReLU[1].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$4746(.Z({ \dot_product_and_ReLU[1].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$4747(.Z({ \dot_product_and_ReLU[1].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$4748(.Z({ \dot_product_and_ReLU[1].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$4749(.Z({ \dot_product_and_ReLU[1].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$4750(.Z({ \dot_product_and_ReLU[1].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$4751(.Z({ \dot_product_and_ReLU[1].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$4752(.Z({ \dot_product_and_ReLU[1].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$4753(.Z({ \dot_product_and_ReLU[1].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$4754(.Z({ \dot_product_and_ReLU[1].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$4755(.Z({ \dot_product_and_ReLU[1].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$4756(.Z({ \dot_product_and_ReLU[1].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$4757(.Z({ \dot_product_and_ReLU[1].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$4758(.Z({ \dot_product_and_ReLU[1].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$4759(.Z({ \dot_product_and_ReLU[1].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$4760(.Z({ \dot_product_and_ReLU[1].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$4761(.Z({ \dot_product_and_ReLU[1].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$4762(.Z({ \dot_product_and_ReLU[1].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$4763(.Z({ \dot_product_and_ReLU[1].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$4764(.Z({ \dot_product_and_ReLU[1].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$4765(.Z({ \dot_product_and_ReLU[1].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$4766(.Z({ \dot_product_and_ReLU[1].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$4767(.Z({ \dot_product_and_ReLU[1].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$4768(.Z({ \dot_product_and_ReLU[1].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$4769(.Z({ \dot_product_and_ReLU[1].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$4770(.Z({ \dot_product_and_ReLU[1].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$4771(.Z({ \dot_product_and_ReLU[1].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$4772(.Z({ \dot_product_and_ReLU[1].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$4773(.Z({ \dot_product_and_ReLU[1].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$4774(.Z({ \dot_product_and_ReLU[1].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$4775(.Z({ \dot_product_and_ReLU[1].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$4776(.Z({ \dot_product_and_ReLU[1].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$4777(.Z({ \dot_product_and_ReLU[1].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$4778(.Z({ \dot_product_and_ReLU[1].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$4779(.Z({ \dot_product_and_ReLU[1].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$4780(.Z({ \dot_product_and_ReLU[1].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$4781(.Z({ \dot_product_and_ReLU[1].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$4782(.Z({ \dot_product_and_ReLU[1].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$4783(.Z({ \dot_product_and_ReLU[1].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$4784(.Z({ \dot_product_and_ReLU[1].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$4785(.Z({ \dot_product_and_ReLU[1].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$4786(.Z({ \dot_product_and_ReLU[1].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$4787(.Z({ \dot_product_and_ReLU[1].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$4788(.Z({ \dot_product_and_ReLU[1].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$4789(.Z({ \dot_product_and_ReLU[1].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$4790(.Z({ \dot_product_and_ReLU[1].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$4791(.Z({ \dot_product_and_ReLU[1].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$4792(.Z({ \dot_product_and_ReLU[1].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$4793(.Z({ \dot_product_and_ReLU[1].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$4794(.Z({ \dot_product_and_ReLU[1].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$4795(.Z({ \dot_product_and_ReLU[1].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$4796(.Z({ \dot_product_and_ReLU[1].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$4797(.Z({ \dot_product_and_ReLU[1].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$4798(.Z({ \dot_product_and_ReLU[1].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$4799(.Z({ \dot_product_and_ReLU[1].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$4800(.Z({ \dot_product_and_ReLU[1].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$4801(.Z({ \dot_product_and_ReLU[1].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$4802(.Z({ \dot_product_and_ReLU[1].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$4803(.Z({ \dot_product_and_ReLU[1].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$4804(.Z({ \dot_product_and_ReLU[1].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$4805(.Z({ \dot_product_and_ReLU[1].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$4806(.Z({ \dot_product_and_ReLU[1].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$4807(.Z({ \dot_product_and_ReLU[1].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$4808(.Z({ \dot_product_and_ReLU[1].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$4809(.Z({ \dot_product_and_ReLU[1].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$4810(.Z({ \dot_product_and_ReLU[1].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$4811(.Z({ \dot_product_and_ReLU[1].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$4812(.Z({ \dot_product_and_ReLU[1].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$4813(.Z({ \dot_product_and_ReLU[1].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$4814(.Z({ \dot_product_and_ReLU[1].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$4815(.Z({ \dot_product_and_ReLU[1].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$4816(.Z({ \dot_product_and_ReLU[1].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$4817(.Z({ \dot_product_and_ReLU[1].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$4818(.Z({ \dot_product_and_ReLU[1].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$4819(.Z({ \dot_product_and_ReLU[1].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$4820(.Z({ \dot_product_and_ReLU[1].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$4821(.Z({ \dot_product_and_ReLU[1].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$4822(.Z({ \dot_product_and_ReLU[1].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$4823(.Z({ \dot_product_and_ReLU[1].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$4824(.Z({ \dot_product_and_ReLU[1].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$4825(.Z({ \dot_product_and_ReLU[1].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$4826(.Z({ \dot_product_and_ReLU[1].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$4827(.Z({ \dot_product_and_ReLU[1].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$4828(.Z({ \dot_product_and_ReLU[1].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$4829(.Z({ \dot_product_and_ReLU[1].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$4830(.Z({ \dot_product_and_ReLU[1].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$4831(.Z({ \dot_product_and_ReLU[1].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$4832(.Z({ \dot_product_and_ReLU[1].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$4833(.Z({ \dot_product_and_ReLU[1].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$4834(.Z({ \dot_product_and_ReLU[1].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$4835(.Z({ \dot_product_and_ReLU[1].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$4836(.Z({ \dot_product_and_ReLU[1].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$4837(.Z({ \dot_product_and_ReLU[1].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$4838(.Z({ \dot_product_and_ReLU[1].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$4839(.Z({ \dot_product_and_ReLU[1].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$4840(.Z({ \dot_product_and_ReLU[1].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$4841(.Z({ \dot_product_and_ReLU[1].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$4842(.Z({ \dot_product_and_ReLU[1].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$4843(.Z({ \dot_product_and_ReLU[1].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$4844(.Z({ \dot_product_and_ReLU[1].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$4845(.Z({ \dot_product_and_ReLU[1].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$4846(.Z({ \dot_product_and_ReLU[1].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$4847(.Z({ \dot_product_and_ReLU[1].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$4848(.Z({ \dot_product_and_ReLU[1].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$4849(.Z({ \dot_product_and_ReLU[1].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$4850(.Z({ \dot_product_and_ReLU[1].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$4851(.Z({ \dot_product_and_ReLU[1].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$4852(.Z({ \dot_product_and_ReLU[1].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$4853(.Z({ \dot_product_and_ReLU[1].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$4854(.Z({ \dot_product_and_ReLU[1].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$4855(.Z({ \dot_product_and_ReLU[1].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$4856(.Z({ \dot_product_and_ReLU[1].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$4857(.Z({ \dot_product_and_ReLU[1].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$4858(.Z({ \dot_product_and_ReLU[1].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$4859(.Z({ \dot_product_and_ReLU[1].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$4860(.Z({ \dot_product_and_ReLU[1].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$4861(.Z({ \dot_product_and_ReLU[1].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$4862(.Z({ \dot_product_and_ReLU[1].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$4863(.Z({ \dot_product_and_ReLU[1].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$4864(.Z({ \dot_product_and_ReLU[1].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[1][255] [4:0] }), .S(B[255]));
  VDW_WMUX5 U$4865(.Z({ \dot_product_and_ReLU[0].product_terms[0] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][0] [4:0] }), .S(B[0]));
  VDW_WMUX5 U$4866(.Z({ \dot_product_and_ReLU[0].product_terms[1] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][1] [4:0] }), .S(B[1]));
  VDW_WMUX5 U$4867(.Z({ \dot_product_and_ReLU[0].product_terms[2] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][2] [4:0] }), .S(B[2]));
  VDW_WMUX5 U$4868(.Z({ \dot_product_and_ReLU[0].product_terms[3] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][3] [4:0] }), .S(B[3]));
  VDW_WMUX5 U$4869(.Z({ \dot_product_and_ReLU[0].product_terms[4] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][4] [4:0] }), .S(B[4]));
  VDW_WMUX5 U$4870(.Z({ \dot_product_and_ReLU[0].product_terms[5] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][5] [4:0] }), .S(B[5]));
  VDW_WMUX5 U$4871(.Z({ \dot_product_and_ReLU[0].product_terms[6] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][6] [4:0] }), .S(B[6]));
  VDW_WMUX5 U$4872(.Z({ \dot_product_and_ReLU[0].product_terms[7] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][7] [4:0] }), .S(B[7]));
  VDW_WMUX5 U$4873(.Z({ \dot_product_and_ReLU[0].product_terms[8] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][8] [4:0] }), .S(B[8]));
  VDW_WMUX5 U$4874(.Z({ \dot_product_and_ReLU[0].product_terms[9] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][9] [4:0] }), .S(B[9]));
  VDW_WMUX5 U$4875(.Z({ \dot_product_and_ReLU[0].product_terms[10] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][10] [4:0] }), .S(B[10]));
  VDW_WMUX5 U$4876(.Z({ \dot_product_and_ReLU[0].product_terms[11] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][11] [4:0] }), .S(B[11]));
  VDW_WMUX5 U$4877(.Z({ \dot_product_and_ReLU[0].product_terms[12] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][12] [4:0] }), .S(B[12]));
  VDW_WMUX5 U$4878(.Z({ \dot_product_and_ReLU[0].product_terms[13] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][13] [4:0] }), .S(B[13]));
  VDW_WMUX5 U$4879(.Z({ \dot_product_and_ReLU[0].product_terms[14] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][14] [4:0] }), .S(B[14]));
  VDW_WMUX5 U$4880(.Z({ \dot_product_and_ReLU[0].product_terms[15] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][15] [4:0] }), .S(B[15]));
  VDW_WMUX5 U$4881(.Z({ \dot_product_and_ReLU[0].product_terms[16] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][16] [4:0] }), .S(B[16]));
  VDW_WMUX5 U$4882(.Z({ \dot_product_and_ReLU[0].product_terms[17] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][17] [4:0] }), .S(B[17]));
  VDW_WMUX5 U$4883(.Z({ \dot_product_and_ReLU[0].product_terms[18] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][18] [4:0] }), .S(B[18]));
  VDW_WMUX5 U$4884(.Z({ \dot_product_and_ReLU[0].product_terms[19] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][19] [4:0] }), .S(B[19]));
  VDW_WMUX5 U$4885(.Z({ \dot_product_and_ReLU[0].product_terms[20] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][20] [4:0] }), .S(B[20]));
  VDW_WMUX5 U$4886(.Z({ \dot_product_and_ReLU[0].product_terms[21] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][21] [4:0] }), .S(B[21]));
  VDW_WMUX5 U$4887(.Z({ \dot_product_and_ReLU[0].product_terms[22] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][22] [4:0] }), .S(B[22]));
  VDW_WMUX5 U$4888(.Z({ \dot_product_and_ReLU[0].product_terms[23] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][23] [4:0] }), .S(B[23]));
  VDW_WMUX5 U$4889(.Z({ \dot_product_and_ReLU[0].product_terms[24] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][24] [4:0] }), .S(B[24]));
  VDW_WMUX5 U$4890(.Z({ \dot_product_and_ReLU[0].product_terms[25] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][25] [4:0] }), .S(B[25]));
  VDW_WMUX5 U$4891(.Z({ \dot_product_and_ReLU[0].product_terms[26] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][26] [4:0] }), .S(B[26]));
  VDW_WMUX5 U$4892(.Z({ \dot_product_and_ReLU[0].product_terms[27] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][27] [4:0] }), .S(B[27]));
  VDW_WMUX5 U$4893(.Z({ \dot_product_and_ReLU[0].product_terms[28] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][28] [4:0] }), .S(B[28]));
  VDW_WMUX5 U$4894(.Z({ \dot_product_and_ReLU[0].product_terms[29] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][29] [4:0] }), .S(B[29]));
  VDW_WMUX5 U$4895(.Z({ \dot_product_and_ReLU[0].product_terms[30] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][30] [4:0] }), .S(B[30]));
  VDW_WMUX5 U$4896(.Z({ \dot_product_and_ReLU[0].product_terms[31] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][31] [4:0] }), .S(B[31]));
  VDW_WMUX5 U$4897(.Z({ \dot_product_and_ReLU[0].product_terms[32] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][32] [4:0] }), .S(B[32]));
  VDW_WMUX5 U$4898(.Z({ \dot_product_and_ReLU[0].product_terms[33] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][33] [4:0] }), .S(B[33]));
  VDW_WMUX5 U$4899(.Z({ \dot_product_and_ReLU[0].product_terms[34] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][34] [4:0] }), .S(B[34]));
  VDW_WMUX5 U$4900(.Z({ \dot_product_and_ReLU[0].product_terms[35] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][35] [4:0] }), .S(B[35]));
  VDW_WMUX5 U$4901(.Z({ \dot_product_and_ReLU[0].product_terms[36] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][36] [4:0] }), .S(B[36]));
  VDW_WMUX5 U$4902(.Z({ \dot_product_and_ReLU[0].product_terms[37] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][37] [4:0] }), .S(B[37]));
  VDW_WMUX5 U$4903(.Z({ \dot_product_and_ReLU[0].product_terms[38] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][38] [4:0] }), .S(B[38]));
  VDW_WMUX5 U$4904(.Z({ \dot_product_and_ReLU[0].product_terms[39] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][39] [4:0] }), .S(B[39]));
  VDW_WMUX5 U$4905(.Z({ \dot_product_and_ReLU[0].product_terms[40] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][40] [4:0] }), .S(B[40]));
  VDW_WMUX5 U$4906(.Z({ \dot_product_and_ReLU[0].product_terms[41] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][41] [4:0] }), .S(B[41]));
  VDW_WMUX5 U$4907(.Z({ \dot_product_and_ReLU[0].product_terms[42] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][42] [4:0] }), .S(B[42]));
  VDW_WMUX5 U$4908(.Z({ \dot_product_and_ReLU[0].product_terms[43] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][43] [4:0] }), .S(B[43]));
  VDW_WMUX5 U$4909(.Z({ \dot_product_and_ReLU[0].product_terms[44] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][44] [4:0] }), .S(B[44]));
  VDW_WMUX5 U$4910(.Z({ \dot_product_and_ReLU[0].product_terms[45] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][45] [4:0] }), .S(B[45]));
  VDW_WMUX5 U$4911(.Z({ \dot_product_and_ReLU[0].product_terms[46] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][46] [4:0] }), .S(B[46]));
  VDW_WMUX5 U$4912(.Z({ \dot_product_and_ReLU[0].product_terms[47] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][47] [4:0] }), .S(B[47]));
  VDW_WMUX5 U$4913(.Z({ \dot_product_and_ReLU[0].product_terms[48] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][48] [4:0] }), .S(B[48]));
  VDW_WMUX5 U$4914(.Z({ \dot_product_and_ReLU[0].product_terms[49] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][49] [4:0] }), .S(B[49]));
  VDW_WMUX5 U$4915(.Z({ \dot_product_and_ReLU[0].product_terms[50] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][50] [4:0] }), .S(B[50]));
  VDW_WMUX5 U$4916(.Z({ \dot_product_and_ReLU[0].product_terms[51] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][51] [4:0] }), .S(B[51]));
  VDW_WMUX5 U$4917(.Z({ \dot_product_and_ReLU[0].product_terms[52] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][52] [4:0] }), .S(B[52]));
  VDW_WMUX5 U$4918(.Z({ \dot_product_and_ReLU[0].product_terms[53] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][53] [4:0] }), .S(B[53]));
  VDW_WMUX5 U$4919(.Z({ \dot_product_and_ReLU[0].product_terms[54] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][54] [4:0] }), .S(B[54]));
  VDW_WMUX5 U$4920(.Z({ \dot_product_and_ReLU[0].product_terms[55] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][55] [4:0] }), .S(B[55]));
  VDW_WMUX5 U$4921(.Z({ \dot_product_and_ReLU[0].product_terms[56] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][56] [4:0] }), .S(B[56]));
  VDW_WMUX5 U$4922(.Z({ \dot_product_and_ReLU[0].product_terms[57] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][57] [4:0] }), .S(B[57]));
  VDW_WMUX5 U$4923(.Z({ \dot_product_and_ReLU[0].product_terms[58] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][58] [4:0] }), .S(B[58]));
  VDW_WMUX5 U$4924(.Z({ \dot_product_and_ReLU[0].product_terms[59] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][59] [4:0] }), .S(B[59]));
  VDW_WMUX5 U$4925(.Z({ \dot_product_and_ReLU[0].product_terms[60] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][60] [4:0] }), .S(B[60]));
  VDW_WMUX5 U$4926(.Z({ \dot_product_and_ReLU[0].product_terms[61] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][61] [4:0] }), .S(B[61]));
  VDW_WMUX5 U$4927(.Z({ \dot_product_and_ReLU[0].product_terms[62] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][62] [4:0] }), .S(B[62]));
  VDW_WMUX5 U$4928(.Z({ \dot_product_and_ReLU[0].product_terms[63] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][63] [4:0] }), .S(B[63]));
  VDW_WMUX5 U$4929(.Z({ \dot_product_and_ReLU[0].product_terms[64] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][64] [4:0] }), .S(B[64]));
  VDW_WMUX5 U$4930(.Z({ \dot_product_and_ReLU[0].product_terms[65] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][65] [4:0] }), .S(B[65]));
  VDW_WMUX5 U$4931(.Z({ \dot_product_and_ReLU[0].product_terms[66] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][66] [4:0] }), .S(B[66]));
  VDW_WMUX5 U$4932(.Z({ \dot_product_and_ReLU[0].product_terms[67] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][67] [4:0] }), .S(B[67]));
  VDW_WMUX5 U$4933(.Z({ \dot_product_and_ReLU[0].product_terms[68] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][68] [4:0] }), .S(B[68]));
  VDW_WMUX5 U$4934(.Z({ \dot_product_and_ReLU[0].product_terms[69] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][69] [4:0] }), .S(B[69]));
  VDW_WMUX5 U$4935(.Z({ \dot_product_and_ReLU[0].product_terms[70] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][70] [4:0] }), .S(B[70]));
  VDW_WMUX5 U$4936(.Z({ \dot_product_and_ReLU[0].product_terms[71] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][71] [4:0] }), .S(B[71]));
  VDW_WMUX5 U$4937(.Z({ \dot_product_and_ReLU[0].product_terms[72] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][72] [4:0] }), .S(B[72]));
  VDW_WMUX5 U$4938(.Z({ \dot_product_and_ReLU[0].product_terms[73] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][73] [4:0] }), .S(B[73]));
  VDW_WMUX5 U$4939(.Z({ \dot_product_and_ReLU[0].product_terms[74] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][74] [4:0] }), .S(B[74]));
  VDW_WMUX5 U$4940(.Z({ \dot_product_and_ReLU[0].product_terms[75] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][75] [4:0] }), .S(B[75]));
  VDW_WMUX5 U$4941(.Z({ \dot_product_and_ReLU[0].product_terms[76] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][76] [4:0] }), .S(B[76]));
  VDW_WMUX5 U$4942(.Z({ \dot_product_and_ReLU[0].product_terms[77] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][77] [4:0] }), .S(B[77]));
  VDW_WMUX5 U$4943(.Z({ \dot_product_and_ReLU[0].product_terms[78] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][78] [4:0] }), .S(B[78]));
  VDW_WMUX5 U$4944(.Z({ \dot_product_and_ReLU[0].product_terms[79] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][79] [4:0] }), .S(B[79]));
  VDW_WMUX5 U$4945(.Z({ \dot_product_and_ReLU[0].product_terms[80] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][80] [4:0] }), .S(B[80]));
  VDW_WMUX5 U$4946(.Z({ \dot_product_and_ReLU[0].product_terms[81] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][81] [4:0] }), .S(B[81]));
  VDW_WMUX5 U$4947(.Z({ \dot_product_and_ReLU[0].product_terms[82] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][82] [4:0] }), .S(B[82]));
  VDW_WMUX5 U$4948(.Z({ \dot_product_and_ReLU[0].product_terms[83] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][83] [4:0] }), .S(B[83]));
  VDW_WMUX5 U$4949(.Z({ \dot_product_and_ReLU[0].product_terms[84] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][84] [4:0] }), .S(B[84]));
  VDW_WMUX5 U$4950(.Z({ \dot_product_and_ReLU[0].product_terms[85] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][85] [4:0] }), .S(B[85]));
  VDW_WMUX5 U$4951(.Z({ \dot_product_and_ReLU[0].product_terms[86] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][86] [4:0] }), .S(B[86]));
  VDW_WMUX5 U$4952(.Z({ \dot_product_and_ReLU[0].product_terms[87] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][87] [4:0] }), .S(B[87]));
  VDW_WMUX5 U$4953(.Z({ \dot_product_and_ReLU[0].product_terms[88] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][88] [4:0] }), .S(B[88]));
  VDW_WMUX5 U$4954(.Z({ \dot_product_and_ReLU[0].product_terms[89] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][89] [4:0] }), .S(B[89]));
  VDW_WMUX5 U$4955(.Z({ \dot_product_and_ReLU[0].product_terms[90] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][90] [4:0] }), .S(B[90]));
  VDW_WMUX5 U$4956(.Z({ \dot_product_and_ReLU[0].product_terms[91] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][91] [4:0] }), .S(B[91]));
  VDW_WMUX5 U$4957(.Z({ \dot_product_and_ReLU[0].product_terms[92] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][92] [4:0] }), .S(B[92]));
  VDW_WMUX5 U$4958(.Z({ \dot_product_and_ReLU[0].product_terms[93] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][93] [4:0] }), .S(B[93]));
  VDW_WMUX5 U$4959(.Z({ \dot_product_and_ReLU[0].product_terms[94] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][94] [4:0] }), .S(B[94]));
  VDW_WMUX5 U$4960(.Z({ \dot_product_and_ReLU[0].product_terms[95] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][95] [4:0] }), .S(B[95]));
  VDW_WMUX5 U$4961(.Z({ \dot_product_and_ReLU[0].product_terms[96] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][96] [4:0] }), .S(B[96]));
  VDW_WMUX5 U$4962(.Z({ \dot_product_and_ReLU[0].product_terms[97] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][97] [4:0] }), .S(B[97]));
  VDW_WMUX5 U$4963(.Z({ \dot_product_and_ReLU[0].product_terms[98] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][98] [4:0] }), .S(B[98]));
  VDW_WMUX5 U$4964(.Z({ \dot_product_and_ReLU[0].product_terms[99] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][99] [4:0] }), .S(B[99]));
  VDW_WMUX5 U$4965(.Z({ \dot_product_and_ReLU[0].product_terms[100] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][100] [4:0] }), .S(B[100]));
  VDW_WMUX5 U$4966(.Z({ \dot_product_and_ReLU[0].product_terms[101] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][101] [4:0] }), .S(B[101]));
  VDW_WMUX5 U$4967(.Z({ \dot_product_and_ReLU[0].product_terms[102] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][102] [4:0] }), .S(B[102]));
  VDW_WMUX5 U$4968(.Z({ \dot_product_and_ReLU[0].product_terms[103] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][103] [4:0] }), .S(B[103]));
  VDW_WMUX5 U$4969(.Z({ \dot_product_and_ReLU[0].product_terms[104] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][104] [4:0] }), .S(B[104]));
  VDW_WMUX5 U$4970(.Z({ \dot_product_and_ReLU[0].product_terms[105] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][105] [4:0] }), .S(B[105]));
  VDW_WMUX5 U$4971(.Z({ \dot_product_and_ReLU[0].product_terms[106] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][106] [4:0] }), .S(B[106]));
  VDW_WMUX5 U$4972(.Z({ \dot_product_and_ReLU[0].product_terms[107] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][107] [4:0] }), .S(B[107]));
  VDW_WMUX5 U$4973(.Z({ \dot_product_and_ReLU[0].product_terms[108] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][108] [4:0] }), .S(B[108]));
  VDW_WMUX5 U$4974(.Z({ \dot_product_and_ReLU[0].product_terms[109] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][109] [4:0] }), .S(B[109]));
  VDW_WMUX5 U$4975(.Z({ \dot_product_and_ReLU[0].product_terms[110] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][110] [4:0] }), .S(B[110]));
  VDW_WMUX5 U$4976(.Z({ \dot_product_and_ReLU[0].product_terms[111] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][111] [4:0] }), .S(B[111]));
  VDW_WMUX5 U$4977(.Z({ \dot_product_and_ReLU[0].product_terms[112] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][112] [4:0] }), .S(B[112]));
  VDW_WMUX5 U$4978(.Z({ \dot_product_and_ReLU[0].product_terms[113] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][113] [4:0] }), .S(B[113]));
  VDW_WMUX5 U$4979(.Z({ \dot_product_and_ReLU[0].product_terms[114] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][114] [4:0] }), .S(B[114]));
  VDW_WMUX5 U$4980(.Z({ \dot_product_and_ReLU[0].product_terms[115] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][115] [4:0] }), .S(B[115]));
  VDW_WMUX5 U$4981(.Z({ \dot_product_and_ReLU[0].product_terms[116] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][116] [4:0] }), .S(B[116]));
  VDW_WMUX5 U$4982(.Z({ \dot_product_and_ReLU[0].product_terms[117] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][117] [4:0] }), .S(B[117]));
  VDW_WMUX5 U$4983(.Z({ \dot_product_and_ReLU[0].product_terms[118] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][118] [4:0] }), .S(B[118]));
  VDW_WMUX5 U$4984(.Z({ \dot_product_and_ReLU[0].product_terms[119] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][119] [4:0] }), .S(B[119]));
  VDW_WMUX5 U$4985(.Z({ \dot_product_and_ReLU[0].product_terms[120] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][120] [4:0] }), .S(B[120]));
  VDW_WMUX5 U$4986(.Z({ \dot_product_and_ReLU[0].product_terms[121] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][121] [4:0] }), .S(B[121]));
  VDW_WMUX5 U$4987(.Z({ \dot_product_and_ReLU[0].product_terms[122] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][122] [4:0] }), .S(B[122]));
  VDW_WMUX5 U$4988(.Z({ \dot_product_and_ReLU[0].product_terms[123] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][123] [4:0] }), .S(B[123]));
  VDW_WMUX5 U$4989(.Z({ \dot_product_and_ReLU[0].product_terms[124] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][124] [4:0] }), .S(B[124]));
  VDW_WMUX5 U$4990(.Z({ \dot_product_and_ReLU[0].product_terms[125] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][125] [4:0] }), .S(B[125]));
  VDW_WMUX5 U$4991(.Z({ \dot_product_and_ReLU[0].product_terms[126] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][126] [4:0] }), .S(B[126]));
  VDW_WMUX5 U$4992(.Z({ \dot_product_and_ReLU[0].product_terms[127] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][127] [4:0] }), .S(B[127]));
  VDW_WMUX5 U$4993(.Z({ \dot_product_and_ReLU[0].product_terms[128] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][128] [4:0] }), .S(B[128]));
  VDW_WMUX5 U$4994(.Z({ \dot_product_and_ReLU[0].product_terms[129] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][129] [4:0] }), .S(B[129]));
  VDW_WMUX5 U$4995(.Z({ \dot_product_and_ReLU[0].product_terms[130] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][130] [4:0] }), .S(B[130]));
  VDW_WMUX5 U$4996(.Z({ \dot_product_and_ReLU[0].product_terms[131] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][131] [4:0] }), .S(B[131]));
  VDW_WMUX5 U$4997(.Z({ \dot_product_and_ReLU[0].product_terms[132] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][132] [4:0] }), .S(B[132]));
  VDW_WMUX5 U$4998(.Z({ \dot_product_and_ReLU[0].product_terms[133] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][133] [4:0] }), .S(B[133]));
  VDW_WMUX5 U$4999(.Z({ \dot_product_and_ReLU[0].product_terms[134] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][134] [4:0] }), .S(B[134]));
  VDW_WMUX5 U$5000(.Z({ \dot_product_and_ReLU[0].product_terms[135] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][135] [4:0] }), .S(B[135]));
  VDW_WMUX5 U$5001(.Z({ \dot_product_and_ReLU[0].product_terms[136] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][136] [4:0] }), .S(B[136]));
  VDW_WMUX5 U$5002(.Z({ \dot_product_and_ReLU[0].product_terms[137] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][137] [4:0] }), .S(B[137]));
  VDW_WMUX5 U$5003(.Z({ \dot_product_and_ReLU[0].product_terms[138] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][138] [4:0] }), .S(B[138]));
  VDW_WMUX5 U$5004(.Z({ \dot_product_and_ReLU[0].product_terms[139] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][139] [4:0] }), .S(B[139]));
  VDW_WMUX5 U$5005(.Z({ \dot_product_and_ReLU[0].product_terms[140] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][140] [4:0] }), .S(B[140]));
  VDW_WMUX5 U$5006(.Z({ \dot_product_and_ReLU[0].product_terms[141] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][141] [4:0] }), .S(B[141]));
  VDW_WMUX5 U$5007(.Z({ \dot_product_and_ReLU[0].product_terms[142] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][142] [4:0] }), .S(B[142]));
  VDW_WMUX5 U$5008(.Z({ \dot_product_and_ReLU[0].product_terms[143] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][143] [4:0] }), .S(B[143]));
  VDW_WMUX5 U$5009(.Z({ \dot_product_and_ReLU[0].product_terms[144] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][144] [4:0] }), .S(B[144]));
  VDW_WMUX5 U$5010(.Z({ \dot_product_and_ReLU[0].product_terms[145] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][145] [4:0] }), .S(B[145]));
  VDW_WMUX5 U$5011(.Z({ \dot_product_and_ReLU[0].product_terms[146] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][146] [4:0] }), .S(B[146]));
  VDW_WMUX5 U$5012(.Z({ \dot_product_and_ReLU[0].product_terms[147] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][147] [4:0] }), .S(B[147]));
  VDW_WMUX5 U$5013(.Z({ \dot_product_and_ReLU[0].product_terms[148] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][148] [4:0] }), .S(B[148]));
  VDW_WMUX5 U$5014(.Z({ \dot_product_and_ReLU[0].product_terms[149] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][149] [4:0] }), .S(B[149]));
  VDW_WMUX5 U$5015(.Z({ \dot_product_and_ReLU[0].product_terms[150] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][150] [4:0] }), .S(B[150]));
  VDW_WMUX5 U$5016(.Z({ \dot_product_and_ReLU[0].product_terms[151] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][151] [4:0] }), .S(B[151]));
  VDW_WMUX5 U$5017(.Z({ \dot_product_and_ReLU[0].product_terms[152] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][152] [4:0] }), .S(B[152]));
  VDW_WMUX5 U$5018(.Z({ \dot_product_and_ReLU[0].product_terms[153] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][153] [4:0] }), .S(B[153]));
  VDW_WMUX5 U$5019(.Z({ \dot_product_and_ReLU[0].product_terms[154] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][154] [4:0] }), .S(B[154]));
  VDW_WMUX5 U$5020(.Z({ \dot_product_and_ReLU[0].product_terms[155] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][155] [4:0] }), .S(B[155]));
  VDW_WMUX5 U$5021(.Z({ \dot_product_and_ReLU[0].product_terms[156] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][156] [4:0] }), .S(B[156]));
  VDW_WMUX5 U$5022(.Z({ \dot_product_and_ReLU[0].product_terms[157] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][157] [4:0] }), .S(B[157]));
  VDW_WMUX5 U$5023(.Z({ \dot_product_and_ReLU[0].product_terms[158] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][158] [4:0] }), .S(B[158]));
  VDW_WMUX5 U$5024(.Z({ \dot_product_and_ReLU[0].product_terms[159] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][159] [4:0] }), .S(B[159]));
  VDW_WMUX5 U$5025(.Z({ \dot_product_and_ReLU[0].product_terms[160] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][160] [4:0] }), .S(B[160]));
  VDW_WMUX5 U$5026(.Z({ \dot_product_and_ReLU[0].product_terms[161] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][161] [4:0] }), .S(B[161]));
  VDW_WMUX5 U$5027(.Z({ \dot_product_and_ReLU[0].product_terms[162] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][162] [4:0] }), .S(B[162]));
  VDW_WMUX5 U$5028(.Z({ \dot_product_and_ReLU[0].product_terms[163] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][163] [4:0] }), .S(B[163]));
  VDW_WMUX5 U$5029(.Z({ \dot_product_and_ReLU[0].product_terms[164] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][164] [4:0] }), .S(B[164]));
  VDW_WMUX5 U$5030(.Z({ \dot_product_and_ReLU[0].product_terms[165] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][165] [4:0] }), .S(B[165]));
  VDW_WMUX5 U$5031(.Z({ \dot_product_and_ReLU[0].product_terms[166] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][166] [4:0] }), .S(B[166]));
  VDW_WMUX5 U$5032(.Z({ \dot_product_and_ReLU[0].product_terms[167] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][167] [4:0] }), .S(B[167]));
  VDW_WMUX5 U$5033(.Z({ \dot_product_and_ReLU[0].product_terms[168] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][168] [4:0] }), .S(B[168]));
  VDW_WMUX5 U$5034(.Z({ \dot_product_and_ReLU[0].product_terms[169] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][169] [4:0] }), .S(B[169]));
  VDW_WMUX5 U$5035(.Z({ \dot_product_and_ReLU[0].product_terms[170] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][170] [4:0] }), .S(B[170]));
  VDW_WMUX5 U$5036(.Z({ \dot_product_and_ReLU[0].product_terms[171] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][171] [4:0] }), .S(B[171]));
  VDW_WMUX5 U$5037(.Z({ \dot_product_and_ReLU[0].product_terms[172] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][172] [4:0] }), .S(B[172]));
  VDW_WMUX5 U$5038(.Z({ \dot_product_and_ReLU[0].product_terms[173] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][173] [4:0] }), .S(B[173]));
  VDW_WMUX5 U$5039(.Z({ \dot_product_and_ReLU[0].product_terms[174] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][174] [4:0] }), .S(B[174]));
  VDW_WMUX5 U$5040(.Z({ \dot_product_and_ReLU[0].product_terms[175] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][175] [4:0] }), .S(B[175]));
  VDW_WMUX5 U$5041(.Z({ \dot_product_and_ReLU[0].product_terms[176] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][176] [4:0] }), .S(B[176]));
  VDW_WMUX5 U$5042(.Z({ \dot_product_and_ReLU[0].product_terms[177] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][177] [4:0] }), .S(B[177]));
  VDW_WMUX5 U$5043(.Z({ \dot_product_and_ReLU[0].product_terms[178] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][178] [4:0] }), .S(B[178]));
  VDW_WMUX5 U$5044(.Z({ \dot_product_and_ReLU[0].product_terms[179] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][179] [4:0] }), .S(B[179]));
  VDW_WMUX5 U$5045(.Z({ \dot_product_and_ReLU[0].product_terms[180] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][180] [4:0] }), .S(B[180]));
  VDW_WMUX5 U$5046(.Z({ \dot_product_and_ReLU[0].product_terms[181] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][181] [4:0] }), .S(B[181]));
  VDW_WMUX5 U$5047(.Z({ \dot_product_and_ReLU[0].product_terms[182] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][182] [4:0] }), .S(B[182]));
  VDW_WMUX5 U$5048(.Z({ \dot_product_and_ReLU[0].product_terms[183] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][183] [4:0] }), .S(B[183]));
  VDW_WMUX5 U$5049(.Z({ \dot_product_and_ReLU[0].product_terms[184] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][184] [4:0] }), .S(B[184]));
  VDW_WMUX5 U$5050(.Z({ \dot_product_and_ReLU[0].product_terms[185] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][185] [4:0] }), .S(B[185]));
  VDW_WMUX5 U$5051(.Z({ \dot_product_and_ReLU[0].product_terms[186] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][186] [4:0] }), .S(B[186]));
  VDW_WMUX5 U$5052(.Z({ \dot_product_and_ReLU[0].product_terms[187] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][187] [4:0] }), .S(B[187]));
  VDW_WMUX5 U$5053(.Z({ \dot_product_and_ReLU[0].product_terms[188] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][188] [4:0] }), .S(B[188]));
  VDW_WMUX5 U$5054(.Z({ \dot_product_and_ReLU[0].product_terms[189] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][189] [4:0] }), .S(B[189]));
  VDW_WMUX5 U$5055(.Z({ \dot_product_and_ReLU[0].product_terms[190] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][190] [4:0] }), .S(B[190]));
  VDW_WMUX5 U$5056(.Z({ \dot_product_and_ReLU[0].product_terms[191] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][191] [4:0] }), .S(B[191]));
  VDW_WMUX5 U$5057(.Z({ \dot_product_and_ReLU[0].product_terms[192] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][192] [4:0] }), .S(B[192]));
  VDW_WMUX5 U$5058(.Z({ \dot_product_and_ReLU[0].product_terms[193] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][193] [4:0] }), .S(B[193]));
  VDW_WMUX5 U$5059(.Z({ \dot_product_and_ReLU[0].product_terms[194] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][194] [4:0] }), .S(B[194]));
  VDW_WMUX5 U$5060(.Z({ \dot_product_and_ReLU[0].product_terms[195] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][195] [4:0] }), .S(B[195]));
  VDW_WMUX5 U$5061(.Z({ \dot_product_and_ReLU[0].product_terms[196] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][196] [4:0] }), .S(B[196]));
  VDW_WMUX5 U$5062(.Z({ \dot_product_and_ReLU[0].product_terms[197] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][197] [4:0] }), .S(B[197]));
  VDW_WMUX5 U$5063(.Z({ \dot_product_and_ReLU[0].product_terms[198] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][198] [4:0] }), .S(B[198]));
  VDW_WMUX5 U$5064(.Z({ \dot_product_and_ReLU[0].product_terms[199] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][199] [4:0] }), .S(B[199]));
  VDW_WMUX5 U$5065(.Z({ \dot_product_and_ReLU[0].product_terms[200] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][200] [4:0] }), .S(B[200]));
  VDW_WMUX5 U$5066(.Z({ \dot_product_and_ReLU[0].product_terms[201] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][201] [4:0] }), .S(B[201]));
  VDW_WMUX5 U$5067(.Z({ \dot_product_and_ReLU[0].product_terms[202] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][202] [4:0] }), .S(B[202]));
  VDW_WMUX5 U$5068(.Z({ \dot_product_and_ReLU[0].product_terms[203] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][203] [4:0] }), .S(B[203]));
  VDW_WMUX5 U$5069(.Z({ \dot_product_and_ReLU[0].product_terms[204] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][204] [4:0] }), .S(B[204]));
  VDW_WMUX5 U$5070(.Z({ \dot_product_and_ReLU[0].product_terms[205] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][205] [4:0] }), .S(B[205]));
  VDW_WMUX5 U$5071(.Z({ \dot_product_and_ReLU[0].product_terms[206] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][206] [4:0] }), .S(B[206]));
  VDW_WMUX5 U$5072(.Z({ \dot_product_and_ReLU[0].product_terms[207] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][207] [4:0] }), .S(B[207]));
  VDW_WMUX5 U$5073(.Z({ \dot_product_and_ReLU[0].product_terms[208] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][208] [4:0] }), .S(B[208]));
  VDW_WMUX5 U$5074(.Z({ \dot_product_and_ReLU[0].product_terms[209] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][209] [4:0] }), .S(B[209]));
  VDW_WMUX5 U$5075(.Z({ \dot_product_and_ReLU[0].product_terms[210] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][210] [4:0] }), .S(B[210]));
  VDW_WMUX5 U$5076(.Z({ \dot_product_and_ReLU[0].product_terms[211] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][211] [4:0] }), .S(B[211]));
  VDW_WMUX5 U$5077(.Z({ \dot_product_and_ReLU[0].product_terms[212] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][212] [4:0] }), .S(B[212]));
  VDW_WMUX5 U$5078(.Z({ \dot_product_and_ReLU[0].product_terms[213] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][213] [4:0] }), .S(B[213]));
  VDW_WMUX5 U$5079(.Z({ \dot_product_and_ReLU[0].product_terms[214] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][214] [4:0] }), .S(B[214]));
  VDW_WMUX5 U$5080(.Z({ \dot_product_and_ReLU[0].product_terms[215] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][215] [4:0] }), .S(B[215]));
  VDW_WMUX5 U$5081(.Z({ \dot_product_and_ReLU[0].product_terms[216] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][216] [4:0] }), .S(B[216]));
  VDW_WMUX5 U$5082(.Z({ \dot_product_and_ReLU[0].product_terms[217] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][217] [4:0] }), .S(B[217]));
  VDW_WMUX5 U$5083(.Z({ \dot_product_and_ReLU[0].product_terms[218] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][218] [4:0] }), .S(B[218]));
  VDW_WMUX5 U$5084(.Z({ \dot_product_and_ReLU[0].product_terms[219] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][219] [4:0] }), .S(B[219]));
  VDW_WMUX5 U$5085(.Z({ \dot_product_and_ReLU[0].product_terms[220] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][220] [4:0] }), .S(B[220]));
  VDW_WMUX5 U$5086(.Z({ \dot_product_and_ReLU[0].product_terms[221] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][221] [4:0] }), .S(B[221]));
  VDW_WMUX5 U$5087(.Z({ \dot_product_and_ReLU[0].product_terms[222] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][222] [4:0] }), .S(B[222]));
  VDW_WMUX5 U$5088(.Z({ \dot_product_and_ReLU[0].product_terms[223] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][223] [4:0] }), .S(B[223]));
  VDW_WMUX5 U$5089(.Z({ \dot_product_and_ReLU[0].product_terms[224] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][224] [4:0] }), .S(B[224]));
  VDW_WMUX5 U$5090(.Z({ \dot_product_and_ReLU[0].product_terms[225] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][225] [4:0] }), .S(B[225]));
  VDW_WMUX5 U$5091(.Z({ \dot_product_and_ReLU[0].product_terms[226] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][226] [4:0] }), .S(B[226]));
  VDW_WMUX5 U$5092(.Z({ \dot_product_and_ReLU[0].product_terms[227] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][227] [4:0] }), .S(B[227]));
  VDW_WMUX5 U$5093(.Z({ \dot_product_and_ReLU[0].product_terms[228] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][228] [4:0] }), .S(B[228]));
  VDW_WMUX5 U$5094(.Z({ \dot_product_and_ReLU[0].product_terms[229] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][229] [4:0] }), .S(B[229]));
  VDW_WMUX5 U$5095(.Z({ \dot_product_and_ReLU[0].product_terms[230] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][230] [4:0] }), .S(B[230]));
  VDW_WMUX5 U$5096(.Z({ \dot_product_and_ReLU[0].product_terms[231] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][231] [4:0] }), .S(B[231]));
  VDW_WMUX5 U$5097(.Z({ \dot_product_and_ReLU[0].product_terms[232] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][232] [4:0] }), .S(B[232]));
  VDW_WMUX5 U$5098(.Z({ \dot_product_and_ReLU[0].product_terms[233] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][233] [4:0] }), .S(B[233]));
  VDW_WMUX5 U$5099(.Z({ \dot_product_and_ReLU[0].product_terms[234] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][234] [4:0] }), .S(B[234]));
  VDW_WMUX5 U$5100(.Z({ \dot_product_and_ReLU[0].product_terms[235] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][235] [4:0] }), .S(B[235]));
  VDW_WMUX5 U$5101(.Z({ \dot_product_and_ReLU[0].product_terms[236] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][236] [4:0] }), .S(B[236]));
  VDW_WMUX5 U$5102(.Z({ \dot_product_and_ReLU[0].product_terms[237] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][237] [4:0] }), .S(B[237]));
  VDW_WMUX5 U$5103(.Z({ \dot_product_and_ReLU[0].product_terms[238] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][238] [4:0] }), .S(B[238]));
  VDW_WMUX5 U$5104(.Z({ \dot_product_and_ReLU[0].product_terms[239] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][239] [4:0] }), .S(B[239]));
  VDW_WMUX5 U$5105(.Z({ \dot_product_and_ReLU[0].product_terms[240] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][240] [4:0] }), .S(B[240]));
  VDW_WMUX5 U$5106(.Z({ \dot_product_and_ReLU[0].product_terms[241] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][241] [4:0] }), .S(B[241]));
  VDW_WMUX5 U$5107(.Z({ \dot_product_and_ReLU[0].product_terms[242] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][242] [4:0] }), .S(B[242]));
  VDW_WMUX5 U$5108(.Z({ \dot_product_and_ReLU[0].product_terms[243] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][243] [4:0] }), .S(B[243]));
  VDW_WMUX5 U$5109(.Z({ \dot_product_and_ReLU[0].product_terms[244] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][244] [4:0] }), .S(B[244]));
  VDW_WMUX5 U$5110(.Z({ \dot_product_and_ReLU[0].product_terms[245] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][245] [4:0] }), .S(B[245]));
  VDW_WMUX5 U$5111(.Z({ \dot_product_and_ReLU[0].product_terms[246] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][246] [4:0] }), .S(B[246]));
  VDW_WMUX5 U$5112(.Z({ \dot_product_and_ReLU[0].product_terms[247] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][247] [4:0] }), .S(B[247]));
  VDW_WMUX5 U$5113(.Z({ \dot_product_and_ReLU[0].product_terms[248] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][248] [4:0] }), .S(B[248]));
  VDW_WMUX5 U$5114(.Z({ \dot_product_and_ReLU[0].product_terms[249] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][249] [4:0] }), .S(B[249]));
  VDW_WMUX5 U$5115(.Z({ \dot_product_and_ReLU[0].product_terms[250] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][250] [4:0] }), .S(B[250]));
  VDW_WMUX5 U$5116(.Z({ \dot_product_and_ReLU[0].product_terms[251] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][251] [4:0] }), .S(B[251]));
  VDW_WMUX5 U$5117(.Z({ \dot_product_and_ReLU[0].product_terms[252] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][252] [4:0] }), .S(B[252]));
  VDW_WMUX5 U$5118(.Z({ \dot_product_and_ReLU[0].product_terms[253] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][253] [4:0] }), .S(B[253]));
  VDW_WMUX5 U$5119(.Z({ \dot_product_and_ReLU[0].product_terms[254] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][254] [4:0] }), .S(B[254]));
  VDW_WMUX5 U$5120(.Z({ \dot_product_and_ReLU[0].product_terms[255] [4:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ \A[0][255] [4:0] }), .S(B[255]));
  _HDFF_verplex \out_reg_reg[0][8] (.Q(\out_reg[0] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[0] [8]));
  _HDFF_verplex \out_reg_reg[0][7] (.Q(\out_reg[0] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[0] [7]));
  _HDFF_verplex \out_reg_reg[0][6] (.Q(\out_reg[0] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[0] [6]));
  _HDFF_verplex \out_reg_reg[0][5] (.Q(\out_reg[0] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[0] [5]));
  _HDFF_verplex \out_reg_reg[0][4] (.Q(\out_reg[0] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[0] [4]));
  _HDFF_verplex \out_reg_reg[0][3] (.Q(\out_reg[0] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[0] [3]));
  _HDFF_verplex \out_reg_reg[0][2] (.Q(\out_reg[0] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[0] [2]));
  _HDFF_verplex \out_reg_reg[0][1] (.Q(\out_reg[0] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[0] [1]));
  _HDFF_verplex \out_reg_reg[0][0] (.Q(\out_reg[0] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[0] [0]));
  _HDFF_verplex \out_reg_reg[1][8] (.Q(\out_reg[1] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[1] [8]));
  _HDFF_verplex \out_reg_reg[1][7] (.Q(\out_reg[1] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[1] [7]));
  _HDFF_verplex \out_reg_reg[1][6] (.Q(\out_reg[1] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[1] [6]));
  _HDFF_verplex \out_reg_reg[1][5] (.Q(\out_reg[1] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[1] [5]));
  _HDFF_verplex \out_reg_reg[1][4] (.Q(\out_reg[1] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[1] [4]));
  _HDFF_verplex \out_reg_reg[1][3] (.Q(\out_reg[1] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[1] [3]));
  _HDFF_verplex \out_reg_reg[1][2] (.Q(\out_reg[1] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[1] [2]));
  _HDFF_verplex \out_reg_reg[1][1] (.Q(\out_reg[1] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[1] [1]));
  _HDFF_verplex \out_reg_reg[1][0] (.Q(\out_reg[1] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[1] [0]));
  _HDFF_verplex \out_reg_reg[2][8] (.Q(\out_reg[2] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[2] [8]));
  _HDFF_verplex \out_reg_reg[2][7] (.Q(\out_reg[2] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[2] [7]));
  _HDFF_verplex \out_reg_reg[2][6] (.Q(\out_reg[2] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[2] [6]));
  _HDFF_verplex \out_reg_reg[2][5] (.Q(\out_reg[2] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[2] [5]));
  _HDFF_verplex \out_reg_reg[2][4] (.Q(\out_reg[2] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[2] [4]));
  _HDFF_verplex \out_reg_reg[2][3] (.Q(\out_reg[2] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[2] [3]));
  _HDFF_verplex \out_reg_reg[2][2] (.Q(\out_reg[2] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[2] [2]));
  _HDFF_verplex \out_reg_reg[2][1] (.Q(\out_reg[2] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[2] [1]));
  _HDFF_verplex \out_reg_reg[2][0] (.Q(\out_reg[2] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[2] [0]));
  _HDFF_verplex \out_reg_reg[3][8] (.Q(\out_reg[3] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[3] [8]));
  _HDFF_verplex \out_reg_reg[3][7] (.Q(\out_reg[3] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[3] [7]));
  _HDFF_verplex \out_reg_reg[3][6] (.Q(\out_reg[3] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[3] [6]));
  _HDFF_verplex \out_reg_reg[3][5] (.Q(\out_reg[3] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[3] [5]));
  _HDFF_verplex \out_reg_reg[3][4] (.Q(\out_reg[3] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[3] [4]));
  _HDFF_verplex \out_reg_reg[3][3] (.Q(\out_reg[3] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[3] [3]));
  _HDFF_verplex \out_reg_reg[3][2] (.Q(\out_reg[3] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[3] [2]));
  _HDFF_verplex \out_reg_reg[3][1] (.Q(\out_reg[3] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[3] [1]));
  _HDFF_verplex \out_reg_reg[3][0] (.Q(\out_reg[3] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[3] [0]));
  _HDFF_verplex \out_reg_reg[4][8] (.Q(\out_reg[4] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[4] [8]));
  _HDFF_verplex \out_reg_reg[4][7] (.Q(\out_reg[4] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[4] [7]));
  _HDFF_verplex \out_reg_reg[4][6] (.Q(\out_reg[4] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[4] [6]));
  _HDFF_verplex \out_reg_reg[4][5] (.Q(\out_reg[4] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[4] [5]));
  _HDFF_verplex \out_reg_reg[4][4] (.Q(\out_reg[4] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[4] [4]));
  _HDFF_verplex \out_reg_reg[4][3] (.Q(\out_reg[4] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[4] [3]));
  _HDFF_verplex \out_reg_reg[4][2] (.Q(\out_reg[4] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[4] [2]));
  _HDFF_verplex \out_reg_reg[4][1] (.Q(\out_reg[4] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[4] [1]));
  _HDFF_verplex \out_reg_reg[4][0] (.Q(\out_reg[4] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[4] [0]));
  _HDFF_verplex \out_reg_reg[5][8] (.Q(\out_reg[5] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[5] [8]));
  _HDFF_verplex \out_reg_reg[5][7] (.Q(\out_reg[5] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[5] [7]));
  _HDFF_verplex \out_reg_reg[5][6] (.Q(\out_reg[5] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[5] [6]));
  _HDFF_verplex \out_reg_reg[5][5] (.Q(\out_reg[5] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[5] [5]));
  _HDFF_verplex \out_reg_reg[5][4] (.Q(\out_reg[5] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[5] [4]));
  _HDFF_verplex \out_reg_reg[5][3] (.Q(\out_reg[5] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[5] [3]));
  _HDFF_verplex \out_reg_reg[5][2] (.Q(\out_reg[5] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[5] [2]));
  _HDFF_verplex \out_reg_reg[5][1] (.Q(\out_reg[5] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[5] [1]));
  _HDFF_verplex \out_reg_reg[5][0] (.Q(\out_reg[5] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[5] [0]));
  _HDFF_verplex \out_reg_reg[6][8] (.Q(\out_reg[6] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[6] [8]));
  _HDFF_verplex \out_reg_reg[6][7] (.Q(\out_reg[6] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[6] [7]));
  _HDFF_verplex \out_reg_reg[6][6] (.Q(\out_reg[6] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[6] [6]));
  _HDFF_verplex \out_reg_reg[6][5] (.Q(\out_reg[6] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[6] [5]));
  _HDFF_verplex \out_reg_reg[6][4] (.Q(\out_reg[6] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[6] [4]));
  _HDFF_verplex \out_reg_reg[6][3] (.Q(\out_reg[6] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[6] [3]));
  _HDFF_verplex \out_reg_reg[6][2] (.Q(\out_reg[6] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[6] [2]));
  _HDFF_verplex \out_reg_reg[6][1] (.Q(\out_reg[6] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[6] [1]));
  _HDFF_verplex \out_reg_reg[6][0] (.Q(\out_reg[6] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[6] [0]));
  _HDFF_verplex \out_reg_reg[7][8] (.Q(\out_reg[7] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[7] [8]));
  _HDFF_verplex \out_reg_reg[7][7] (.Q(\out_reg[7] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[7] [7]));
  _HDFF_verplex \out_reg_reg[7][6] (.Q(\out_reg[7] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[7] [6]));
  _HDFF_verplex \out_reg_reg[7][5] (.Q(\out_reg[7] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[7] [5]));
  _HDFF_verplex \out_reg_reg[7][4] (.Q(\out_reg[7] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[7] [4]));
  _HDFF_verplex \out_reg_reg[7][3] (.Q(\out_reg[7] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[7] [3]));
  _HDFF_verplex \out_reg_reg[7][2] (.Q(\out_reg[7] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[7] [2]));
  _HDFF_verplex \out_reg_reg[7][1] (.Q(\out_reg[7] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[7] [1]));
  _HDFF_verplex \out_reg_reg[7][0] (.Q(\out_reg[7] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[7] [0]));
  _HDFF_verplex \out_reg_reg[8][8] (.Q(\out_reg[8] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[8] [8]));
  _HDFF_verplex \out_reg_reg[8][7] (.Q(\out_reg[8] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[8] [7]));
  _HDFF_verplex \out_reg_reg[8][6] (.Q(\out_reg[8] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[8] [6]));
  _HDFF_verplex \out_reg_reg[8][5] (.Q(\out_reg[8] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[8] [5]));
  _HDFF_verplex \out_reg_reg[8][4] (.Q(\out_reg[8] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[8] [4]));
  _HDFF_verplex \out_reg_reg[8][3] (.Q(\out_reg[8] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[8] [3]));
  _HDFF_verplex \out_reg_reg[8][2] (.Q(\out_reg[8] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[8] [2]));
  _HDFF_verplex \out_reg_reg[8][1] (.Q(\out_reg[8] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[8] [1]));
  _HDFF_verplex \out_reg_reg[8][0] (.Q(\out_reg[8] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[8] [0]));
  _HDFF_verplex \out_reg_reg[9][8] (.Q(\out_reg[9] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[9] [8]));
  _HDFF_verplex \out_reg_reg[9][7] (.Q(\out_reg[9] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[9] [7]));
  _HDFF_verplex \out_reg_reg[9][6] (.Q(\out_reg[9] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[9] [6]));
  _HDFF_verplex \out_reg_reg[9][5] (.Q(\out_reg[9] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[9] [5]));
  _HDFF_verplex \out_reg_reg[9][4] (.Q(\out_reg[9] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[9] [4]));
  _HDFF_verplex \out_reg_reg[9][3] (.Q(\out_reg[9] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[9] [3]));
  _HDFF_verplex \out_reg_reg[9][2] (.Q(\out_reg[9] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[9] [2]));
  _HDFF_verplex \out_reg_reg[9][1] (.Q(\out_reg[9] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[9] [1]));
  _HDFF_verplex \out_reg_reg[9][0] (.Q(\out_reg[9] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[9] [0]));
  _HDFF_verplex \out_reg_reg[10][8] (.Q(\out_reg[10] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[10] [8]));
  _HDFF_verplex \out_reg_reg[10][7] (.Q(\out_reg[10] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[10] [7]));
  _HDFF_verplex \out_reg_reg[10][6] (.Q(\out_reg[10] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[10] [6]));
  _HDFF_verplex \out_reg_reg[10][5] (.Q(\out_reg[10] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[10] [5]));
  _HDFF_verplex \out_reg_reg[10][4] (.Q(\out_reg[10] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[10] [4]));
  _HDFF_verplex \out_reg_reg[10][3] (.Q(\out_reg[10] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[10] [3]));
  _HDFF_verplex \out_reg_reg[10][2] (.Q(\out_reg[10] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[10] [2]));
  _HDFF_verplex \out_reg_reg[10][1] (.Q(\out_reg[10] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[10] [1]));
  _HDFF_verplex \out_reg_reg[10][0] (.Q(\out_reg[10] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[10] [0]));
  _HDFF_verplex \out_reg_reg[11][8] (.Q(\out_reg[11] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[11] [8]));
  _HDFF_verplex \out_reg_reg[11][7] (.Q(\out_reg[11] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[11] [7]));
  _HDFF_verplex \out_reg_reg[11][6] (.Q(\out_reg[11] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[11] [6]));
  _HDFF_verplex \out_reg_reg[11][5] (.Q(\out_reg[11] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[11] [5]));
  _HDFF_verplex \out_reg_reg[11][4] (.Q(\out_reg[11] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[11] [4]));
  _HDFF_verplex \out_reg_reg[11][3] (.Q(\out_reg[11] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[11] [3]));
  _HDFF_verplex \out_reg_reg[11][2] (.Q(\out_reg[11] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[11] [2]));
  _HDFF_verplex \out_reg_reg[11][1] (.Q(\out_reg[11] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[11] [1]));
  _HDFF_verplex \out_reg_reg[11][0] (.Q(\out_reg[11] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[11] [0]));
  _HDFF_verplex \out_reg_reg[12][8] (.Q(\out_reg[12] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[12] [8]));
  _HDFF_verplex \out_reg_reg[12][7] (.Q(\out_reg[12] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[12] [7]));
  _HDFF_verplex \out_reg_reg[12][6] (.Q(\out_reg[12] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[12] [6]));
  _HDFF_verplex \out_reg_reg[12][5] (.Q(\out_reg[12] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[12] [5]));
  _HDFF_verplex \out_reg_reg[12][4] (.Q(\out_reg[12] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[12] [4]));
  _HDFF_verplex \out_reg_reg[12][3] (.Q(\out_reg[12] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[12] [3]));
  _HDFF_verplex \out_reg_reg[12][2] (.Q(\out_reg[12] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[12] [2]));
  _HDFF_verplex \out_reg_reg[12][1] (.Q(\out_reg[12] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[12] [1]));
  _HDFF_verplex \out_reg_reg[12][0] (.Q(\out_reg[12] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[12] [0]));
  _HDFF_verplex \out_reg_reg[13][8] (.Q(\out_reg[13] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[13] [8]));
  _HDFF_verplex \out_reg_reg[13][7] (.Q(\out_reg[13] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[13] [7]));
  _HDFF_verplex \out_reg_reg[13][6] (.Q(\out_reg[13] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[13] [6]));
  _HDFF_verplex \out_reg_reg[13][5] (.Q(\out_reg[13] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[13] [5]));
  _HDFF_verplex \out_reg_reg[13][4] (.Q(\out_reg[13] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[13] [4]));
  _HDFF_verplex \out_reg_reg[13][3] (.Q(\out_reg[13] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[13] [3]));
  _HDFF_verplex \out_reg_reg[13][2] (.Q(\out_reg[13] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[13] [2]));
  _HDFF_verplex \out_reg_reg[13][1] (.Q(\out_reg[13] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[13] [1]));
  _HDFF_verplex \out_reg_reg[13][0] (.Q(\out_reg[13] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[13] [0]));
  _HDFF_verplex \out_reg_reg[14][8] (.Q(\out_reg[14] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[14] [8]));
  _HDFF_verplex \out_reg_reg[14][7] (.Q(\out_reg[14] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[14] [7]));
  _HDFF_verplex \out_reg_reg[14][6] (.Q(\out_reg[14] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[14] [6]));
  _HDFF_verplex \out_reg_reg[14][5] (.Q(\out_reg[14] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[14] [5]));
  _HDFF_verplex \out_reg_reg[14][4] (.Q(\out_reg[14] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[14] [4]));
  _HDFF_verplex \out_reg_reg[14][3] (.Q(\out_reg[14] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[14] [3]));
  _HDFF_verplex \out_reg_reg[14][2] (.Q(\out_reg[14] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[14] [2]));
  _HDFF_verplex \out_reg_reg[14][1] (.Q(\out_reg[14] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[14] [1]));
  _HDFF_verplex \out_reg_reg[14][0] (.Q(\out_reg[14] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[14] [0]));
  _HDFF_verplex \out_reg_reg[15][8] (.Q(\out_reg[15] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[15] [8]));
  _HDFF_verplex \out_reg_reg[15][7] (.Q(\out_reg[15] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[15] [7]));
  _HDFF_verplex \out_reg_reg[15][6] (.Q(\out_reg[15] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[15] [6]));
  _HDFF_verplex \out_reg_reg[15][5] (.Q(\out_reg[15] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[15] [5]));
  _HDFF_verplex \out_reg_reg[15][4] (.Q(\out_reg[15] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[15] [4]));
  _HDFF_verplex \out_reg_reg[15][3] (.Q(\out_reg[15] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[15] [3]));
  _HDFF_verplex \out_reg_reg[15][2] (.Q(\out_reg[15] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[15] [2]));
  _HDFF_verplex \out_reg_reg[15][1] (.Q(\out_reg[15] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[15] [1]));
  _HDFF_verplex \out_reg_reg[15][0] (.Q(\out_reg[15] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[15] [0]));
  _HDFF_verplex \out_reg_reg[16][8] (.Q(\out_reg[16] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[16] [8]));
  _HDFF_verplex \out_reg_reg[16][7] (.Q(\out_reg[16] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[16] [7]));
  _HDFF_verplex \out_reg_reg[16][6] (.Q(\out_reg[16] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[16] [6]));
  _HDFF_verplex \out_reg_reg[16][5] (.Q(\out_reg[16] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[16] [5]));
  _HDFF_verplex \out_reg_reg[16][4] (.Q(\out_reg[16] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[16] [4]));
  _HDFF_verplex \out_reg_reg[16][3] (.Q(\out_reg[16] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[16] [3]));
  _HDFF_verplex \out_reg_reg[16][2] (.Q(\out_reg[16] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[16] [2]));
  _HDFF_verplex \out_reg_reg[16][1] (.Q(\out_reg[16] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[16] [1]));
  _HDFF_verplex \out_reg_reg[16][0] (.Q(\out_reg[16] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[16] [0]));
  _HDFF_verplex \out_reg_reg[17][8] (.Q(\out_reg[17] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[17] [8]));
  _HDFF_verplex \out_reg_reg[17][7] (.Q(\out_reg[17] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[17] [7]));
  _HDFF_verplex \out_reg_reg[17][6] (.Q(\out_reg[17] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[17] [6]));
  _HDFF_verplex \out_reg_reg[17][5] (.Q(\out_reg[17] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[17] [5]));
  _HDFF_verplex \out_reg_reg[17][4] (.Q(\out_reg[17] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[17] [4]));
  _HDFF_verplex \out_reg_reg[17][3] (.Q(\out_reg[17] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[17] [3]));
  _HDFF_verplex \out_reg_reg[17][2] (.Q(\out_reg[17] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[17] [2]));
  _HDFF_verplex \out_reg_reg[17][1] (.Q(\out_reg[17] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[17] [1]));
  _HDFF_verplex \out_reg_reg[17][0] (.Q(\out_reg[17] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[17] [0]));
  _HDFF_verplex \out_reg_reg[18][8] (.Q(\out_reg[18] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[18] [8]));
  _HDFF_verplex \out_reg_reg[18][7] (.Q(\out_reg[18] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[18] [7]));
  _HDFF_verplex \out_reg_reg[18][6] (.Q(\out_reg[18] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[18] [6]));
  _HDFF_verplex \out_reg_reg[18][5] (.Q(\out_reg[18] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[18] [5]));
  _HDFF_verplex \out_reg_reg[18][4] (.Q(\out_reg[18] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[18] [4]));
  _HDFF_verplex \out_reg_reg[18][3] (.Q(\out_reg[18] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[18] [3]));
  _HDFF_verplex \out_reg_reg[18][2] (.Q(\out_reg[18] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[18] [2]));
  _HDFF_verplex \out_reg_reg[18][1] (.Q(\out_reg[18] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[18] [1]));
  _HDFF_verplex \out_reg_reg[18][0] (.Q(\out_reg[18] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[18] [0]));
  _HDFF_verplex \out_reg_reg[19][8] (.Q(\out_reg[19] [8]), .QN( ), .S(N$9), .R(
    n5413), .CK(clk), .D(\out_sig[19] [8]));
  _HDFF_verplex \out_reg_reg[19][7] (.Q(\out_reg[19] [7]), .QN( ), .S(N$8), .R(
    n5413), .CK(clk), .D(\out_sig[19] [7]));
  _HDFF_verplex \out_reg_reg[19][6] (.Q(\out_reg[19] [6]), .QN( ), .S(N$7), .R(
    n5413), .CK(clk), .D(\out_sig[19] [6]));
  _HDFF_verplex \out_reg_reg[19][5] (.Q(\out_reg[19] [5]), .QN( ), .S(N$6), .R(
    n5413), .CK(clk), .D(\out_sig[19] [5]));
  _HDFF_verplex \out_reg_reg[19][4] (.Q(\out_reg[19] [4]), .QN( ), .S(N$5), .R(
    n5413), .CK(clk), .D(\out_sig[19] [4]));
  _HDFF_verplex \out_reg_reg[19][3] (.Q(\out_reg[19] [3]), .QN( ), .S(N$4), .R(
    n5413), .CK(clk), .D(\out_sig[19] [3]));
  _HDFF_verplex \out_reg_reg[19][2] (.Q(\out_reg[19] [2]), .QN( ), .S(N$3), .R(
    n5413), .CK(clk), .D(\out_sig[19] [2]));
  _HDFF_verplex \out_reg_reg[19][1] (.Q(\out_reg[19] [1]), .QN( ), .S(N$2), .R(
    n5413), .CK(clk), .D(\out_sig[19] [1]));
  _HDFF_verplex \out_reg_reg[19][0] (.Q(\out_reg[19] [0]), .QN( ), .S(N$1), .R(
    n5413), .CK(clk), .D(\out_sig[19] [0]));
  VDW_ADD_10_1_0 add_5494_52_I1(.SUM({ \final_sums[0] [9:0] }), .A({ \level_8_sums[0] [9:0] }), .B({ \biases_l1_ext[0] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I2(.SUM({ \final_sums[1] [9:0] }), .A({ \level_8_sums[1] [9:0] }), .B({ \biases_l1_ext[1] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I3(.SUM({ \final_sums[2] [9:0] }), .A({ \level_8_sums[2] [9:0] }), .B({ \biases_l1_ext[2] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I4(.SUM({ \final_sums[3] [9:0] }), .A({ \level_8_sums[3] [9:0] }), .B({ \biases_l1_ext[3] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I5(.SUM({ \final_sums[4] [9:0] }), .A({ \level_8_sums[4] [9:0] }), .B({ \biases_l1_ext[4] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I6(.SUM({ \final_sums[5] [9:0] }), .A({ \level_8_sums[5] [9:0] }), .B({ \biases_l1_ext[5] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I7(.SUM({ \final_sums[6] [9:0] }), .A({ \level_8_sums[6] [9:0] }), .B({ \biases_l1_ext[6] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I8(.SUM({ \final_sums[7] [9:0] }), .A({ \level_8_sums[7] [9:0] }), .B({ \biases_l1_ext[7] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I9(.SUM({ \final_sums[8] [9:0] }), .A({ \level_8_sums[8] [9:0] }), .B({ \biases_l1_ext[8] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I10(.SUM({ \final_sums[9] [9:0] }), .A({ \level_8_sums[9] [9:0] }), .B({ \biases_l1_ext[9] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I11(.SUM({ \final_sums[10] [9:0] }), .A({ \level_8_sums[10] [9:0] }), .B({ \biases_l1_ext[10] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I12(.SUM({ \final_sums[11] [9:0] }), .A({ \level_8_sums[11] [9:0] }), .B({ \biases_l1_ext[11] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I13(.SUM({ \final_sums[12] [9:0] }), .A({ \level_8_sums[12] [9:0] }), .B({ \biases_l1_ext[12] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I14(.SUM({ \final_sums[13] [9:0] }), .A({ \level_8_sums[13] [9:0] }), .B({ \biases_l1_ext[13] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I15(.SUM({ \final_sums[14] [9:0] }), .A({ \level_8_sums[14] [9:0] }), .B({ \biases_l1_ext[14] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I16(.SUM({ \final_sums[15] [9:0] }), .A({ \level_8_sums[15] [9:0] }), .B({ \biases_l1_ext[15] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I17(.SUM({ \final_sums[16] [9:0] }), .A({ \level_8_sums[16] [9:0] }), .B({ \biases_l1_ext[16] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I18(.SUM({ \final_sums[17] [9:0] }), .A({ \level_8_sums[17] [9:0] }), .B({ \biases_l1_ext[17] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I19(.SUM({ \final_sums[18] [9:0] }), .A({ \level_8_sums[18] [9:0] }), .B({ \biases_l1_ext[18] [9:0] }));
  VDW_ADD_10_1_0 add_5494_52_I20(.SUM({ \final_sums[19] [9:0] }), .A({ \level_8_sums[19] [9:0] }), .B({ \biases_l1_ext[19] [9:0] }));
  assign \biases_l1_ext[0] [9] = \biases_l1[0] [6];
  assign \biases_l1_ext[0] [8] = \biases_l1[0] [6];
  assign \biases_l1_ext[0] [7] = \biases_l1[0] [6];
  assign \biases_l1_ext[0] [6] = \biases_l1[0] [6];
  assign \biases_l1_ext[0] [5] = \biases_l1[0] [5];
  assign \biases_l1_ext[0] [4] = \biases_l1[0] [4];
  assign \biases_l1_ext[0] [3] = \biases_l1[0] [3];
  assign \biases_l1_ext[0] [2] = \biases_l1[0] [2];
  assign \biases_l1_ext[0] [1] = \biases_l1[0] [1];
  assign \biases_l1_ext[0] [0] = \biases_l1[0] [0];
  assign \biases_l1_ext[1] [9] = \biases_l1[1] [6];
  assign \biases_l1_ext[1] [8] = \biases_l1[1] [6];
  assign \biases_l1_ext[1] [7] = \biases_l1[1] [6];
  assign \biases_l1_ext[1] [6] = \biases_l1[1] [6];
  assign \biases_l1_ext[1] [5] = \biases_l1[1] [5];
  assign \biases_l1_ext[1] [4] = \biases_l1[1] [4];
  assign \biases_l1_ext[1] [3] = \biases_l1[1] [3];
  assign \biases_l1_ext[1] [2] = \biases_l1[1] [2];
  assign \biases_l1_ext[1] [1] = \biases_l1[1] [1];
  assign \biases_l1_ext[1] [0] = \biases_l1[1] [0];
  assign \biases_l1_ext[2] [9] = \biases_l1[2] [6];
  assign \biases_l1_ext[2] [8] = \biases_l1[2] [6];
  assign \biases_l1_ext[2] [7] = \biases_l1[2] [6];
  assign \biases_l1_ext[2] [6] = \biases_l1[2] [6];
  assign \biases_l1_ext[2] [5] = \biases_l1[2] [5];
  assign \biases_l1_ext[2] [4] = \biases_l1[2] [4];
  assign \biases_l1_ext[2] [3] = \biases_l1[2] [3];
  assign \biases_l1_ext[2] [2] = \biases_l1[2] [2];
  assign \biases_l1_ext[2] [1] = \biases_l1[2] [1];
  assign \biases_l1_ext[2] [0] = \biases_l1[2] [0];
  assign \biases_l1_ext[3] [9] = \biases_l1[3] [6];
  assign \biases_l1_ext[3] [8] = \biases_l1[3] [6];
  assign \biases_l1_ext[3] [7] = \biases_l1[3] [6];
  assign \biases_l1_ext[3] [6] = \biases_l1[3] [6];
  assign \biases_l1_ext[3] [5] = \biases_l1[3] [5];
  assign \biases_l1_ext[3] [4] = \biases_l1[3] [4];
  assign \biases_l1_ext[3] [3] = \biases_l1[3] [3];
  assign \biases_l1_ext[3] [2] = \biases_l1[3] [2];
  assign \biases_l1_ext[3] [1] = \biases_l1[3] [1];
  assign \biases_l1_ext[3] [0] = \biases_l1[3] [0];
  assign \biases_l1_ext[4] [9] = \biases_l1[4] [6];
  assign \biases_l1_ext[4] [8] = \biases_l1[4] [6];
  assign \biases_l1_ext[4] [7] = \biases_l1[4] [6];
  assign \biases_l1_ext[4] [6] = \biases_l1[4] [6];
  assign \biases_l1_ext[4] [5] = \biases_l1[4] [5];
  assign \biases_l1_ext[4] [4] = \biases_l1[4] [4];
  assign \biases_l1_ext[4] [3] = \biases_l1[4] [3];
  assign \biases_l1_ext[4] [2] = \biases_l1[4] [2];
  assign \biases_l1_ext[4] [1] = \biases_l1[4] [1];
  assign \biases_l1_ext[4] [0] = \biases_l1[4] [0];
  assign \biases_l1_ext[5] [9] = \biases_l1[5] [6];
  assign \biases_l1_ext[5] [8] = \biases_l1[5] [6];
  assign \biases_l1_ext[5] [7] = \biases_l1[5] [6];
  assign \biases_l1_ext[5] [6] = \biases_l1[5] [6];
  assign \biases_l1_ext[5] [5] = \biases_l1[5] [5];
  assign \biases_l1_ext[5] [4] = \biases_l1[5] [4];
  assign \biases_l1_ext[5] [3] = \biases_l1[5] [3];
  assign \biases_l1_ext[5] [2] = \biases_l1[5] [2];
  assign \biases_l1_ext[5] [1] = \biases_l1[5] [1];
  assign \biases_l1_ext[5] [0] = \biases_l1[5] [0];
  assign \biases_l1_ext[6] [9] = \biases_l1[6] [6];
  assign \biases_l1_ext[6] [8] = \biases_l1[6] [6];
  assign \biases_l1_ext[6] [7] = \biases_l1[6] [6];
  assign \biases_l1_ext[6] [6] = \biases_l1[6] [6];
  assign \biases_l1_ext[6] [5] = \biases_l1[6] [5];
  assign \biases_l1_ext[6] [4] = \biases_l1[6] [4];
  assign \biases_l1_ext[6] [3] = \biases_l1[6] [3];
  assign \biases_l1_ext[6] [2] = \biases_l1[6] [2];
  assign \biases_l1_ext[6] [1] = \biases_l1[6] [1];
  assign \biases_l1_ext[6] [0] = \biases_l1[6] [0];
  assign \biases_l1_ext[7] [9] = \biases_l1[7] [6];
  assign \biases_l1_ext[7] [8] = \biases_l1[7] [6];
  assign \biases_l1_ext[7] [7] = \biases_l1[7] [6];
  assign \biases_l1_ext[7] [6] = \biases_l1[7] [6];
  assign \biases_l1_ext[7] [5] = \biases_l1[7] [5];
  assign \biases_l1_ext[7] [4] = \biases_l1[7] [4];
  assign \biases_l1_ext[7] [3] = \biases_l1[7] [3];
  assign \biases_l1_ext[7] [2] = \biases_l1[7] [2];
  assign \biases_l1_ext[7] [1] = \biases_l1[7] [1];
  assign \biases_l1_ext[7] [0] = \biases_l1[7] [0];
  assign \biases_l1_ext[8] [9] = \biases_l1[8] [6];
  assign \biases_l1_ext[8] [8] = \biases_l1[8] [6];
  assign \biases_l1_ext[8] [7] = \biases_l1[8] [6];
  assign \biases_l1_ext[8] [6] = \biases_l1[8] [6];
  assign \biases_l1_ext[8] [5] = \biases_l1[8] [5];
  assign \biases_l1_ext[8] [4] = \biases_l1[8] [4];
  assign \biases_l1_ext[8] [3] = \biases_l1[8] [3];
  assign \biases_l1_ext[8] [2] = \biases_l1[8] [2];
  assign \biases_l1_ext[8] [1] = \biases_l1[8] [1];
  assign \biases_l1_ext[8] [0] = \biases_l1[8] [0];
  assign \biases_l1_ext[9] [9] = \biases_l1[9] [6];
  assign \biases_l1_ext[9] [8] = \biases_l1[9] [6];
  assign \biases_l1_ext[9] [7] = \biases_l1[9] [6];
  assign \biases_l1_ext[9] [6] = \biases_l1[9] [6];
  assign \biases_l1_ext[9] [5] = \biases_l1[9] [5];
  assign \biases_l1_ext[9] [4] = \biases_l1[9] [4];
  assign \biases_l1_ext[9] [3] = \biases_l1[9] [3];
  assign \biases_l1_ext[9] [2] = \biases_l1[9] [2];
  assign \biases_l1_ext[9] [1] = \biases_l1[9] [1];
  assign \biases_l1_ext[9] [0] = \biases_l1[9] [0];
  assign \biases_l1_ext[10] [9] = \biases_l1[10] [6];
  assign \biases_l1_ext[10] [8] = \biases_l1[10] [6];
  assign \biases_l1_ext[10] [7] = \biases_l1[10] [6];
  assign \biases_l1_ext[10] [6] = \biases_l1[10] [6];
  assign \biases_l1_ext[10] [5] = \biases_l1[10] [5];
  assign \biases_l1_ext[10] [4] = \biases_l1[10] [4];
  assign \biases_l1_ext[10] [3] = \biases_l1[10] [3];
  assign \biases_l1_ext[10] [2] = \biases_l1[10] [2];
  assign \biases_l1_ext[10] [1] = \biases_l1[10] [1];
  assign \biases_l1_ext[10] [0] = \biases_l1[10] [0];
  assign \biases_l1_ext[11] [9] = \biases_l1[11] [6];
  assign \biases_l1_ext[11] [8] = \biases_l1[11] [6];
  assign \biases_l1_ext[11] [7] = \biases_l1[11] [6];
  assign \biases_l1_ext[11] [6] = \biases_l1[11] [6];
  assign \biases_l1_ext[11] [5] = \biases_l1[11] [5];
  assign \biases_l1_ext[11] [4] = \biases_l1[11] [4];
  assign \biases_l1_ext[11] [3] = \biases_l1[11] [3];
  assign \biases_l1_ext[11] [2] = \biases_l1[11] [2];
  assign \biases_l1_ext[11] [1] = \biases_l1[11] [1];
  assign \biases_l1_ext[11] [0] = \biases_l1[11] [0];
  assign \biases_l1_ext[12] [9] = \biases_l1[12] [6];
  assign \biases_l1_ext[12] [8] = \biases_l1[12] [6];
  assign \biases_l1_ext[12] [7] = \biases_l1[12] [6];
  assign \biases_l1_ext[12] [6] = \biases_l1[12] [6];
  assign \biases_l1_ext[12] [5] = \biases_l1[12] [5];
  assign \biases_l1_ext[12] [4] = \biases_l1[12] [4];
  assign \biases_l1_ext[12] [3] = \biases_l1[12] [3];
  assign \biases_l1_ext[12] [2] = \biases_l1[12] [2];
  assign \biases_l1_ext[12] [1] = \biases_l1[12] [1];
  assign \biases_l1_ext[12] [0] = \biases_l1[12] [0];
  assign \biases_l1_ext[13] [9] = \biases_l1[13] [6];
  assign \biases_l1_ext[13] [8] = \biases_l1[13] [6];
  assign \biases_l1_ext[13] [7] = \biases_l1[13] [6];
  assign \biases_l1_ext[13] [6] = \biases_l1[13] [6];
  assign \biases_l1_ext[13] [5] = \biases_l1[13] [5];
  assign \biases_l1_ext[13] [4] = \biases_l1[13] [4];
  assign \biases_l1_ext[13] [3] = \biases_l1[13] [3];
  assign \biases_l1_ext[13] [2] = \biases_l1[13] [2];
  assign \biases_l1_ext[13] [1] = \biases_l1[13] [1];
  assign \biases_l1_ext[13] [0] = \biases_l1[13] [0];
  assign \biases_l1_ext[14] [9] = \biases_l1[14] [6];
  assign \biases_l1_ext[14] [8] = \biases_l1[14] [6];
  assign \biases_l1_ext[14] [7] = \biases_l1[14] [6];
  assign \biases_l1_ext[14] [6] = \biases_l1[14] [6];
  assign \biases_l1_ext[14] [5] = \biases_l1[14] [5];
  assign \biases_l1_ext[14] [4] = \biases_l1[14] [4];
  assign \biases_l1_ext[14] [3] = \biases_l1[14] [3];
  assign \biases_l1_ext[14] [2] = \biases_l1[14] [2];
  assign \biases_l1_ext[14] [1] = \biases_l1[14] [1];
  assign \biases_l1_ext[14] [0] = \biases_l1[14] [0];
  assign \biases_l1_ext[15] [9] = \biases_l1[15] [6];
  assign \biases_l1_ext[15] [8] = \biases_l1[15] [6];
  assign \biases_l1_ext[15] [7] = \biases_l1[15] [6];
  assign \biases_l1_ext[15] [6] = \biases_l1[15] [6];
  assign \biases_l1_ext[15] [5] = \biases_l1[15] [5];
  assign \biases_l1_ext[15] [4] = \biases_l1[15] [4];
  assign \biases_l1_ext[15] [3] = \biases_l1[15] [3];
  assign \biases_l1_ext[15] [2] = \biases_l1[15] [2];
  assign \biases_l1_ext[15] [1] = \biases_l1[15] [1];
  assign \biases_l1_ext[15] [0] = \biases_l1[15] [0];
  assign \biases_l1_ext[16] [9] = \biases_l1[16] [6];
  assign \biases_l1_ext[16] [8] = \biases_l1[16] [6];
  assign \biases_l1_ext[16] [7] = \biases_l1[16] [6];
  assign \biases_l1_ext[16] [6] = \biases_l1[16] [6];
  assign \biases_l1_ext[16] [5] = \biases_l1[16] [5];
  assign \biases_l1_ext[16] [4] = \biases_l1[16] [4];
  assign \biases_l1_ext[16] [3] = \biases_l1[16] [3];
  assign \biases_l1_ext[16] [2] = \biases_l1[16] [2];
  assign \biases_l1_ext[16] [1] = \biases_l1[16] [1];
  assign \biases_l1_ext[16] [0] = \biases_l1[16] [0];
  assign \biases_l1_ext[17] [9] = \biases_l1[17] [6];
  assign \biases_l1_ext[17] [8] = \biases_l1[17] [6];
  assign \biases_l1_ext[17] [7] = \biases_l1[17] [6];
  assign \biases_l1_ext[17] [6] = \biases_l1[17] [6];
  assign \biases_l1_ext[17] [5] = \biases_l1[17] [5];
  assign \biases_l1_ext[17] [4] = \biases_l1[17] [4];
  assign \biases_l1_ext[17] [3] = \biases_l1[17] [3];
  assign \biases_l1_ext[17] [2] = \biases_l1[17] [2];
  assign \biases_l1_ext[17] [1] = \biases_l1[17] [1];
  assign \biases_l1_ext[17] [0] = \biases_l1[17] [0];
  assign \biases_l1_ext[18] [9] = \biases_l1[18] [6];
  assign \biases_l1_ext[18] [8] = \biases_l1[18] [6];
  assign \biases_l1_ext[18] [7] = \biases_l1[18] [6];
  assign \biases_l1_ext[18] [6] = \biases_l1[18] [6];
  assign \biases_l1_ext[18] [5] = \biases_l1[18] [5];
  assign \biases_l1_ext[18] [4] = \biases_l1[18] [4];
  assign \biases_l1_ext[18] [3] = \biases_l1[18] [3];
  assign \biases_l1_ext[18] [2] = \biases_l1[18] [2];
  assign \biases_l1_ext[18] [1] = \biases_l1[18] [1];
  assign \biases_l1_ext[18] [0] = \biases_l1[18] [0];
  assign \biases_l1_ext[19] [9] = \biases_l1[19] [6];
  assign \biases_l1_ext[19] [8] = \biases_l1[19] [6];
  assign \biases_l1_ext[19] [7] = \biases_l1[19] [6];
  assign \biases_l1_ext[19] [6] = \biases_l1[19] [6];
  assign \biases_l1_ext[19] [5] = \biases_l1[19] [5];
  assign \biases_l1_ext[19] [4] = \biases_l1[19] [4];
  assign \biases_l1_ext[19] [3] = \biases_l1[19] [3];
  assign \biases_l1_ext[19] [2] = \biases_l1[19] [2];
  assign \biases_l1_ext[19] [1] = \biases_l1[19] [1];
  assign \biases_l1_ext[19] [0] = \biases_l1[19] [0];
  _HDFF_verplex \B_reg[0] (.Q(B[0]), .QN( ), .S(N$265), .R(n5413), .CK(clk), .D(
    n5418[255]));
  _HDFF_verplex \B_reg[1] (.Q(B[1]), .QN( ), .S(N$264), .R(n5413), .CK(clk), .D(
    n5418[254]));
  _HDFF_verplex \B_reg[2] (.Q(B[2]), .QN( ), .S(N$263), .R(n5413), .CK(clk), .D(
    n5418[253]));
  _HDFF_verplex \B_reg[3] (.Q(B[3]), .QN( ), .S(N$262), .R(n5413), .CK(clk), .D(
    n5418[252]));
  _HDFF_verplex \B_reg[4] (.Q(B[4]), .QN( ), .S(N$261), .R(n5413), .CK(clk), .D(
    n5418[251]));
  _HDFF_verplex \B_reg[5] (.Q(B[5]), .QN( ), .S(N$260), .R(n5413), .CK(clk), .D(
    n5418[250]));
  _HDFF_verplex \B_reg[6] (.Q(B[6]), .QN( ), .S(N$259), .R(n5413), .CK(clk), .D(
    n5418[249]));
  _HDFF_verplex \B_reg[7] (.Q(B[7]), .QN( ), .S(N$258), .R(n5413), .CK(clk), .D(
    n5418[248]));
  _HDFF_verplex \B_reg[8] (.Q(B[8]), .QN( ), .S(N$257), .R(n5413), .CK(clk), .D(
    n5418[247]));
  _HDFF_verplex \B_reg[9] (.Q(B[9]), .QN( ), .S(N$256), .R(n5413), .CK(clk), .D(
    n5418[246]));
  _HDFF_verplex \B_reg[10] (.Q(B[10]), .QN( ), .S(N$255), .R(n5413), .CK(clk)
    , .D(n5418[245]));
  _HDFF_verplex \B_reg[11] (.Q(B[11]), .QN( ), .S(N$254), .R(n5413), .CK(clk)
    , .D(n5418[244]));
  _HDFF_verplex \B_reg[12] (.Q(B[12]), .QN( ), .S(N$253), .R(n5413), .CK(clk)
    , .D(n5418[243]));
  _HDFF_verplex \B_reg[13] (.Q(B[13]), .QN( ), .S(N$252), .R(n5413), .CK(clk)
    , .D(n5418[242]));
  _HDFF_verplex \B_reg[14] (.Q(B[14]), .QN( ), .S(N$251), .R(n5413), .CK(clk)
    , .D(n5418[241]));
  _HDFF_verplex \B_reg[15] (.Q(B[15]), .QN( ), .S(N$250), .R(n5413), .CK(clk)
    , .D(n5418[240]));
  _HDFF_verplex \B_reg[16] (.Q(B[16]), .QN( ), .S(N$249), .R(n5413), .CK(clk)
    , .D(n5418[239]));
  _HDFF_verplex \B_reg[17] (.Q(B[17]), .QN( ), .S(N$248), .R(n5413), .CK(clk)
    , .D(n5418[238]));
  _HDFF_verplex \B_reg[18] (.Q(B[18]), .QN( ), .S(N$247), .R(n5413), .CK(clk)
    , .D(n5418[237]));
  _HDFF_verplex \B_reg[19] (.Q(B[19]), .QN( ), .S(N$246), .R(n5413), .CK(clk)
    , .D(n5418[236]));
  _HDFF_verplex \B_reg[20] (.Q(B[20]), .QN( ), .S(N$245), .R(n5413), .CK(clk)
    , .D(n5418[235]));
  _HDFF_verplex \B_reg[21] (.Q(B[21]), .QN( ), .S(N$244), .R(n5413), .CK(clk)
    , .D(n5418[234]));
  _HDFF_verplex \B_reg[22] (.Q(B[22]), .QN( ), .S(N$243), .R(n5413), .CK(clk)
    , .D(n5418[233]));
  _HDFF_verplex \B_reg[23] (.Q(B[23]), .QN( ), .S(N$242), .R(n5413), .CK(clk)
    , .D(n5418[232]));
  _HDFF_verplex \B_reg[24] (.Q(B[24]), .QN( ), .S(N$241), .R(n5413), .CK(clk)
    , .D(n5418[231]));
  _HDFF_verplex \B_reg[25] (.Q(B[25]), .QN( ), .S(N$240), .R(n5413), .CK(clk)
    , .D(n5418[230]));
  _HDFF_verplex \B_reg[26] (.Q(B[26]), .QN( ), .S(N$239), .R(n5413), .CK(clk)
    , .D(n5418[229]));
  _HDFF_verplex \B_reg[27] (.Q(B[27]), .QN( ), .S(N$238), .R(n5413), .CK(clk)
    , .D(n5418[228]));
  _HDFF_verplex \B_reg[28] (.Q(B[28]), .QN( ), .S(N$237), .R(n5413), .CK(clk)
    , .D(n5418[227]));
  _HDFF_verplex \B_reg[29] (.Q(B[29]), .QN( ), .S(N$236), .R(n5413), .CK(clk)
    , .D(n5418[226]));
  _HDFF_verplex \B_reg[30] (.Q(B[30]), .QN( ), .S(N$235), .R(n5413), .CK(clk)
    , .D(n5418[225]));
  _HDFF_verplex \B_reg[31] (.Q(B[31]), .QN( ), .S(N$234), .R(n5413), .CK(clk)
    , .D(n5418[224]));
  _HDFF_verplex \B_reg[32] (.Q(B[32]), .QN( ), .S(N$233), .R(n5413), .CK(clk)
    , .D(n5418[223]));
  _HDFF_verplex \B_reg[33] (.Q(B[33]), .QN( ), .S(N$232), .R(n5413), .CK(clk)
    , .D(n5418[222]));
  _HDFF_verplex \B_reg[34] (.Q(B[34]), .QN( ), .S(N$231), .R(n5413), .CK(clk)
    , .D(n5418[221]));
  _HDFF_verplex \B_reg[35] (.Q(B[35]), .QN( ), .S(N$230), .R(n5413), .CK(clk)
    , .D(n5418[220]));
  _HDFF_verplex \B_reg[36] (.Q(B[36]), .QN( ), .S(N$229), .R(n5413), .CK(clk)
    , .D(n5418[219]));
  _HDFF_verplex \B_reg[37] (.Q(B[37]), .QN( ), .S(N$228), .R(n5413), .CK(clk)
    , .D(n5418[218]));
  _HDFF_verplex \B_reg[38] (.Q(B[38]), .QN( ), .S(N$227), .R(n5413), .CK(clk)
    , .D(n5418[217]));
  _HDFF_verplex \B_reg[39] (.Q(B[39]), .QN( ), .S(N$226), .R(n5413), .CK(clk)
    , .D(n5418[216]));
  _HDFF_verplex \B_reg[40] (.Q(B[40]), .QN( ), .S(N$225), .R(n5413), .CK(clk)
    , .D(n5418[215]));
  _HDFF_verplex \B_reg[41] (.Q(B[41]), .QN( ), .S(N$224), .R(n5413), .CK(clk)
    , .D(n5418[214]));
  _HDFF_verplex \B_reg[42] (.Q(B[42]), .QN( ), .S(N$223), .R(n5413), .CK(clk)
    , .D(n5418[213]));
  _HDFF_verplex \B_reg[43] (.Q(B[43]), .QN( ), .S(N$222), .R(n5413), .CK(clk)
    , .D(n5418[212]));
  _HDFF_verplex \B_reg[44] (.Q(B[44]), .QN( ), .S(N$221), .R(n5413), .CK(clk)
    , .D(n5418[211]));
  _HDFF_verplex \B_reg[45] (.Q(B[45]), .QN( ), .S(N$220), .R(n5413), .CK(clk)
    , .D(n5418[210]));
  _HDFF_verplex \B_reg[46] (.Q(B[46]), .QN( ), .S(N$219), .R(n5413), .CK(clk)
    , .D(n5418[209]));
  _HDFF_verplex \B_reg[47] (.Q(B[47]), .QN( ), .S(N$218), .R(n5413), .CK(clk)
    , .D(n5418[208]));
  _HDFF_verplex \B_reg[48] (.Q(B[48]), .QN( ), .S(N$217), .R(n5413), .CK(clk)
    , .D(n5418[207]));
  _HDFF_verplex \B_reg[49] (.Q(B[49]), .QN( ), .S(N$216), .R(n5413), .CK(clk)
    , .D(n5418[206]));
  _HDFF_verplex \B_reg[50] (.Q(B[50]), .QN( ), .S(N$215), .R(n5413), .CK(clk)
    , .D(n5418[205]));
  _HDFF_verplex \B_reg[51] (.Q(B[51]), .QN( ), .S(N$214), .R(n5413), .CK(clk)
    , .D(n5418[204]));
  _HDFF_verplex \B_reg[52] (.Q(B[52]), .QN( ), .S(N$213), .R(n5413), .CK(clk)
    , .D(n5418[203]));
  _HDFF_verplex \B_reg[53] (.Q(B[53]), .QN( ), .S(N$212), .R(n5413), .CK(clk)
    , .D(n5418[202]));
  _HDFF_verplex \B_reg[54] (.Q(B[54]), .QN( ), .S(N$211), .R(n5413), .CK(clk)
    , .D(n5418[201]));
  _HDFF_verplex \B_reg[55] (.Q(B[55]), .QN( ), .S(N$210), .R(n5413), .CK(clk)
    , .D(n5418[200]));
  _HDFF_verplex \B_reg[56] (.Q(B[56]), .QN( ), .S(N$209), .R(n5413), .CK(clk)
    , .D(n5418[199]));
  _HDFF_verplex \B_reg[57] (.Q(B[57]), .QN( ), .S(N$208), .R(n5413), .CK(clk)
    , .D(n5418[198]));
  _HDFF_verplex \B_reg[58] (.Q(B[58]), .QN( ), .S(N$207), .R(n5413), .CK(clk)
    , .D(n5418[197]));
  _HDFF_verplex \B_reg[59] (.Q(B[59]), .QN( ), .S(N$206), .R(n5413), .CK(clk)
    , .D(n5418[196]));
  _HDFF_verplex \B_reg[60] (.Q(B[60]), .QN( ), .S(N$205), .R(n5413), .CK(clk)
    , .D(n5418[195]));
  _HDFF_verplex \B_reg[61] (.Q(B[61]), .QN( ), .S(N$204), .R(n5413), .CK(clk)
    , .D(n5418[194]));
  _HDFF_verplex \B_reg[62] (.Q(B[62]), .QN( ), .S(N$203), .R(n5413), .CK(clk)
    , .D(n5418[193]));
  _HDFF_verplex \B_reg[63] (.Q(B[63]), .QN( ), .S(N$202), .R(n5413), .CK(clk)
    , .D(n5418[192]));
  _HDFF_verplex \B_reg[64] (.Q(B[64]), .QN( ), .S(N$201), .R(n5413), .CK(clk)
    , .D(n5418[191]));
  _HDFF_verplex \B_reg[65] (.Q(B[65]), .QN( ), .S(N$200), .R(n5413), .CK(clk)
    , .D(n5418[190]));
  _HDFF_verplex \B_reg[66] (.Q(B[66]), .QN( ), .S(N$199), .R(n5413), .CK(clk)
    , .D(n5418[189]));
  _HDFF_verplex \B_reg[67] (.Q(B[67]), .QN( ), .S(N$198), .R(n5413), .CK(clk)
    , .D(n5418[188]));
  _HDFF_verplex \B_reg[68] (.Q(B[68]), .QN( ), .S(N$197), .R(n5413), .CK(clk)
    , .D(n5418[187]));
  _HDFF_verplex \B_reg[69] (.Q(B[69]), .QN( ), .S(N$196), .R(n5413), .CK(clk)
    , .D(n5418[186]));
  _HDFF_verplex \B_reg[70] (.Q(B[70]), .QN( ), .S(N$195), .R(n5413), .CK(clk)
    , .D(n5418[185]));
  _HDFF_verplex \B_reg[71] (.Q(B[71]), .QN( ), .S(N$194), .R(n5413), .CK(clk)
    , .D(n5418[184]));
  _HDFF_verplex \B_reg[72] (.Q(B[72]), .QN( ), .S(N$193), .R(n5413), .CK(clk)
    , .D(n5418[183]));
  _HDFF_verplex \B_reg[73] (.Q(B[73]), .QN( ), .S(N$192), .R(n5413), .CK(clk)
    , .D(n5418[182]));
  _HDFF_verplex \B_reg[74] (.Q(B[74]), .QN( ), .S(N$191), .R(n5413), .CK(clk)
    , .D(n5418[181]));
  _HDFF_verplex \B_reg[75] (.Q(B[75]), .QN( ), .S(N$190), .R(n5413), .CK(clk)
    , .D(n5418[180]));
  _HDFF_verplex \B_reg[76] (.Q(B[76]), .QN( ), .S(N$189), .R(n5413), .CK(clk)
    , .D(n5418[179]));
  _HDFF_verplex \B_reg[77] (.Q(B[77]), .QN( ), .S(N$188), .R(n5413), .CK(clk)
    , .D(n5418[178]));
  _HDFF_verplex \B_reg[78] (.Q(B[78]), .QN( ), .S(N$187), .R(n5413), .CK(clk)
    , .D(n5418[177]));
  _HDFF_verplex \B_reg[79] (.Q(B[79]), .QN( ), .S(N$186), .R(n5413), .CK(clk)
    , .D(n5418[176]));
  _HDFF_verplex \B_reg[80] (.Q(B[80]), .QN( ), .S(N$185), .R(n5413), .CK(clk)
    , .D(n5418[175]));
  _HDFF_verplex \B_reg[81] (.Q(B[81]), .QN( ), .S(N$184), .R(n5413), .CK(clk)
    , .D(n5418[174]));
  _HDFF_verplex \B_reg[82] (.Q(B[82]), .QN( ), .S(N$183), .R(n5413), .CK(clk)
    , .D(n5418[173]));
  _HDFF_verplex \B_reg[83] (.Q(B[83]), .QN( ), .S(N$182), .R(n5413), .CK(clk)
    , .D(n5418[172]));
  _HDFF_verplex \B_reg[84] (.Q(B[84]), .QN( ), .S(N$181), .R(n5413), .CK(clk)
    , .D(n5418[171]));
  _HDFF_verplex \B_reg[85] (.Q(B[85]), .QN( ), .S(N$180), .R(n5413), .CK(clk)
    , .D(n5418[170]));
  _HDFF_verplex \B_reg[86] (.Q(B[86]), .QN( ), .S(N$179), .R(n5413), .CK(clk)
    , .D(n5418[169]));
  _HDFF_verplex \B_reg[87] (.Q(B[87]), .QN( ), .S(N$178), .R(n5413), .CK(clk)
    , .D(n5418[168]));
  _HDFF_verplex \B_reg[88] (.Q(B[88]), .QN( ), .S(N$177), .R(n5413), .CK(clk)
    , .D(n5418[167]));
  _HDFF_verplex \B_reg[89] (.Q(B[89]), .QN( ), .S(N$176), .R(n5413), .CK(clk)
    , .D(n5418[166]));
  _HDFF_verplex \B_reg[90] (.Q(B[90]), .QN( ), .S(N$175), .R(n5413), .CK(clk)
    , .D(n5418[165]));
  _HDFF_verplex \B_reg[91] (.Q(B[91]), .QN( ), .S(N$174), .R(n5413), .CK(clk)
    , .D(n5418[164]));
  _HDFF_verplex \B_reg[92] (.Q(B[92]), .QN( ), .S(N$173), .R(n5413), .CK(clk)
    , .D(n5418[163]));
  _HDFF_verplex \B_reg[93] (.Q(B[93]), .QN( ), .S(N$172), .R(n5413), .CK(clk)
    , .D(n5418[162]));
  _HDFF_verplex \B_reg[94] (.Q(B[94]), .QN( ), .S(N$171), .R(n5413), .CK(clk)
    , .D(n5418[161]));
  _HDFF_verplex \B_reg[95] (.Q(B[95]), .QN( ), .S(N$170), .R(n5413), .CK(clk)
    , .D(n5418[160]));
  _HDFF_verplex \B_reg[96] (.Q(B[96]), .QN( ), .S(N$169), .R(n5413), .CK(clk)
    , .D(n5418[159]));
  _HDFF_verplex \B_reg[97] (.Q(B[97]), .QN( ), .S(N$168), .R(n5413), .CK(clk)
    , .D(n5418[158]));
  _HDFF_verplex \B_reg[98] (.Q(B[98]), .QN( ), .S(N$167), .R(n5413), .CK(clk)
    , .D(n5418[157]));
  _HDFF_verplex \B_reg[99] (.Q(B[99]), .QN( ), .S(N$166), .R(n5413), .CK(clk)
    , .D(n5418[156]));
  _HDFF_verplex \B_reg[100] (.Q(B[100]), .QN( ), .S(N$165), .R(n5413), .CK(clk)
    , .D(n5418[155]));
  _HDFF_verplex \B_reg[101] (.Q(B[101]), .QN( ), .S(N$164), .R(n5413), .CK(clk)
    , .D(n5418[154]));
  _HDFF_verplex \B_reg[102] (.Q(B[102]), .QN( ), .S(N$163), .R(n5413), .CK(clk)
    , .D(n5418[153]));
  _HDFF_verplex \B_reg[103] (.Q(B[103]), .QN( ), .S(N$162), .R(n5413), .CK(clk)
    , .D(n5418[152]));
  _HDFF_verplex \B_reg[104] (.Q(B[104]), .QN( ), .S(N$161), .R(n5413), .CK(clk)
    , .D(n5418[151]));
  _HDFF_verplex \B_reg[105] (.Q(B[105]), .QN( ), .S(N$160), .R(n5413), .CK(clk)
    , .D(n5418[150]));
  _HDFF_verplex \B_reg[106] (.Q(B[106]), .QN( ), .S(N$159), .R(n5413), .CK(clk)
    , .D(n5418[149]));
  _HDFF_verplex \B_reg[107] (.Q(B[107]), .QN( ), .S(N$158), .R(n5413), .CK(clk)
    , .D(n5418[148]));
  _HDFF_verplex \B_reg[108] (.Q(B[108]), .QN( ), .S(N$157), .R(n5413), .CK(clk)
    , .D(n5418[147]));
  _HDFF_verplex \B_reg[109] (.Q(B[109]), .QN( ), .S(N$156), .R(n5413), .CK(clk)
    , .D(n5418[146]));
  _HDFF_verplex \B_reg[110] (.Q(B[110]), .QN( ), .S(N$155), .R(n5413), .CK(clk)
    , .D(n5418[145]));
  _HDFF_verplex \B_reg[111] (.Q(B[111]), .QN( ), .S(N$154), .R(n5413), .CK(clk)
    , .D(n5418[144]));
  _HDFF_verplex \B_reg[112] (.Q(B[112]), .QN( ), .S(N$153), .R(n5413), .CK(clk)
    , .D(n5418[143]));
  _HDFF_verplex \B_reg[113] (.Q(B[113]), .QN( ), .S(N$152), .R(n5413), .CK(clk)
    , .D(n5418[142]));
  _HDFF_verplex \B_reg[114] (.Q(B[114]), .QN( ), .S(N$151), .R(n5413), .CK(clk)
    , .D(n5418[141]));
  _HDFF_verplex \B_reg[115] (.Q(B[115]), .QN( ), .S(N$150), .R(n5413), .CK(clk)
    , .D(n5418[140]));
  _HDFF_verplex \B_reg[116] (.Q(B[116]), .QN( ), .S(N$149), .R(n5413), .CK(clk)
    , .D(n5418[139]));
  _HDFF_verplex \B_reg[117] (.Q(B[117]), .QN( ), .S(N$148), .R(n5413), .CK(clk)
    , .D(n5418[138]));
  _HDFF_verplex \B_reg[118] (.Q(B[118]), .QN( ), .S(N$147), .R(n5413), .CK(clk)
    , .D(n5418[137]));
  _HDFF_verplex \B_reg[119] (.Q(B[119]), .QN( ), .S(N$146), .R(n5413), .CK(clk)
    , .D(n5418[136]));
  _HDFF_verplex \B_reg[120] (.Q(B[120]), .QN( ), .S(N$145), .R(n5413), .CK(clk)
    , .D(n5418[135]));
  _HDFF_verplex \B_reg[121] (.Q(B[121]), .QN( ), .S(N$144), .R(n5413), .CK(clk)
    , .D(n5418[134]));
  _HDFF_verplex \B_reg[122] (.Q(B[122]), .QN( ), .S(N$143), .R(n5413), .CK(clk)
    , .D(n5418[133]));
  _HDFF_verplex \B_reg[123] (.Q(B[123]), .QN( ), .S(N$142), .R(n5413), .CK(clk)
    , .D(n5418[132]));
  _HDFF_verplex \B_reg[124] (.Q(B[124]), .QN( ), .S(N$141), .R(n5413), .CK(clk)
    , .D(n5418[131]));
  _HDFF_verplex \B_reg[125] (.Q(B[125]), .QN( ), .S(N$140), .R(n5413), .CK(clk)
    , .D(n5418[130]));
  _HDFF_verplex \B_reg[126] (.Q(B[126]), .QN( ), .S(N$139), .R(n5413), .CK(clk)
    , .D(n5418[129]));
  _HDFF_verplex \B_reg[127] (.Q(B[127]), .QN( ), .S(N$138), .R(n5413), .CK(clk)
    , .D(n5418[128]));
  _HDFF_verplex \B_reg[128] (.Q(B[128]), .QN( ), .S(N$137), .R(n5413), .CK(clk)
    , .D(n5418[127]));
  _HDFF_verplex \B_reg[129] (.Q(B[129]), .QN( ), .S(N$136), .R(n5413), .CK(clk)
    , .D(n5418[126]));
  _HDFF_verplex \B_reg[130] (.Q(B[130]), .QN( ), .S(N$135), .R(n5413), .CK(clk)
    , .D(n5418[125]));
  _HDFF_verplex \B_reg[131] (.Q(B[131]), .QN( ), .S(N$134), .R(n5413), .CK(clk)
    , .D(n5418[124]));
  _HDFF_verplex \B_reg[132] (.Q(B[132]), .QN( ), .S(N$133), .R(n5413), .CK(clk)
    , .D(n5418[123]));
  _HDFF_verplex \B_reg[133] (.Q(B[133]), .QN( ), .S(N$132), .R(n5413), .CK(clk)
    , .D(n5418[122]));
  _HDFF_verplex \B_reg[134] (.Q(B[134]), .QN( ), .S(N$131), .R(n5413), .CK(clk)
    , .D(n5418[121]));
  _HDFF_verplex \B_reg[135] (.Q(B[135]), .QN( ), .S(N$130), .R(n5413), .CK(clk)
    , .D(n5418[120]));
  _HDFF_verplex \B_reg[136] (.Q(B[136]), .QN( ), .S(N$129), .R(n5413), .CK(clk)
    , .D(n5418[119]));
  _HDFF_verplex \B_reg[137] (.Q(B[137]), .QN( ), .S(N$128), .R(n5413), .CK(clk)
    , .D(n5418[118]));
  _HDFF_verplex \B_reg[138] (.Q(B[138]), .QN( ), .S(N$127), .R(n5413), .CK(clk)
    , .D(n5418[117]));
  _HDFF_verplex \B_reg[139] (.Q(B[139]), .QN( ), .S(N$126), .R(n5413), .CK(clk)
    , .D(n5418[116]));
  _HDFF_verplex \B_reg[140] (.Q(B[140]), .QN( ), .S(N$125), .R(n5413), .CK(clk)
    , .D(n5418[115]));
  _HDFF_verplex \B_reg[141] (.Q(B[141]), .QN( ), .S(N$124), .R(n5413), .CK(clk)
    , .D(n5418[114]));
  _HDFF_verplex \B_reg[142] (.Q(B[142]), .QN( ), .S(N$123), .R(n5413), .CK(clk)
    , .D(n5418[113]));
  _HDFF_verplex \B_reg[143] (.Q(B[143]), .QN( ), .S(N$122), .R(n5413), .CK(clk)
    , .D(n5418[112]));
  _HDFF_verplex \B_reg[144] (.Q(B[144]), .QN( ), .S(N$121), .R(n5413), .CK(clk)
    , .D(n5418[111]));
  _HDFF_verplex \B_reg[145] (.Q(B[145]), .QN( ), .S(N$120), .R(n5413), .CK(clk)
    , .D(n5418[110]));
  _HDFF_verplex \B_reg[146] (.Q(B[146]), .QN( ), .S(N$119), .R(n5413), .CK(clk)
    , .D(n5418[109]));
  _HDFF_verplex \B_reg[147] (.Q(B[147]), .QN( ), .S(N$118), .R(n5413), .CK(clk)
    , .D(n5418[108]));
  _HDFF_verplex \B_reg[148] (.Q(B[148]), .QN( ), .S(N$117), .R(n5413), .CK(clk)
    , .D(n5418[107]));
  _HDFF_verplex \B_reg[149] (.Q(B[149]), .QN( ), .S(N$116), .R(n5413), .CK(clk)
    , .D(n5418[106]));
  _HDFF_verplex \B_reg[150] (.Q(B[150]), .QN( ), .S(N$115), .R(n5413), .CK(clk)
    , .D(n5418[105]));
  _HDFF_verplex \B_reg[151] (.Q(B[151]), .QN( ), .S(N$114), .R(n5413), .CK(clk)
    , .D(n5418[104]));
  _HDFF_verplex \B_reg[152] (.Q(B[152]), .QN( ), .S(N$113), .R(n5413), .CK(clk)
    , .D(n5418[103]));
  _HDFF_verplex \B_reg[153] (.Q(B[153]), .QN( ), .S(N$112), .R(n5413), .CK(clk)
    , .D(n5418[102]));
  _HDFF_verplex \B_reg[154] (.Q(B[154]), .QN( ), .S(N$111), .R(n5413), .CK(clk)
    , .D(n5418[101]));
  _HDFF_verplex \B_reg[155] (.Q(B[155]), .QN( ), .S(N$110), .R(n5413), .CK(clk)
    , .D(n5418[100]));
  _HDFF_verplex \B_reg[156] (.Q(B[156]), .QN( ), .S(N$109), .R(n5413), .CK(clk)
    , .D(n5418[99]));
  _HDFF_verplex \B_reg[157] (.Q(B[157]), .QN( ), .S(N$108), .R(n5413), .CK(clk)
    , .D(n5418[98]));
  _HDFF_verplex \B_reg[158] (.Q(B[158]), .QN( ), .S(N$107), .R(n5413), .CK(clk)
    , .D(n5418[97]));
  _HDFF_verplex \B_reg[159] (.Q(B[159]), .QN( ), .S(N$106), .R(n5413), .CK(clk)
    , .D(n5418[96]));
  _HDFF_verplex \B_reg[160] (.Q(B[160]), .QN( ), .S(N$105), .R(n5413), .CK(clk)
    , .D(n5418[95]));
  _HDFF_verplex \B_reg[161] (.Q(B[161]), .QN( ), .S(N$104), .R(n5413), .CK(clk)
    , .D(n5418[94]));
  _HDFF_verplex \B_reg[162] (.Q(B[162]), .QN( ), .S(N$103), .R(n5413), .CK(clk)
    , .D(n5418[93]));
  _HDFF_verplex \B_reg[163] (.Q(B[163]), .QN( ), .S(N$102), .R(n5413), .CK(clk)
    , .D(n5418[92]));
  _HDFF_verplex \B_reg[164] (.Q(B[164]), .QN( ), .S(N$101), .R(n5413), .CK(clk)
    , .D(n5418[91]));
  _HDFF_verplex \B_reg[165] (.Q(B[165]), .QN( ), .S(N$100), .R(n5413), .CK(clk)
    , .D(n5418[90]));
  _HDFF_verplex \B_reg[166] (.Q(B[166]), .QN( ), .S(N$99), .R(n5413), .CK(clk)
    , .D(n5418[89]));
  _HDFF_verplex \B_reg[167] (.Q(B[167]), .QN( ), .S(N$98), .R(n5413), .CK(clk)
    , .D(n5418[88]));
  _HDFF_verplex \B_reg[168] (.Q(B[168]), .QN( ), .S(N$97), .R(n5413), .CK(clk)
    , .D(n5418[87]));
  _HDFF_verplex \B_reg[169] (.Q(B[169]), .QN( ), .S(N$96), .R(n5413), .CK(clk)
    , .D(n5418[86]));
  _HDFF_verplex \B_reg[170] (.Q(B[170]), .QN( ), .S(N$95), .R(n5413), .CK(clk)
    , .D(n5418[85]));
  _HDFF_verplex \B_reg[171] (.Q(B[171]), .QN( ), .S(N$94), .R(n5413), .CK(clk)
    , .D(n5418[84]));
  _HDFF_verplex \B_reg[172] (.Q(B[172]), .QN( ), .S(N$93), .R(n5413), .CK(clk)
    , .D(n5418[83]));
  _HDFF_verplex \B_reg[173] (.Q(B[173]), .QN( ), .S(N$92), .R(n5413), .CK(clk)
    , .D(n5418[82]));
  _HDFF_verplex \B_reg[174] (.Q(B[174]), .QN( ), .S(N$91), .R(n5413), .CK(clk)
    , .D(n5418[81]));
  _HDFF_verplex \B_reg[175] (.Q(B[175]), .QN( ), .S(N$90), .R(n5413), .CK(clk)
    , .D(n5418[80]));
  _HDFF_verplex \B_reg[176] (.Q(B[176]), .QN( ), .S(N$89), .R(n5413), .CK(clk)
    , .D(n5418[79]));
  _HDFF_verplex \B_reg[177] (.Q(B[177]), .QN( ), .S(N$88), .R(n5413), .CK(clk)
    , .D(n5418[78]));
  _HDFF_verplex \B_reg[178] (.Q(B[178]), .QN( ), .S(N$87), .R(n5413), .CK(clk)
    , .D(n5418[77]));
  _HDFF_verplex \B_reg[179] (.Q(B[179]), .QN( ), .S(N$86), .R(n5413), .CK(clk)
    , .D(n5418[76]));
  _HDFF_verplex \B_reg[180] (.Q(B[180]), .QN( ), .S(N$85), .R(n5413), .CK(clk)
    , .D(n5418[75]));
  _HDFF_verplex \B_reg[181] (.Q(B[181]), .QN( ), .S(N$84), .R(n5413), .CK(clk)
    , .D(n5418[74]));
  _HDFF_verplex \B_reg[182] (.Q(B[182]), .QN( ), .S(N$83), .R(n5413), .CK(clk)
    , .D(n5418[73]));
  _HDFF_verplex \B_reg[183] (.Q(B[183]), .QN( ), .S(N$82), .R(n5413), .CK(clk)
    , .D(n5418[72]));
  _HDFF_verplex \B_reg[184] (.Q(B[184]), .QN( ), .S(N$81), .R(n5413), .CK(clk)
    , .D(n5418[71]));
  _HDFF_verplex \B_reg[185] (.Q(B[185]), .QN( ), .S(N$80), .R(n5413), .CK(clk)
    , .D(n5418[70]));
  _HDFF_verplex \B_reg[186] (.Q(B[186]), .QN( ), .S(N$79), .R(n5413), .CK(clk)
    , .D(n5418[69]));
  _HDFF_verplex \B_reg[187] (.Q(B[187]), .QN( ), .S(N$78), .R(n5413), .CK(clk)
    , .D(n5418[68]));
  _HDFF_verplex \B_reg[188] (.Q(B[188]), .QN( ), .S(N$77), .R(n5413), .CK(clk)
    , .D(n5418[67]));
  _HDFF_verplex \B_reg[189] (.Q(B[189]), .QN( ), .S(N$76), .R(n5413), .CK(clk)
    , .D(n5418[66]));
  _HDFF_verplex \B_reg[190] (.Q(B[190]), .QN( ), .S(N$75), .R(n5413), .CK(clk)
    , .D(n5418[65]));
  _HDFF_verplex \B_reg[191] (.Q(B[191]), .QN( ), .S(N$74), .R(n5413), .CK(clk)
    , .D(n5418[64]));
  _HDFF_verplex \B_reg[192] (.Q(B[192]), .QN( ), .S(N$73), .R(n5413), .CK(clk)
    , .D(n5418[63]));
  _HDFF_verplex \B_reg[193] (.Q(B[193]), .QN( ), .S(N$72), .R(n5413), .CK(clk)
    , .D(n5418[62]));
  _HDFF_verplex \B_reg[194] (.Q(B[194]), .QN( ), .S(N$71), .R(n5413), .CK(clk)
    , .D(n5418[61]));
  _HDFF_verplex \B_reg[195] (.Q(B[195]), .QN( ), .S(N$70), .R(n5413), .CK(clk)
    , .D(n5418[60]));
  _HDFF_verplex \B_reg[196] (.Q(B[196]), .QN( ), .S(N$69), .R(n5413), .CK(clk)
    , .D(n5418[59]));
  _HDFF_verplex \B_reg[197] (.Q(B[197]), .QN( ), .S(N$68), .R(n5413), .CK(clk)
    , .D(n5418[58]));
  _HDFF_verplex \B_reg[198] (.Q(B[198]), .QN( ), .S(N$67), .R(n5413), .CK(clk)
    , .D(n5418[57]));
  _HDFF_verplex \B_reg[199] (.Q(B[199]), .QN( ), .S(N$66), .R(n5413), .CK(clk)
    , .D(n5418[56]));
  _HDFF_verplex \B_reg[200] (.Q(B[200]), .QN( ), .S(N$65), .R(n5413), .CK(clk)
    , .D(n5418[55]));
  _HDFF_verplex \B_reg[201] (.Q(B[201]), .QN( ), .S(N$64), .R(n5413), .CK(clk)
    , .D(n5418[54]));
  _HDFF_verplex \B_reg[202] (.Q(B[202]), .QN( ), .S(N$63), .R(n5413), .CK(clk)
    , .D(n5418[53]));
  _HDFF_verplex \B_reg[203] (.Q(B[203]), .QN( ), .S(N$62), .R(n5413), .CK(clk)
    , .D(n5418[52]));
  _HDFF_verplex \B_reg[204] (.Q(B[204]), .QN( ), .S(N$61), .R(n5413), .CK(clk)
    , .D(n5418[51]));
  _HDFF_verplex \B_reg[205] (.Q(B[205]), .QN( ), .S(N$60), .R(n5413), .CK(clk)
    , .D(n5418[50]));
  _HDFF_verplex \B_reg[206] (.Q(B[206]), .QN( ), .S(N$59), .R(n5413), .CK(clk)
    , .D(n5418[49]));
  _HDFF_verplex \B_reg[207] (.Q(B[207]), .QN( ), .S(N$58), .R(n5413), .CK(clk)
    , .D(n5418[48]));
  _HDFF_verplex \B_reg[208] (.Q(B[208]), .QN( ), .S(N$57), .R(n5413), .CK(clk)
    , .D(n5418[47]));
  _HDFF_verplex \B_reg[209] (.Q(B[209]), .QN( ), .S(N$56), .R(n5413), .CK(clk)
    , .D(n5418[46]));
  _HDFF_verplex \B_reg[210] (.Q(B[210]), .QN( ), .S(N$55), .R(n5413), .CK(clk)
    , .D(n5418[45]));
  _HDFF_verplex \B_reg[211] (.Q(B[211]), .QN( ), .S(N$54), .R(n5413), .CK(clk)
    , .D(n5418[44]));
  _HDFF_verplex \B_reg[212] (.Q(B[212]), .QN( ), .S(N$53), .R(n5413), .CK(clk)
    , .D(n5418[43]));
  _HDFF_verplex \B_reg[213] (.Q(B[213]), .QN( ), .S(N$52), .R(n5413), .CK(clk)
    , .D(n5418[42]));
  _HDFF_verplex \B_reg[214] (.Q(B[214]), .QN( ), .S(N$51), .R(n5413), .CK(clk)
    , .D(n5418[41]));
  _HDFF_verplex \B_reg[215] (.Q(B[215]), .QN( ), .S(N$50), .R(n5413), .CK(clk)
    , .D(n5418[40]));
  _HDFF_verplex \B_reg[216] (.Q(B[216]), .QN( ), .S(N$49), .R(n5413), .CK(clk)
    , .D(n5418[39]));
  _HDFF_verplex \B_reg[217] (.Q(B[217]), .QN( ), .S(N$48), .R(n5413), .CK(clk)
    , .D(n5418[38]));
  _HDFF_verplex \B_reg[218] (.Q(B[218]), .QN( ), .S(N$47), .R(n5413), .CK(clk)
    , .D(n5418[37]));
  _HDFF_verplex \B_reg[219] (.Q(B[219]), .QN( ), .S(N$46), .R(n5413), .CK(clk)
    , .D(n5418[36]));
  _HDFF_verplex \B_reg[220] (.Q(B[220]), .QN( ), .S(N$45), .R(n5413), .CK(clk)
    , .D(n5418[35]));
  _HDFF_verplex \B_reg[221] (.Q(B[221]), .QN( ), .S(N$44), .R(n5413), .CK(clk)
    , .D(n5418[34]));
  _HDFF_verplex \B_reg[222] (.Q(B[222]), .QN( ), .S(N$43), .R(n5413), .CK(clk)
    , .D(n5418[33]));
  _HDFF_verplex \B_reg[223] (.Q(B[223]), .QN( ), .S(N$42), .R(n5413), .CK(clk)
    , .D(n5418[32]));
  _HDFF_verplex \B_reg[224] (.Q(B[224]), .QN( ), .S(N$41), .R(n5413), .CK(clk)
    , .D(n5418[31]));
  _HDFF_verplex \B_reg[225] (.Q(B[225]), .QN( ), .S(N$40), .R(n5413), .CK(clk)
    , .D(n5418[30]));
  _HDFF_verplex \B_reg[226] (.Q(B[226]), .QN( ), .S(N$39), .R(n5413), .CK(clk)
    , .D(n5418[29]));
  _HDFF_verplex \B_reg[227] (.Q(B[227]), .QN( ), .S(N$38), .R(n5413), .CK(clk)
    , .D(n5418[28]));
  _HDFF_verplex \B_reg[228] (.Q(B[228]), .QN( ), .S(N$37), .R(n5413), .CK(clk)
    , .D(n5418[27]));
  _HDFF_verplex \B_reg[229] (.Q(B[229]), .QN( ), .S(N$36), .R(n5413), .CK(clk)
    , .D(n5418[26]));
  _HDFF_verplex \B_reg[230] (.Q(B[230]), .QN( ), .S(N$35), .R(n5413), .CK(clk)
    , .D(n5418[25]));
  _HDFF_verplex \B_reg[231] (.Q(B[231]), .QN( ), .S(N$34), .R(n5413), .CK(clk)
    , .D(n5418[24]));
  _HDFF_verplex \B_reg[232] (.Q(B[232]), .QN( ), .S(N$33), .R(n5413), .CK(clk)
    , .D(n5418[23]));
  _HDFF_verplex \B_reg[233] (.Q(B[233]), .QN( ), .S(N$32), .R(n5413), .CK(clk)
    , .D(n5418[22]));
  _HDFF_verplex \B_reg[234] (.Q(B[234]), .QN( ), .S(N$31), .R(n5413), .CK(clk)
    , .D(n5418[21]));
  _HDFF_verplex \B_reg[235] (.Q(B[235]), .QN( ), .S(N$30), .R(n5413), .CK(clk)
    , .D(n5418[20]));
  _HDFF_verplex \B_reg[236] (.Q(B[236]), .QN( ), .S(N$29), .R(n5413), .CK(clk)
    , .D(n5418[19]));
  _HDFF_verplex \B_reg[237] (.Q(B[237]), .QN( ), .S(N$28), .R(n5413), .CK(clk)
    , .D(n5418[18]));
  _HDFF_verplex \B_reg[238] (.Q(B[238]), .QN( ), .S(N$27), .R(n5413), .CK(clk)
    , .D(n5418[17]));
  _HDFF_verplex \B_reg[239] (.Q(B[239]), .QN( ), .S(N$26), .R(n5413), .CK(clk)
    , .D(n5418[16]));
  _HDFF_verplex \B_reg[240] (.Q(B[240]), .QN( ), .S(N$25), .R(n5413), .CK(clk)
    , .D(n5418[15]));
  _HDFF_verplex \B_reg[241] (.Q(B[241]), .QN( ), .S(N$24), .R(n5413), .CK(clk)
    , .D(n5418[14]));
  _HDFF_verplex \B_reg[242] (.Q(B[242]), .QN( ), .S(N$23), .R(n5413), .CK(clk)
    , .D(n5418[13]));
  _HDFF_verplex \B_reg[243] (.Q(B[243]), .QN( ), .S(N$22), .R(n5413), .CK(clk)
    , .D(n5418[12]));
  _HDFF_verplex \B_reg[244] (.Q(B[244]), .QN( ), .S(N$21), .R(n5413), .CK(clk)
    , .D(n5418[11]));
  _HDFF_verplex \B_reg[245] (.Q(B[245]), .QN( ), .S(N$20), .R(n5413), .CK(clk)
    , .D(n5418[10]));
  _HDFF_verplex \B_reg[246] (.Q(B[246]), .QN( ), .S(N$19), .R(n5413), .CK(clk)
    , .D(n5418[9]));
  _HDFF_verplex \B_reg[247] (.Q(B[247]), .QN( ), .S(N$18), .R(n5413), .CK(clk)
    , .D(n5418[8]));
  _HDFF_verplex \B_reg[248] (.Q(B[248]), .QN( ), .S(N$17), .R(n5413), .CK(clk)
    , .D(n5418[7]));
  _HDFF_verplex \B_reg[249] (.Q(B[249]), .QN( ), .S(N$16), .R(n5413), .CK(clk)
    , .D(n5418[6]));
  _HDFF_verplex \B_reg[250] (.Q(B[250]), .QN( ), .S(N$15), .R(n5413), .CK(clk)
    , .D(n5418[5]));
  _HDFF_verplex \B_reg[251] (.Q(B[251]), .QN( ), .S(N$14), .R(n5413), .CK(clk)
    , .D(n5418[4]));
  _HDFF_verplex \B_reg[252] (.Q(B[252]), .QN( ), .S(N$13), .R(n5413), .CK(clk)
    , .D(n5418[3]));
  _HDFF_verplex \B_reg[253] (.Q(B[253]), .QN( ), .S(N$12), .R(n5413), .CK(clk)
    , .D(n5418[2]));
  _HDFF_verplex \B_reg[254] (.Q(B[254]), .QN( ), .S(N$11), .R(n5413), .CK(clk)
    , .D(n5418[1]));
  _HDFF_verplex \B_reg[255] (.Q(B[255]), .QN( ), .S(N$10), .R(n5413), .CK(clk)
    , .D(n5418[0]));
  VDW_WMUX256 U$5321(.Z({ n5418[255:0] }), .A({ in[0:127] ,  B[128:255] }), .B({ B[0:127] ,  in[0:127] }), .S(updown));
  not U$5322(n5413, rst_n);
  assign out[179] = \out_reg[19] [8];
  assign out[178] = \out_reg[19] [7];
  assign out[177] = \out_reg[19] [6];
  assign out[176] = \out_reg[19] [5];
  assign out[175] = \out_reg[19] [4];
  assign out[174] = \out_reg[19] [3];
  assign out[173] = \out_reg[19] [2];
  assign out[172] = \out_reg[19] [1];
  assign out[171] = \out_reg[19] [0];
  assign out[170] = \out_reg[18] [8];
  assign out[169] = \out_reg[18] [7];
  assign out[168] = \out_reg[18] [6];
  assign out[167] = \out_reg[18] [5];
  assign out[166] = \out_reg[18] [4];
  assign out[165] = \out_reg[18] [3];
  assign out[164] = \out_reg[18] [2];
  assign out[163] = \out_reg[18] [1];
  assign out[162] = \out_reg[18] [0];
  assign out[161] = \out_reg[17] [8];
  assign out[160] = \out_reg[17] [7];
  assign out[159] = \out_reg[17] [6];
  assign out[158] = \out_reg[17] [5];
  assign out[157] = \out_reg[17] [4];
  assign out[156] = \out_reg[17] [3];
  assign out[155] = \out_reg[17] [2];
  assign out[154] = \out_reg[17] [1];
  assign out[153] = \out_reg[17] [0];
  assign out[152] = \out_reg[16] [8];
  assign out[151] = \out_reg[16] [7];
  assign out[150] = \out_reg[16] [6];
  assign out[149] = \out_reg[16] [5];
  assign out[148] = \out_reg[16] [4];
  assign out[147] = \out_reg[16] [3];
  assign out[146] = \out_reg[16] [2];
  assign out[145] = \out_reg[16] [1];
  assign out[144] = \out_reg[16] [0];
  assign out[143] = \out_reg[15] [8];
  assign out[142] = \out_reg[15] [7];
  assign out[141] = \out_reg[15] [6];
  assign out[140] = \out_reg[15] [5];
  assign out[139] = \out_reg[15] [4];
  assign out[138] = \out_reg[15] [3];
  assign out[137] = \out_reg[15] [2];
  assign out[136] = \out_reg[15] [1];
  assign out[135] = \out_reg[15] [0];
  assign out[134] = \out_reg[14] [8];
  assign out[133] = \out_reg[14] [7];
  assign out[132] = \out_reg[14] [6];
  assign out[131] = \out_reg[14] [5];
  assign out[130] = \out_reg[14] [4];
  assign out[129] = \out_reg[14] [3];
  assign out[128] = \out_reg[14] [2];
  assign out[127] = \out_reg[14] [1];
  assign out[126] = \out_reg[14] [0];
  assign out[125] = \out_reg[13] [8];
  assign out[124] = \out_reg[13] [7];
  assign out[123] = \out_reg[13] [6];
  assign out[122] = \out_reg[13] [5];
  assign out[121] = \out_reg[13] [4];
  assign out[120] = \out_reg[13] [3];
  assign out[119] = \out_reg[13] [2];
  assign out[118] = \out_reg[13] [1];
  assign out[117] = \out_reg[13] [0];
  assign out[116] = \out_reg[12] [8];
  assign out[115] = \out_reg[12] [7];
  assign out[114] = \out_reg[12] [6];
  assign out[113] = \out_reg[12] [5];
  assign out[112] = \out_reg[12] [4];
  assign out[111] = \out_reg[12] [3];
  assign out[110] = \out_reg[12] [2];
  assign out[109] = \out_reg[12] [1];
  assign out[108] = \out_reg[12] [0];
  assign out[107] = \out_reg[11] [8];
  assign out[106] = \out_reg[11] [7];
  assign out[105] = \out_reg[11] [6];
  assign out[104] = \out_reg[11] [5];
  assign out[103] = \out_reg[11] [4];
  assign out[102] = \out_reg[11] [3];
  assign out[101] = \out_reg[11] [2];
  assign out[100] = \out_reg[11] [1];
  assign out[99] = \out_reg[11] [0];
  assign out[98] = \out_reg[10] [8];
  assign out[97] = \out_reg[10] [7];
  assign out[96] = \out_reg[10] [6];
  assign out[95] = \out_reg[10] [5];
  assign out[94] = \out_reg[10] [4];
  assign out[93] = \out_reg[10] [3];
  assign out[92] = \out_reg[10] [2];
  assign out[91] = \out_reg[10] [1];
  assign out[90] = \out_reg[10] [0];
  assign out[89] = \out_reg[9] [8];
  assign out[88] = \out_reg[9] [7];
  assign out[87] = \out_reg[9] [6];
  assign out[86] = \out_reg[9] [5];
  assign out[85] = \out_reg[9] [4];
  assign out[84] = \out_reg[9] [3];
  assign out[83] = \out_reg[9] [2];
  assign out[82] = \out_reg[9] [1];
  assign out[81] = \out_reg[9] [0];
  assign out[80] = \out_reg[8] [8];
  assign out[79] = \out_reg[8] [7];
  assign out[78] = \out_reg[8] [6];
  assign out[77] = \out_reg[8] [5];
  assign out[76] = \out_reg[8] [4];
  assign out[75] = \out_reg[8] [3];
  assign out[74] = \out_reg[8] [2];
  assign out[73] = \out_reg[8] [1];
  assign out[72] = \out_reg[8] [0];
  assign out[71] = \out_reg[7] [8];
  assign out[70] = \out_reg[7] [7];
  assign out[69] = \out_reg[7] [6];
  assign out[68] = \out_reg[7] [5];
  assign out[67] = \out_reg[7] [4];
  assign out[66] = \out_reg[7] [3];
  assign out[65] = \out_reg[7] [2];
  assign out[64] = \out_reg[7] [1];
  assign out[63] = \out_reg[7] [0];
  assign out[62] = \out_reg[6] [8];
  assign out[61] = \out_reg[6] [7];
  assign out[60] = \out_reg[6] [6];
  assign out[59] = \out_reg[6] [5];
  assign out[58] = \out_reg[6] [4];
  assign out[57] = \out_reg[6] [3];
  assign out[56] = \out_reg[6] [2];
  assign out[55] = \out_reg[6] [1];
  assign out[54] = \out_reg[6] [0];
  assign out[53] = \out_reg[5] [8];
  assign out[52] = \out_reg[5] [7];
  assign out[51] = \out_reg[5] [6];
  assign out[50] = \out_reg[5] [5];
  assign out[49] = \out_reg[5] [4];
  assign out[48] = \out_reg[5] [3];
  assign out[47] = \out_reg[5] [2];
  assign out[46] = \out_reg[5] [1];
  assign out[45] = \out_reg[5] [0];
  assign out[44] = \out_reg[4] [8];
  assign out[43] = \out_reg[4] [7];
  assign out[42] = \out_reg[4] [6];
  assign out[41] = \out_reg[4] [5];
  assign out[40] = \out_reg[4] [4];
  assign out[39] = \out_reg[4] [3];
  assign out[38] = \out_reg[4] [2];
  assign out[37] = \out_reg[4] [1];
  assign out[36] = \out_reg[4] [0];
  assign out[35] = \out_reg[3] [8];
  assign out[34] = \out_reg[3] [7];
  assign out[33] = \out_reg[3] [6];
  assign out[32] = \out_reg[3] [5];
  assign out[31] = \out_reg[3] [4];
  assign out[30] = \out_reg[3] [3];
  assign out[29] = \out_reg[3] [2];
  assign out[28] = \out_reg[3] [1];
  assign out[27] = \out_reg[3] [0];
  assign out[26] = \out_reg[2] [8];
  assign out[25] = \out_reg[2] [7];
  assign out[24] = \out_reg[2] [6];
  assign out[23] = \out_reg[2] [5];
  assign out[22] = \out_reg[2] [4];
  assign out[21] = \out_reg[2] [3];
  assign out[20] = \out_reg[2] [2];
  assign out[19] = \out_reg[2] [1];
  assign out[18] = \out_reg[2] [0];
  assign out[17] = \out_reg[1] [8];
  assign out[16] = \out_reg[1] [7];
  assign out[15] = \out_reg[1] [6];
  assign out[14] = \out_reg[1] [5];
  assign out[13] = \out_reg[1] [4];
  assign out[12] = \out_reg[1] [3];
  assign out[11] = \out_reg[1] [2];
  assign out[10] = \out_reg[1] [1];
  assign out[9] = \out_reg[1] [0];
  assign out[8] = \out_reg[0] [8];
  assign out[7] = \out_reg[0] [7];
  assign out[6] = \out_reg[0] [6];
  assign out[5] = \out_reg[0] [5];
  assign out[4] = \out_reg[0] [4];
  assign out[3] = \out_reg[0] [3];
  assign out[2] = \out_reg[0] [2];
  assign out[1] = \out_reg[0] [1];
  assign out[0] = \out_reg[0] [0];
  ReLU_10bit \dot_product_and_ReLU[0].relu_inst (.in_data({ \final_sums[0] [9:0] }), .out_data({ \out_sig[0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[1] [4:0] }), .sum({ \level_1_sums[0][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[3] [4:0] }), .sum({ \level_1_sums[0][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[0][1] [5:0] }),
     .b({ \level_1_sums[0][0] [5:0] }), .sum({ \level_2_sums[0][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[5] [4:0] }), .sum({ \level_1_sums[0][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[7] [4:0] }), .sum({ \level_1_sums[0][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[0][3] [5:0] }),
     .b({ \level_1_sums[0][2] [5:0] }), .sum({ \level_2_sums[0][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[0][1] [6:0] }),
     .b({ \level_2_sums[0][0] [6:0] }), .sum({ \level_3_sums[0][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[9] [4:0] }), .sum({ \level_1_sums[0][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[11] [4:0] }), .sum({ \level_1_sums[0][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[0][5] [5:0] }),
     .b({ \level_1_sums[0][4] [5:0] }), .sum({ \level_2_sums[0][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[13] [4:0] }), .sum({ \level_1_sums[0][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[15] [4:0] }), .sum({ \level_1_sums[0][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[0][7] [5:0] }),
     .b({ \level_1_sums[0][6] [5:0] }), .sum({ \level_2_sums[0][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[0][3] [6:0] }),
     .b({ \level_2_sums[0][2] [6:0] }), .sum({ \level_3_sums[0][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[0][1] [7:0] }),
     .b({ \level_3_sums[0][0] [7:0] }), .sum({ \level_4_sums[0][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[17] [4:0] }), .sum({ \level_1_sums[0][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[19] [4:0] }), .sum({ \level_1_sums[0][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[0][9] [5:0] }),
     .b({ \level_1_sums[0][8] [5:0] }), .sum({ \level_2_sums[0][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[21] [4:0] }), .sum({ \level_1_sums[0][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[23] [4:0] }), .sum({ \level_1_sums[0][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[0][11] [5:0] }),
     .b({ \level_1_sums[0][10] [5:0] }), .sum({ \level_2_sums[0][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[0][5] [6:0] }),
     .b({ \level_2_sums[0][4] [6:0] }), .sum({ \level_3_sums[0][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[25] [4:0] }), .sum({ \level_1_sums[0][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[27] [4:0] }), .sum({ \level_1_sums[0][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[0][13] [5:0] }),
     .b({ \level_1_sums[0][12] [5:0] }), .sum({ \level_2_sums[0][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[29] [4:0] }), .sum({ \level_1_sums[0][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[31] [4:0] }), .sum({ \level_1_sums[0][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[0][15] [5:0] }),
     .b({ \level_1_sums[0][14] [5:0] }), .sum({ \level_2_sums[0][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[0][7] [6:0] }),
     .b({ \level_2_sums[0][6] [6:0] }), .sum({ \level_3_sums[0][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[0][3] [7:0] }),
     .b({ \level_3_sums[0][2] [7:0] }), .sum({ \level_4_sums[0][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[0][1] [8:0] }),
     .b({ \level_4_sums[0][0] [8:0] }), .sum({ \level_5_sums[0][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[33] [4:0] }), .sum({ \level_1_sums[0][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[35] [4:0] }), .sum({ \level_1_sums[0][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[0][17] [5:0] }),
     .b({ \level_1_sums[0][16] [5:0] }), .sum({ \level_2_sums[0][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[37] [4:0] }), .sum({ \level_1_sums[0][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[39] [4:0] }), .sum({ \level_1_sums[0][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[0][19] [5:0] }),
     .b({ \level_1_sums[0][18] [5:0] }), .sum({ \level_2_sums[0][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[0][9] [6:0] }),
     .b({ \level_2_sums[0][8] [6:0] }), .sum({ \level_3_sums[0][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[41] [4:0] }), .sum({ \level_1_sums[0][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[43] [4:0] }), .sum({ \level_1_sums[0][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[0][21] [5:0] }),
     .b({ \level_1_sums[0][20] [5:0] }), .sum({ \level_2_sums[0][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[45] [4:0] }), .sum({ \level_1_sums[0][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[47] [4:0] }), .sum({ \level_1_sums[0][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[0][23] [5:0] }),
     .b({ \level_1_sums[0][22] [5:0] }), .sum({ \level_2_sums[0][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[0][11] [6:0] }),
     .b({ \level_2_sums[0][10] [6:0] }), .sum({ \level_3_sums[0][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[0][5] [7:0] }),
     .b({ \level_3_sums[0][4] [7:0] }), .sum({ \level_4_sums[0][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[49] [4:0] }), .sum({ \level_1_sums[0][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[51] [4:0] }), .sum({ \level_1_sums[0][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[0][25] [5:0] }),
     .b({ \level_1_sums[0][24] [5:0] }), .sum({ \level_2_sums[0][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[53] [4:0] }), .sum({ \level_1_sums[0][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[55] [4:0] }), .sum({ \level_1_sums[0][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[0][27] [5:0] }),
     .b({ \level_1_sums[0][26] [5:0] }), .sum({ \level_2_sums[0][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[0][13] [6:0] }),
     .b({ \level_2_sums[0][12] [6:0] }), .sum({ \level_3_sums[0][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[57] [4:0] }), .sum({ \level_1_sums[0][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[59] [4:0] }), .sum({ \level_1_sums[0][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[0][29] [5:0] }),
     .b({ \level_1_sums[0][28] [5:0] }), .sum({ \level_2_sums[0][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[61] [4:0] }), .sum({ \level_1_sums[0][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[63] [4:0] }), .sum({ \level_1_sums[0][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[0][31] [5:0] }),
     .b({ \level_1_sums[0][30] [5:0] }), .sum({ \level_2_sums[0][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[0][15] [6:0] }),
     .b({ \level_2_sums[0][14] [6:0] }), .sum({ \level_3_sums[0][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[0][7] [7:0] }),
     .b({ \level_3_sums[0][6] [7:0] }), .sum({ \level_4_sums[0][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[0][3] [8:0] }),
     .b({ \level_4_sums[0][2] [8:0] }), .sum({ \level_5_sums[0][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[0][1] [9:0] }),
     .b({ \level_5_sums[0][0] [9:0] }), .sum({ \level_6_sums[0][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[65] [4:0] }), .sum({ \level_1_sums[0][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[67] [4:0] }), .sum({ \level_1_sums[0][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[0][33] [5:0] }),
     .b({ \level_1_sums[0][32] [5:0] }), .sum({ \level_2_sums[0][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[69] [4:0] }), .sum({ \level_1_sums[0][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[71] [4:0] }), .sum({ \level_1_sums[0][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[0][35] [5:0] }),
     .b({ \level_1_sums[0][34] [5:0] }), .sum({ \level_2_sums[0][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[0][17] [6:0] }),
     .b({ \level_2_sums[0][16] [6:0] }), .sum({ \level_3_sums[0][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[73] [4:0] }), .sum({ \level_1_sums[0][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[75] [4:0] }), .sum({ \level_1_sums[0][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[0][37] [5:0] }),
     .b({ \level_1_sums[0][36] [5:0] }), .sum({ \level_2_sums[0][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[77] [4:0] }), .sum({ \level_1_sums[0][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[79] [4:0] }), .sum({ \level_1_sums[0][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[0][39] [5:0] }),
     .b({ \level_1_sums[0][38] [5:0] }), .sum({ \level_2_sums[0][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[0][19] [6:0] }),
     .b({ \level_2_sums[0][18] [6:0] }), .sum({ \level_3_sums[0][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[0][9] [7:0] }),
     .b({ \level_3_sums[0][8] [7:0] }), .sum({ \level_4_sums[0][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[81] [4:0] }), .sum({ \level_1_sums[0][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[83] [4:0] }), .sum({ \level_1_sums[0][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[0][41] [5:0] }),
     .b({ \level_1_sums[0][40] [5:0] }), .sum({ \level_2_sums[0][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[85] [4:0] }), .sum({ \level_1_sums[0][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[87] [4:0] }), .sum({ \level_1_sums[0][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[0][43] [5:0] }),
     .b({ \level_1_sums[0][42] [5:0] }), .sum({ \level_2_sums[0][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[0][21] [6:0] }),
     .b({ \level_2_sums[0][20] [6:0] }), .sum({ \level_3_sums[0][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[89] [4:0] }), .sum({ \level_1_sums[0][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[91] [4:0] }), .sum({ \level_1_sums[0][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[0][45] [5:0] }),
     .b({ \level_1_sums[0][44] [5:0] }), .sum({ \level_2_sums[0][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[93] [4:0] }), .sum({ \level_1_sums[0][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[95] [4:0] }), .sum({ \level_1_sums[0][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[0][47] [5:0] }),
     .b({ \level_1_sums[0][46] [5:0] }), .sum({ \level_2_sums[0][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[0][23] [6:0] }),
     .b({ \level_2_sums[0][22] [6:0] }), .sum({ \level_3_sums[0][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[0][11] [7:0] }),
     .b({ \level_3_sums[0][10] [7:0] }), .sum({ \level_4_sums[0][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[0][5] [8:0] }),
     .b({ \level_4_sums[0][4] [8:0] }), .sum({ \level_5_sums[0][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[97] [4:0] }), .sum({ \level_1_sums[0][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[99] [4:0] }), .sum({ \level_1_sums[0][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[0][49] [5:0] }),
     .b({ \level_1_sums[0][48] [5:0] }), .sum({ \level_2_sums[0][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[101] [4:0] }), .sum({ \level_1_sums[0][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[103] [4:0] }), .sum({ \level_1_sums[0][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[0][51] [5:0] }),
     .b({ \level_1_sums[0][50] [5:0] }), .sum({ \level_2_sums[0][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[0][25] [6:0] }),
     .b({ \level_2_sums[0][24] [6:0] }), .sum({ \level_3_sums[0][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[105] [4:0] }), .sum({ \level_1_sums[0][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[107] [4:0] }), .sum({ \level_1_sums[0][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[0][53] [5:0] }),
     .b({ \level_1_sums[0][52] [5:0] }), .sum({ \level_2_sums[0][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[109] [4:0] }), .sum({ \level_1_sums[0][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[111] [4:0] }), .sum({ \level_1_sums[0][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[0][55] [5:0] }),
     .b({ \level_1_sums[0][54] [5:0] }), .sum({ \level_2_sums[0][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[0][27] [6:0] }),
     .b({ \level_2_sums[0][26] [6:0] }), .sum({ \level_3_sums[0][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[0][13] [7:0] }),
     .b({ \level_3_sums[0][12] [7:0] }), .sum({ \level_4_sums[0][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[113] [4:0] }), .sum({ \level_1_sums[0][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[115] [4:0] }), .sum({ \level_1_sums[0][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[0][57] [5:0] }),
     .b({ \level_1_sums[0][56] [5:0] }), .sum({ \level_2_sums[0][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[117] [4:0] }), .sum({ \level_1_sums[0][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[119] [4:0] }), .sum({ \level_1_sums[0][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[0][59] [5:0] }),
     .b({ \level_1_sums[0][58] [5:0] }), .sum({ \level_2_sums[0][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[0][29] [6:0] }),
     .b({ \level_2_sums[0][28] [6:0] }), .sum({ \level_3_sums[0][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[121] [4:0] }), .sum({ \level_1_sums[0][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[123] [4:0] }), .sum({ \level_1_sums[0][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[0][61] [5:0] }),
     .b({ \level_1_sums[0][60] [5:0] }), .sum({ \level_2_sums[0][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[125] [4:0] }), .sum({ \level_1_sums[0][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[127] [4:0] }), .sum({ \level_1_sums[0][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[0][63] [5:0] }),
     .b({ \level_1_sums[0][62] [5:0] }), .sum({ \level_2_sums[0][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[0][31] [6:0] }),
     .b({ \level_2_sums[0][30] [6:0] }), .sum({ \level_3_sums[0][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[0][15] [7:0] }),
     .b({ \level_3_sums[0][14] [7:0] }), .sum({ \level_4_sums[0][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[0][7] [8:0] }),
     .b({ \level_4_sums[0][6] [8:0] }), .sum({ \level_5_sums[0][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[0][3] [9:0] }),
     .b({ \level_5_sums[0][2] [9:0] }), .sum({ \level_6_sums[0][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[0][1] [9:0] }),
     .b({ \level_6_sums[0][0] [9:0] }), .sum({ \level_7_sums[0][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[129] [4:0] }), .sum({ \level_1_sums[0][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[131] [4:0] }), .sum({ \level_1_sums[0][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[0][65] [5:0] }),
     .b({ \level_1_sums[0][64] [5:0] }), .sum({ \level_2_sums[0][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[133] [4:0] }), .sum({ \level_1_sums[0][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[135] [4:0] }), .sum({ \level_1_sums[0][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[0][67] [5:0] }),
     .b({ \level_1_sums[0][66] [5:0] }), .sum({ \level_2_sums[0][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[0][33] [6:0] }),
     .b({ \level_2_sums[0][32] [6:0] }), .sum({ \level_3_sums[0][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[137] [4:0] }), .sum({ \level_1_sums[0][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[139] [4:0] }), .sum({ \level_1_sums[0][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[0][69] [5:0] }),
     .b({ \level_1_sums[0][68] [5:0] }), .sum({ \level_2_sums[0][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[141] [4:0] }), .sum({ \level_1_sums[0][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[143] [4:0] }), .sum({ \level_1_sums[0][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[0][71] [5:0] }),
     .b({ \level_1_sums[0][70] [5:0] }), .sum({ \level_2_sums[0][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[0][35] [6:0] }),
     .b({ \level_2_sums[0][34] [6:0] }), .sum({ \level_3_sums[0][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[0][17] [7:0] }),
     .b({ \level_3_sums[0][16] [7:0] }), .sum({ \level_4_sums[0][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[145] [4:0] }), .sum({ \level_1_sums[0][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[147] [4:0] }), .sum({ \level_1_sums[0][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[0][73] [5:0] }),
     .b({ \level_1_sums[0][72] [5:0] }), .sum({ \level_2_sums[0][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[149] [4:0] }), .sum({ \level_1_sums[0][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[151] [4:0] }), .sum({ \level_1_sums[0][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[0][75] [5:0] }),
     .b({ \level_1_sums[0][74] [5:0] }), .sum({ \level_2_sums[0][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[0][37] [6:0] }),
     .b({ \level_2_sums[0][36] [6:0] }), .sum({ \level_3_sums[0][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[153] [4:0] }), .sum({ \level_1_sums[0][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[155] [4:0] }), .sum({ \level_1_sums[0][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[0][77] [5:0] }),
     .b({ \level_1_sums[0][76] [5:0] }), .sum({ \level_2_sums[0][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[157] [4:0] }), .sum({ \level_1_sums[0][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[159] [4:0] }), .sum({ \level_1_sums[0][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[0][79] [5:0] }),
     .b({ \level_1_sums[0][78] [5:0] }), .sum({ \level_2_sums[0][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[0][39] [6:0] }),
     .b({ \level_2_sums[0][38] [6:0] }), .sum({ \level_3_sums[0][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[0][19] [7:0] }),
     .b({ \level_3_sums[0][18] [7:0] }), .sum({ \level_4_sums[0][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[0][9] [8:0] }),
     .b({ \level_4_sums[0][8] [8:0] }), .sum({ \level_5_sums[0][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[161] [4:0] }), .sum({ \level_1_sums[0][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[163] [4:0] }), .sum({ \level_1_sums[0][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[0][81] [5:0] }),
     .b({ \level_1_sums[0][80] [5:0] }), .sum({ \level_2_sums[0][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[165] [4:0] }), .sum({ \level_1_sums[0][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[167] [4:0] }), .sum({ \level_1_sums[0][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[0][83] [5:0] }),
     .b({ \level_1_sums[0][82] [5:0] }), .sum({ \level_2_sums[0][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[0][41] [6:0] }),
     .b({ \level_2_sums[0][40] [6:0] }), .sum({ \level_3_sums[0][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[169] [4:0] }), .sum({ \level_1_sums[0][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[171] [4:0] }), .sum({ \level_1_sums[0][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[0][85] [5:0] }),
     .b({ \level_1_sums[0][84] [5:0] }), .sum({ \level_2_sums[0][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[173] [4:0] }), .sum({ \level_1_sums[0][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[175] [4:0] }), .sum({ \level_1_sums[0][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[0][87] [5:0] }),
     .b({ \level_1_sums[0][86] [5:0] }), .sum({ \level_2_sums[0][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[0][43] [6:0] }),
     .b({ \level_2_sums[0][42] [6:0] }), .sum({ \level_3_sums[0][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[0][21] [7:0] }),
     .b({ \level_3_sums[0][20] [7:0] }), .sum({ \level_4_sums[0][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[177] [4:0] }), .sum({ \level_1_sums[0][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[179] [4:0] }), .sum({ \level_1_sums[0][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[0][89] [5:0] }),
     .b({ \level_1_sums[0][88] [5:0] }), .sum({ \level_2_sums[0][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[181] [4:0] }), .sum({ \level_1_sums[0][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[183] [4:0] }), .sum({ \level_1_sums[0][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[0][91] [5:0] }),
     .b({ \level_1_sums[0][90] [5:0] }), .sum({ \level_2_sums[0][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[0][45] [6:0] }),
     .b({ \level_2_sums[0][44] [6:0] }), .sum({ \level_3_sums[0][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[185] [4:0] }), .sum({ \level_1_sums[0][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[187] [4:0] }), .sum({ \level_1_sums[0][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[0][93] [5:0] }),
     .b({ \level_1_sums[0][92] [5:0] }), .sum({ \level_2_sums[0][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[189] [4:0] }), .sum({ \level_1_sums[0][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[191] [4:0] }), .sum({ \level_1_sums[0][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[0][95] [5:0] }),
     .b({ \level_1_sums[0][94] [5:0] }), .sum({ \level_2_sums[0][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[0][47] [6:0] }),
     .b({ \level_2_sums[0][46] [6:0] }), .sum({ \level_3_sums[0][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[0][23] [7:0] }),
     .b({ \level_3_sums[0][22] [7:0] }), .sum({ \level_4_sums[0][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[0][11] [8:0] }),
     .b({ \level_4_sums[0][10] [8:0] }), .sum({ \level_5_sums[0][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[0][5] [9:0] }),
     .b({ \level_5_sums[0][4] [9:0] }), .sum({ \level_6_sums[0][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[193] [4:0] }), .sum({ \level_1_sums[0][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[195] [4:0] }), .sum({ \level_1_sums[0][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[0][97] [5:0] }),
     .b({ \level_1_sums[0][96] [5:0] }), .sum({ \level_2_sums[0][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[197] [4:0] }), .sum({ \level_1_sums[0][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[199] [4:0] }), .sum({ \level_1_sums[0][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[0][99] [5:0] }),
     .b({ \level_1_sums[0][98] [5:0] }), .sum({ \level_2_sums[0][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[0][49] [6:0] }),
     .b({ \level_2_sums[0][48] [6:0] }), .sum({ \level_3_sums[0][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[201] [4:0] }), .sum({ \level_1_sums[0][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[203] [4:0] }), .sum({ \level_1_sums[0][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[0][101] [5:0] }),
     .b({ \level_1_sums[0][100] [5:0] }), .sum({ \level_2_sums[0][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[205] [4:0] }), .sum({ \level_1_sums[0][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[207] [4:0] }), .sum({ \level_1_sums[0][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[0][103] [5:0] }),
     .b({ \level_1_sums[0][102] [5:0] }), .sum({ \level_2_sums[0][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[0][51] [6:0] }),
     .b({ \level_2_sums[0][50] [6:0] }), .sum({ \level_3_sums[0][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[0][25] [7:0] }),
     .b({ \level_3_sums[0][24] [7:0] }), .sum({ \level_4_sums[0][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[209] [4:0] }), .sum({ \level_1_sums[0][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[211] [4:0] }), .sum({ \level_1_sums[0][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[0][105] [5:0] }),
     .b({ \level_1_sums[0][104] [5:0] }), .sum({ \level_2_sums[0][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[213] [4:0] }), .sum({ \level_1_sums[0][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[215] [4:0] }), .sum({ \level_1_sums[0][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[0][107] [5:0] }),
     .b({ \level_1_sums[0][106] [5:0] }), .sum({ \level_2_sums[0][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[0][53] [6:0] }),
     .b({ \level_2_sums[0][52] [6:0] }), .sum({ \level_3_sums[0][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[217] [4:0] }), .sum({ \level_1_sums[0][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[219] [4:0] }), .sum({ \level_1_sums[0][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[0][109] [5:0] }),
     .b({ \level_1_sums[0][108] [5:0] }), .sum({ \level_2_sums[0][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[221] [4:0] }), .sum({ \level_1_sums[0][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[223] [4:0] }), .sum({ \level_1_sums[0][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[0][111] [5:0] }),
     .b({ \level_1_sums[0][110] [5:0] }), .sum({ \level_2_sums[0][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[0][55] [6:0] }),
     .b({ \level_2_sums[0][54] [6:0] }), .sum({ \level_3_sums[0][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[0][27] [7:0] }),
     .b({ \level_3_sums[0][26] [7:0] }), .sum({ \level_4_sums[0][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[0][13] [8:0] }),
     .b({ \level_4_sums[0][12] [8:0] }), .sum({ \level_5_sums[0][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[225] [4:0] }), .sum({ \level_1_sums[0][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[227] [4:0] }), .sum({ \level_1_sums[0][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[0][113] [5:0] }),
     .b({ \level_1_sums[0][112] [5:0] }), .sum({ \level_2_sums[0][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[229] [4:0] }), .sum({ \level_1_sums[0][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[231] [4:0] }), .sum({ \level_1_sums[0][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[0][115] [5:0] }),
     .b({ \level_1_sums[0][114] [5:0] }), .sum({ \level_2_sums[0][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[0][57] [6:0] }),
     .b({ \level_2_sums[0][56] [6:0] }), .sum({ \level_3_sums[0][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[233] [4:0] }), .sum({ \level_1_sums[0][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[235] [4:0] }), .sum({ \level_1_sums[0][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[0][117] [5:0] }),
     .b({ \level_1_sums[0][116] [5:0] }), .sum({ \level_2_sums[0][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[237] [4:0] }), .sum({ \level_1_sums[0][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[239] [4:0] }), .sum({ \level_1_sums[0][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[0][119] [5:0] }),
     .b({ \level_1_sums[0][118] [5:0] }), .sum({ \level_2_sums[0][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[0][59] [6:0] }),
     .b({ \level_2_sums[0][58] [6:0] }), .sum({ \level_3_sums[0][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[0][29] [7:0] }),
     .b({ \level_3_sums[0][28] [7:0] }), .sum({ \level_4_sums[0][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[241] [4:0] }), .sum({ \level_1_sums[0][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[243] [4:0] }), .sum({ \level_1_sums[0][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[0][121] [5:0] }),
     .b({ \level_1_sums[0][120] [5:0] }), .sum({ \level_2_sums[0][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[245] [4:0] }), .sum({ \level_1_sums[0][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[247] [4:0] }), .sum({ \level_1_sums[0][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[0][123] [5:0] }),
     .b({ \level_1_sums[0][122] [5:0] }), .sum({ \level_2_sums[0][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[0][61] [6:0] }),
     .b({ \level_2_sums[0][60] [6:0] }), .sum({ \level_3_sums[0][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[249] [4:0] }), .sum({ \level_1_sums[0][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[251] [4:0] }), .sum({ \level_1_sums[0][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[0][125] [5:0] }),
     .b({ \level_1_sums[0][124] [5:0] }), .sum({ \level_2_sums[0][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[253] [4:0] }), .sum({ \level_1_sums[0][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[0].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[0].product_terms[255] [4:0] }), .sum({ \level_1_sums[0][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[0][127] [5:0] }),
     .b({ \level_1_sums[0][126] [5:0] }), .sum({ \level_2_sums[0][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[0][63] [6:0] }),
     .b({ \level_2_sums[0][62] [6:0] }), .sum({ \level_3_sums[0][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[0][31] [7:0] }),
     .b({ \level_3_sums[0][30] [7:0] }), .sum({ \level_4_sums[0][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[0][15] [8:0] }),
     .b({ \level_4_sums[0][14] [8:0] }), .sum({ \level_5_sums[0][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[0][7] [9:0] }),
     .b({ \level_5_sums[0][6] [9:0] }), .sum({ \level_6_sums[0][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[0][3] [9:0] }),
     .b({ \level_6_sums[0][2] [9:0] }), .sum({ \level_7_sums[0][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[0].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[0][0] [9:0] }),
     .b({ \level_7_sums[0][1] [9:0] }), .sum({ \level_8_sums[0] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[1].relu_inst (.in_data({ \final_sums[1] [9:0] }), .out_data({ \out_sig[1] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[1] [4:0] }), .sum({ \level_1_sums[1][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[3] [4:0] }), .sum({ \level_1_sums[1][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[1][1] [5:0] }),
     .b({ \level_1_sums[1][0] [5:0] }), .sum({ \level_2_sums[1][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[5] [4:0] }), .sum({ \level_1_sums[1][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[7] [4:0] }), .sum({ \level_1_sums[1][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[1][3] [5:0] }),
     .b({ \level_1_sums[1][2] [5:0] }), .sum({ \level_2_sums[1][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[1][1] [6:0] }),
     .b({ \level_2_sums[1][0] [6:0] }), .sum({ \level_3_sums[1][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[9] [4:0] }), .sum({ \level_1_sums[1][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[11] [4:0] }), .sum({ \level_1_sums[1][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[1][5] [5:0] }),
     .b({ \level_1_sums[1][4] [5:0] }), .sum({ \level_2_sums[1][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[13] [4:0] }), .sum({ \level_1_sums[1][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[15] [4:0] }), .sum({ \level_1_sums[1][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[1][7] [5:0] }),
     .b({ \level_1_sums[1][6] [5:0] }), .sum({ \level_2_sums[1][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[1][3] [6:0] }),
     .b({ \level_2_sums[1][2] [6:0] }), .sum({ \level_3_sums[1][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[1][1] [7:0] }),
     .b({ \level_3_sums[1][0] [7:0] }), .sum({ \level_4_sums[1][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[17] [4:0] }), .sum({ \level_1_sums[1][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[19] [4:0] }), .sum({ \level_1_sums[1][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[1][9] [5:0] }),
     .b({ \level_1_sums[1][8] [5:0] }), .sum({ \level_2_sums[1][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[21] [4:0] }), .sum({ \level_1_sums[1][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[23] [4:0] }), .sum({ \level_1_sums[1][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[1][11] [5:0] }),
     .b({ \level_1_sums[1][10] [5:0] }), .sum({ \level_2_sums[1][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[1][5] [6:0] }),
     .b({ \level_2_sums[1][4] [6:0] }), .sum({ \level_3_sums[1][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[25] [4:0] }), .sum({ \level_1_sums[1][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[27] [4:0] }), .sum({ \level_1_sums[1][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[1][13] [5:0] }),
     .b({ \level_1_sums[1][12] [5:0] }), .sum({ \level_2_sums[1][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[29] [4:0] }), .sum({ \level_1_sums[1][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[31] [4:0] }), .sum({ \level_1_sums[1][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[1][15] [5:0] }),
     .b({ \level_1_sums[1][14] [5:0] }), .sum({ \level_2_sums[1][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[1][7] [6:0] }),
     .b({ \level_2_sums[1][6] [6:0] }), .sum({ \level_3_sums[1][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[1][3] [7:0] }),
     .b({ \level_3_sums[1][2] [7:0] }), .sum({ \level_4_sums[1][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[1][1] [8:0] }),
     .b({ \level_4_sums[1][0] [8:0] }), .sum({ \level_5_sums[1][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[33] [4:0] }), .sum({ \level_1_sums[1][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[35] [4:0] }), .sum({ \level_1_sums[1][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[1][17] [5:0] }),
     .b({ \level_1_sums[1][16] [5:0] }), .sum({ \level_2_sums[1][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[37] [4:0] }), .sum({ \level_1_sums[1][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[39] [4:0] }), .sum({ \level_1_sums[1][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[1][19] [5:0] }),
     .b({ \level_1_sums[1][18] [5:0] }), .sum({ \level_2_sums[1][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[1][9] [6:0] }),
     .b({ \level_2_sums[1][8] [6:0] }), .sum({ \level_3_sums[1][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[41] [4:0] }), .sum({ \level_1_sums[1][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[43] [4:0] }), .sum({ \level_1_sums[1][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[1][21] [5:0] }),
     .b({ \level_1_sums[1][20] [5:0] }), .sum({ \level_2_sums[1][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[45] [4:0] }), .sum({ \level_1_sums[1][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[47] [4:0] }), .sum({ \level_1_sums[1][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[1][23] [5:0] }),
     .b({ \level_1_sums[1][22] [5:0] }), .sum({ \level_2_sums[1][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[1][11] [6:0] }),
     .b({ \level_2_sums[1][10] [6:0] }), .sum({ \level_3_sums[1][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[1][5] [7:0] }),
     .b({ \level_3_sums[1][4] [7:0] }), .sum({ \level_4_sums[1][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[49] [4:0] }), .sum({ \level_1_sums[1][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[51] [4:0] }), .sum({ \level_1_sums[1][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[1][25] [5:0] }),
     .b({ \level_1_sums[1][24] [5:0] }), .sum({ \level_2_sums[1][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[53] [4:0] }), .sum({ \level_1_sums[1][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[55] [4:0] }), .sum({ \level_1_sums[1][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[1][27] [5:0] }),
     .b({ \level_1_sums[1][26] [5:0] }), .sum({ \level_2_sums[1][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[1][13] [6:0] }),
     .b({ \level_2_sums[1][12] [6:0] }), .sum({ \level_3_sums[1][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[57] [4:0] }), .sum({ \level_1_sums[1][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[59] [4:0] }), .sum({ \level_1_sums[1][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[1][29] [5:0] }),
     .b({ \level_1_sums[1][28] [5:0] }), .sum({ \level_2_sums[1][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[61] [4:0] }), .sum({ \level_1_sums[1][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[63] [4:0] }), .sum({ \level_1_sums[1][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[1][31] [5:0] }),
     .b({ \level_1_sums[1][30] [5:0] }), .sum({ \level_2_sums[1][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[1][15] [6:0] }),
     .b({ \level_2_sums[1][14] [6:0] }), .sum({ \level_3_sums[1][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[1][7] [7:0] }),
     .b({ \level_3_sums[1][6] [7:0] }), .sum({ \level_4_sums[1][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[1][3] [8:0] }),
     .b({ \level_4_sums[1][2] [8:0] }), .sum({ \level_5_sums[1][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[1][1] [9:0] }),
     .b({ \level_5_sums[1][0] [9:0] }), .sum({ \level_6_sums[1][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[65] [4:0] }), .sum({ \level_1_sums[1][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[67] [4:0] }), .sum({ \level_1_sums[1][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[1][33] [5:0] }),
     .b({ \level_1_sums[1][32] [5:0] }), .sum({ \level_2_sums[1][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[69] [4:0] }), .sum({ \level_1_sums[1][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[71] [4:0] }), .sum({ \level_1_sums[1][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[1][35] [5:0] }),
     .b({ \level_1_sums[1][34] [5:0] }), .sum({ \level_2_sums[1][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[1][17] [6:0] }),
     .b({ \level_2_sums[1][16] [6:0] }), .sum({ \level_3_sums[1][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[73] [4:0] }), .sum({ \level_1_sums[1][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[75] [4:0] }), .sum({ \level_1_sums[1][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[1][37] [5:0] }),
     .b({ \level_1_sums[1][36] [5:0] }), .sum({ \level_2_sums[1][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[77] [4:0] }), .sum({ \level_1_sums[1][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[79] [4:0] }), .sum({ \level_1_sums[1][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[1][39] [5:0] }),
     .b({ \level_1_sums[1][38] [5:0] }), .sum({ \level_2_sums[1][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[1][19] [6:0] }),
     .b({ \level_2_sums[1][18] [6:0] }), .sum({ \level_3_sums[1][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[1][9] [7:0] }),
     .b({ \level_3_sums[1][8] [7:0] }), .sum({ \level_4_sums[1][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[81] [4:0] }), .sum({ \level_1_sums[1][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[83] [4:0] }), .sum({ \level_1_sums[1][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[1][41] [5:0] }),
     .b({ \level_1_sums[1][40] [5:0] }), .sum({ \level_2_sums[1][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[85] [4:0] }), .sum({ \level_1_sums[1][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[87] [4:0] }), .sum({ \level_1_sums[1][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[1][43] [5:0] }),
     .b({ \level_1_sums[1][42] [5:0] }), .sum({ \level_2_sums[1][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[1][21] [6:0] }),
     .b({ \level_2_sums[1][20] [6:0] }), .sum({ \level_3_sums[1][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[89] [4:0] }), .sum({ \level_1_sums[1][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[91] [4:0] }), .sum({ \level_1_sums[1][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[1][45] [5:0] }),
     .b({ \level_1_sums[1][44] [5:0] }), .sum({ \level_2_sums[1][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[93] [4:0] }), .sum({ \level_1_sums[1][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[95] [4:0] }), .sum({ \level_1_sums[1][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[1][47] [5:0] }),
     .b({ \level_1_sums[1][46] [5:0] }), .sum({ \level_2_sums[1][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[1][23] [6:0] }),
     .b({ \level_2_sums[1][22] [6:0] }), .sum({ \level_3_sums[1][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[1][11] [7:0] }),
     .b({ \level_3_sums[1][10] [7:0] }), .sum({ \level_4_sums[1][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[1][5] [8:0] }),
     .b({ \level_4_sums[1][4] [8:0] }), .sum({ \level_5_sums[1][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[97] [4:0] }), .sum({ \level_1_sums[1][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[99] [4:0] }), .sum({ \level_1_sums[1][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[1][49] [5:0] }),
     .b({ \level_1_sums[1][48] [5:0] }), .sum({ \level_2_sums[1][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[101] [4:0] }), .sum({ \level_1_sums[1][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[103] [4:0] }), .sum({ \level_1_sums[1][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[1][51] [5:0] }),
     .b({ \level_1_sums[1][50] [5:0] }), .sum({ \level_2_sums[1][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[1][25] [6:0] }),
     .b({ \level_2_sums[1][24] [6:0] }), .sum({ \level_3_sums[1][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[105] [4:0] }), .sum({ \level_1_sums[1][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[107] [4:0] }), .sum({ \level_1_sums[1][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[1][53] [5:0] }),
     .b({ \level_1_sums[1][52] [5:0] }), .sum({ \level_2_sums[1][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[109] [4:0] }), .sum({ \level_1_sums[1][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[111] [4:0] }), .sum({ \level_1_sums[1][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[1][55] [5:0] }),
     .b({ \level_1_sums[1][54] [5:0] }), .sum({ \level_2_sums[1][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[1][27] [6:0] }),
     .b({ \level_2_sums[1][26] [6:0] }), .sum({ \level_3_sums[1][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[1][13] [7:0] }),
     .b({ \level_3_sums[1][12] [7:0] }), .sum({ \level_4_sums[1][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[113] [4:0] }), .sum({ \level_1_sums[1][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[115] [4:0] }), .sum({ \level_1_sums[1][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[1][57] [5:0] }),
     .b({ \level_1_sums[1][56] [5:0] }), .sum({ \level_2_sums[1][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[117] [4:0] }), .sum({ \level_1_sums[1][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[119] [4:0] }), .sum({ \level_1_sums[1][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[1][59] [5:0] }),
     .b({ \level_1_sums[1][58] [5:0] }), .sum({ \level_2_sums[1][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[1][29] [6:0] }),
     .b({ \level_2_sums[1][28] [6:0] }), .sum({ \level_3_sums[1][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[121] [4:0] }), .sum({ \level_1_sums[1][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[123] [4:0] }), .sum({ \level_1_sums[1][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[1][61] [5:0] }),
     .b({ \level_1_sums[1][60] [5:0] }), .sum({ \level_2_sums[1][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[125] [4:0] }), .sum({ \level_1_sums[1][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[127] [4:0] }), .sum({ \level_1_sums[1][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[1][63] [5:0] }),
     .b({ \level_1_sums[1][62] [5:0] }), .sum({ \level_2_sums[1][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[1][31] [6:0] }),
     .b({ \level_2_sums[1][30] [6:0] }), .sum({ \level_3_sums[1][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[1][15] [7:0] }),
     .b({ \level_3_sums[1][14] [7:0] }), .sum({ \level_4_sums[1][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[1][7] [8:0] }),
     .b({ \level_4_sums[1][6] [8:0] }), .sum({ \level_5_sums[1][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[1][3] [9:0] }),
     .b({ \level_5_sums[1][2] [9:0] }), .sum({ \level_6_sums[1][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[1][1] [9:0] }),
     .b({ \level_6_sums[1][0] [9:0] }), .sum({ \level_7_sums[1][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[129] [4:0] }), .sum({ \level_1_sums[1][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[131] [4:0] }), .sum({ \level_1_sums[1][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[1][65] [5:0] }),
     .b({ \level_1_sums[1][64] [5:0] }), .sum({ \level_2_sums[1][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[133] [4:0] }), .sum({ \level_1_sums[1][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[135] [4:0] }), .sum({ \level_1_sums[1][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[1][67] [5:0] }),
     .b({ \level_1_sums[1][66] [5:0] }), .sum({ \level_2_sums[1][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[1][33] [6:0] }),
     .b({ \level_2_sums[1][32] [6:0] }), .sum({ \level_3_sums[1][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[137] [4:0] }), .sum({ \level_1_sums[1][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[139] [4:0] }), .sum({ \level_1_sums[1][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[1][69] [5:0] }),
     .b({ \level_1_sums[1][68] [5:0] }), .sum({ \level_2_sums[1][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[141] [4:0] }), .sum({ \level_1_sums[1][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[143] [4:0] }), .sum({ \level_1_sums[1][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[1][71] [5:0] }),
     .b({ \level_1_sums[1][70] [5:0] }), .sum({ \level_2_sums[1][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[1][35] [6:0] }),
     .b({ \level_2_sums[1][34] [6:0] }), .sum({ \level_3_sums[1][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[1][17] [7:0] }),
     .b({ \level_3_sums[1][16] [7:0] }), .sum({ \level_4_sums[1][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[145] [4:0] }), .sum({ \level_1_sums[1][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[147] [4:0] }), .sum({ \level_1_sums[1][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[1][73] [5:0] }),
     .b({ \level_1_sums[1][72] [5:0] }), .sum({ \level_2_sums[1][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[149] [4:0] }), .sum({ \level_1_sums[1][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[151] [4:0] }), .sum({ \level_1_sums[1][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[1][75] [5:0] }),
     .b({ \level_1_sums[1][74] [5:0] }), .sum({ \level_2_sums[1][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[1][37] [6:0] }),
     .b({ \level_2_sums[1][36] [6:0] }), .sum({ \level_3_sums[1][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[153] [4:0] }), .sum({ \level_1_sums[1][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[155] [4:0] }), .sum({ \level_1_sums[1][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[1][77] [5:0] }),
     .b({ \level_1_sums[1][76] [5:0] }), .sum({ \level_2_sums[1][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[157] [4:0] }), .sum({ \level_1_sums[1][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[159] [4:0] }), .sum({ \level_1_sums[1][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[1][79] [5:0] }),
     .b({ \level_1_sums[1][78] [5:0] }), .sum({ \level_2_sums[1][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[1][39] [6:0] }),
     .b({ \level_2_sums[1][38] [6:0] }), .sum({ \level_3_sums[1][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[1][19] [7:0] }),
     .b({ \level_3_sums[1][18] [7:0] }), .sum({ \level_4_sums[1][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[1][9] [8:0] }),
     .b({ \level_4_sums[1][8] [8:0] }), .sum({ \level_5_sums[1][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[161] [4:0] }), .sum({ \level_1_sums[1][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[163] [4:0] }), .sum({ \level_1_sums[1][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[1][81] [5:0] }),
     .b({ \level_1_sums[1][80] [5:0] }), .sum({ \level_2_sums[1][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[165] [4:0] }), .sum({ \level_1_sums[1][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[167] [4:0] }), .sum({ \level_1_sums[1][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[1][83] [5:0] }),
     .b({ \level_1_sums[1][82] [5:0] }), .sum({ \level_2_sums[1][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[1][41] [6:0] }),
     .b({ \level_2_sums[1][40] [6:0] }), .sum({ \level_3_sums[1][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[169] [4:0] }), .sum({ \level_1_sums[1][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[171] [4:0] }), .sum({ \level_1_sums[1][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[1][85] [5:0] }),
     .b({ \level_1_sums[1][84] [5:0] }), .sum({ \level_2_sums[1][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[173] [4:0] }), .sum({ \level_1_sums[1][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[175] [4:0] }), .sum({ \level_1_sums[1][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[1][87] [5:0] }),
     .b({ \level_1_sums[1][86] [5:0] }), .sum({ \level_2_sums[1][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[1][43] [6:0] }),
     .b({ \level_2_sums[1][42] [6:0] }), .sum({ \level_3_sums[1][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[1][21] [7:0] }),
     .b({ \level_3_sums[1][20] [7:0] }), .sum({ \level_4_sums[1][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[177] [4:0] }), .sum({ \level_1_sums[1][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[179] [4:0] }), .sum({ \level_1_sums[1][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[1][89] [5:0] }),
     .b({ \level_1_sums[1][88] [5:0] }), .sum({ \level_2_sums[1][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[181] [4:0] }), .sum({ \level_1_sums[1][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[183] [4:0] }), .sum({ \level_1_sums[1][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[1][91] [5:0] }),
     .b({ \level_1_sums[1][90] [5:0] }), .sum({ \level_2_sums[1][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[1][45] [6:0] }),
     .b({ \level_2_sums[1][44] [6:0] }), .sum({ \level_3_sums[1][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[185] [4:0] }), .sum({ \level_1_sums[1][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[187] [4:0] }), .sum({ \level_1_sums[1][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[1][93] [5:0] }),
     .b({ \level_1_sums[1][92] [5:0] }), .sum({ \level_2_sums[1][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[189] [4:0] }), .sum({ \level_1_sums[1][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[191] [4:0] }), .sum({ \level_1_sums[1][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[1][95] [5:0] }),
     .b({ \level_1_sums[1][94] [5:0] }), .sum({ \level_2_sums[1][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[1][47] [6:0] }),
     .b({ \level_2_sums[1][46] [6:0] }), .sum({ \level_3_sums[1][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[1][23] [7:0] }),
     .b({ \level_3_sums[1][22] [7:0] }), .sum({ \level_4_sums[1][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[1][11] [8:0] }),
     .b({ \level_4_sums[1][10] [8:0] }), .sum({ \level_5_sums[1][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[1][5] [9:0] }),
     .b({ \level_5_sums[1][4] [9:0] }), .sum({ \level_6_sums[1][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[193] [4:0] }), .sum({ \level_1_sums[1][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[195] [4:0] }), .sum({ \level_1_sums[1][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[1][97] [5:0] }),
     .b({ \level_1_sums[1][96] [5:0] }), .sum({ \level_2_sums[1][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[197] [4:0] }), .sum({ \level_1_sums[1][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[199] [4:0] }), .sum({ \level_1_sums[1][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[1][99] [5:0] }),
     .b({ \level_1_sums[1][98] [5:0] }), .sum({ \level_2_sums[1][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[1][49] [6:0] }),
     .b({ \level_2_sums[1][48] [6:0] }), .sum({ \level_3_sums[1][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[201] [4:0] }), .sum({ \level_1_sums[1][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[203] [4:0] }), .sum({ \level_1_sums[1][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[1][101] [5:0] }),
     .b({ \level_1_sums[1][100] [5:0] }), .sum({ \level_2_sums[1][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[205] [4:0] }), .sum({ \level_1_sums[1][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[207] [4:0] }), .sum({ \level_1_sums[1][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[1][103] [5:0] }),
     .b({ \level_1_sums[1][102] [5:0] }), .sum({ \level_2_sums[1][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[1][51] [6:0] }),
     .b({ \level_2_sums[1][50] [6:0] }), .sum({ \level_3_sums[1][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[1][25] [7:0] }),
     .b({ \level_3_sums[1][24] [7:0] }), .sum({ \level_4_sums[1][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[209] [4:0] }), .sum({ \level_1_sums[1][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[211] [4:0] }), .sum({ \level_1_sums[1][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[1][105] [5:0] }),
     .b({ \level_1_sums[1][104] [5:0] }), .sum({ \level_2_sums[1][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[213] [4:0] }), .sum({ \level_1_sums[1][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[215] [4:0] }), .sum({ \level_1_sums[1][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[1][107] [5:0] }),
     .b({ \level_1_sums[1][106] [5:0] }), .sum({ \level_2_sums[1][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[1][53] [6:0] }),
     .b({ \level_2_sums[1][52] [6:0] }), .sum({ \level_3_sums[1][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[217] [4:0] }), .sum({ \level_1_sums[1][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[219] [4:0] }), .sum({ \level_1_sums[1][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[1][109] [5:0] }),
     .b({ \level_1_sums[1][108] [5:0] }), .sum({ \level_2_sums[1][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[221] [4:0] }), .sum({ \level_1_sums[1][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[223] [4:0] }), .sum({ \level_1_sums[1][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[1][111] [5:0] }),
     .b({ \level_1_sums[1][110] [5:0] }), .sum({ \level_2_sums[1][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[1][55] [6:0] }),
     .b({ \level_2_sums[1][54] [6:0] }), .sum({ \level_3_sums[1][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[1][27] [7:0] }),
     .b({ \level_3_sums[1][26] [7:0] }), .sum({ \level_4_sums[1][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[1][13] [8:0] }),
     .b({ \level_4_sums[1][12] [8:0] }), .sum({ \level_5_sums[1][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[225] [4:0] }), .sum({ \level_1_sums[1][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[227] [4:0] }), .sum({ \level_1_sums[1][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[1][113] [5:0] }),
     .b({ \level_1_sums[1][112] [5:0] }), .sum({ \level_2_sums[1][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[229] [4:0] }), .sum({ \level_1_sums[1][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[231] [4:0] }), .sum({ \level_1_sums[1][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[1][115] [5:0] }),
     .b({ \level_1_sums[1][114] [5:0] }), .sum({ \level_2_sums[1][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[1][57] [6:0] }),
     .b({ \level_2_sums[1][56] [6:0] }), .sum({ \level_3_sums[1][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[233] [4:0] }), .sum({ \level_1_sums[1][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[235] [4:0] }), .sum({ \level_1_sums[1][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[1][117] [5:0] }),
     .b({ \level_1_sums[1][116] [5:0] }), .sum({ \level_2_sums[1][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[237] [4:0] }), .sum({ \level_1_sums[1][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[239] [4:0] }), .sum({ \level_1_sums[1][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[1][119] [5:0] }),
     .b({ \level_1_sums[1][118] [5:0] }), .sum({ \level_2_sums[1][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[1][59] [6:0] }),
     .b({ \level_2_sums[1][58] [6:0] }), .sum({ \level_3_sums[1][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[1][29] [7:0] }),
     .b({ \level_3_sums[1][28] [7:0] }), .sum({ \level_4_sums[1][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[241] [4:0] }), .sum({ \level_1_sums[1][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[243] [4:0] }), .sum({ \level_1_sums[1][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[1][121] [5:0] }),
     .b({ \level_1_sums[1][120] [5:0] }), .sum({ \level_2_sums[1][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[245] [4:0] }), .sum({ \level_1_sums[1][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[247] [4:0] }), .sum({ \level_1_sums[1][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[1][123] [5:0] }),
     .b({ \level_1_sums[1][122] [5:0] }), .sum({ \level_2_sums[1][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[1][61] [6:0] }),
     .b({ \level_2_sums[1][60] [6:0] }), .sum({ \level_3_sums[1][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[249] [4:0] }), .sum({ \level_1_sums[1][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[251] [4:0] }), .sum({ \level_1_sums[1][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[1][125] [5:0] }),
     .b({ \level_1_sums[1][124] [5:0] }), .sum({ \level_2_sums[1][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[253] [4:0] }), .sum({ \level_1_sums[1][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[1].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[1].product_terms[255] [4:0] }), .sum({ \level_1_sums[1][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[1][127] [5:0] }),
     .b({ \level_1_sums[1][126] [5:0] }), .sum({ \level_2_sums[1][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[1][63] [6:0] }),
     .b({ \level_2_sums[1][62] [6:0] }), .sum({ \level_3_sums[1][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[1][31] [7:0] }),
     .b({ \level_3_sums[1][30] [7:0] }), .sum({ \level_4_sums[1][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[1][15] [8:0] }),
     .b({ \level_4_sums[1][14] [8:0] }), .sum({ \level_5_sums[1][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[1][7] [9:0] }),
     .b({ \level_5_sums[1][6] [9:0] }), .sum({ \level_6_sums[1][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[1][3] [9:0] }),
     .b({ \level_6_sums[1][2] [9:0] }), .sum({ \level_7_sums[1][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[1].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[1][0] [9:0] }),
     .b({ \level_7_sums[1][1] [9:0] }), .sum({ \level_8_sums[1] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[2].relu_inst (.in_data({ \final_sums[2] [9:0] }), .out_data({ \out_sig[2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[1] [4:0] }), .sum({ \level_1_sums[2][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[3] [4:0] }), .sum({ \level_1_sums[2][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[2][1] [5:0] }),
     .b({ \level_1_sums[2][0] [5:0] }), .sum({ \level_2_sums[2][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[5] [4:0] }), .sum({ \level_1_sums[2][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[7] [4:0] }), .sum({ \level_1_sums[2][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[2][3] [5:0] }),
     .b({ \level_1_sums[2][2] [5:0] }), .sum({ \level_2_sums[2][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[2][1] [6:0] }),
     .b({ \level_2_sums[2][0] [6:0] }), .sum({ \level_3_sums[2][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[9] [4:0] }), .sum({ \level_1_sums[2][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[11] [4:0] }), .sum({ \level_1_sums[2][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[2][5] [5:0] }),
     .b({ \level_1_sums[2][4] [5:0] }), .sum({ \level_2_sums[2][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[13] [4:0] }), .sum({ \level_1_sums[2][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[15] [4:0] }), .sum({ \level_1_sums[2][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[2][7] [5:0] }),
     .b({ \level_1_sums[2][6] [5:0] }), .sum({ \level_2_sums[2][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[2][3] [6:0] }),
     .b({ \level_2_sums[2][2] [6:0] }), .sum({ \level_3_sums[2][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[2][1] [7:0] }),
     .b({ \level_3_sums[2][0] [7:0] }), .sum({ \level_4_sums[2][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[17] [4:0] }), .sum({ \level_1_sums[2][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[19] [4:0] }), .sum({ \level_1_sums[2][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[2][9] [5:0] }),
     .b({ \level_1_sums[2][8] [5:0] }), .sum({ \level_2_sums[2][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[21] [4:0] }), .sum({ \level_1_sums[2][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[23] [4:0] }), .sum({ \level_1_sums[2][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[2][11] [5:0] }),
     .b({ \level_1_sums[2][10] [5:0] }), .sum({ \level_2_sums[2][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[2][5] [6:0] }),
     .b({ \level_2_sums[2][4] [6:0] }), .sum({ \level_3_sums[2][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[25] [4:0] }), .sum({ \level_1_sums[2][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[27] [4:0] }), .sum({ \level_1_sums[2][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[2][13] [5:0] }),
     .b({ \level_1_sums[2][12] [5:0] }), .sum({ \level_2_sums[2][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[29] [4:0] }), .sum({ \level_1_sums[2][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[31] [4:0] }), .sum({ \level_1_sums[2][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[2][15] [5:0] }),
     .b({ \level_1_sums[2][14] [5:0] }), .sum({ \level_2_sums[2][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[2][7] [6:0] }),
     .b({ \level_2_sums[2][6] [6:0] }), .sum({ \level_3_sums[2][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[2][3] [7:0] }),
     .b({ \level_3_sums[2][2] [7:0] }), .sum({ \level_4_sums[2][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[2][1] [8:0] }),
     .b({ \level_4_sums[2][0] [8:0] }), .sum({ \level_5_sums[2][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[33] [4:0] }), .sum({ \level_1_sums[2][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[35] [4:0] }), .sum({ \level_1_sums[2][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[2][17] [5:0] }),
     .b({ \level_1_sums[2][16] [5:0] }), .sum({ \level_2_sums[2][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[37] [4:0] }), .sum({ \level_1_sums[2][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[39] [4:0] }), .sum({ \level_1_sums[2][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[2][19] [5:0] }),
     .b({ \level_1_sums[2][18] [5:0] }), .sum({ \level_2_sums[2][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[2][9] [6:0] }),
     .b({ \level_2_sums[2][8] [6:0] }), .sum({ \level_3_sums[2][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[41] [4:0] }), .sum({ \level_1_sums[2][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[43] [4:0] }), .sum({ \level_1_sums[2][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[2][21] [5:0] }),
     .b({ \level_1_sums[2][20] [5:0] }), .sum({ \level_2_sums[2][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[45] [4:0] }), .sum({ \level_1_sums[2][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[47] [4:0] }), .sum({ \level_1_sums[2][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[2][23] [5:0] }),
     .b({ \level_1_sums[2][22] [5:0] }), .sum({ \level_2_sums[2][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[2][11] [6:0] }),
     .b({ \level_2_sums[2][10] [6:0] }), .sum({ \level_3_sums[2][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[2][5] [7:0] }),
     .b({ \level_3_sums[2][4] [7:0] }), .sum({ \level_4_sums[2][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[49] [4:0] }), .sum({ \level_1_sums[2][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[51] [4:0] }), .sum({ \level_1_sums[2][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[2][25] [5:0] }),
     .b({ \level_1_sums[2][24] [5:0] }), .sum({ \level_2_sums[2][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[53] [4:0] }), .sum({ \level_1_sums[2][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[55] [4:0] }), .sum({ \level_1_sums[2][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[2][27] [5:0] }),
     .b({ \level_1_sums[2][26] [5:0] }), .sum({ \level_2_sums[2][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[2][13] [6:0] }),
     .b({ \level_2_sums[2][12] [6:0] }), .sum({ \level_3_sums[2][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[57] [4:0] }), .sum({ \level_1_sums[2][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[59] [4:0] }), .sum({ \level_1_sums[2][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[2][29] [5:0] }),
     .b({ \level_1_sums[2][28] [5:0] }), .sum({ \level_2_sums[2][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[61] [4:0] }), .sum({ \level_1_sums[2][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[63] [4:0] }), .sum({ \level_1_sums[2][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[2][31] [5:0] }),
     .b({ \level_1_sums[2][30] [5:0] }), .sum({ \level_2_sums[2][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[2][15] [6:0] }),
     .b({ \level_2_sums[2][14] [6:0] }), .sum({ \level_3_sums[2][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[2][7] [7:0] }),
     .b({ \level_3_sums[2][6] [7:0] }), .sum({ \level_4_sums[2][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[2][3] [8:0] }),
     .b({ \level_4_sums[2][2] [8:0] }), .sum({ \level_5_sums[2][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[2][1] [9:0] }),
     .b({ \level_5_sums[2][0] [9:0] }), .sum({ \level_6_sums[2][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[65] [4:0] }), .sum({ \level_1_sums[2][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[67] [4:0] }), .sum({ \level_1_sums[2][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[2][33] [5:0] }),
     .b({ \level_1_sums[2][32] [5:0] }), .sum({ \level_2_sums[2][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[69] [4:0] }), .sum({ \level_1_sums[2][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[71] [4:0] }), .sum({ \level_1_sums[2][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[2][35] [5:0] }),
     .b({ \level_1_sums[2][34] [5:0] }), .sum({ \level_2_sums[2][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[2][17] [6:0] }),
     .b({ \level_2_sums[2][16] [6:0] }), .sum({ \level_3_sums[2][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[73] [4:0] }), .sum({ \level_1_sums[2][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[75] [4:0] }), .sum({ \level_1_sums[2][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[2][37] [5:0] }),
     .b({ \level_1_sums[2][36] [5:0] }), .sum({ \level_2_sums[2][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[77] [4:0] }), .sum({ \level_1_sums[2][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[79] [4:0] }), .sum({ \level_1_sums[2][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[2][39] [5:0] }),
     .b({ \level_1_sums[2][38] [5:0] }), .sum({ \level_2_sums[2][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[2][19] [6:0] }),
     .b({ \level_2_sums[2][18] [6:0] }), .sum({ \level_3_sums[2][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[2][9] [7:0] }),
     .b({ \level_3_sums[2][8] [7:0] }), .sum({ \level_4_sums[2][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[81] [4:0] }), .sum({ \level_1_sums[2][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[83] [4:0] }), .sum({ \level_1_sums[2][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[2][41] [5:0] }),
     .b({ \level_1_sums[2][40] [5:0] }), .sum({ \level_2_sums[2][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[85] [4:0] }), .sum({ \level_1_sums[2][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[87] [4:0] }), .sum({ \level_1_sums[2][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[2][43] [5:0] }),
     .b({ \level_1_sums[2][42] [5:0] }), .sum({ \level_2_sums[2][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[2][21] [6:0] }),
     .b({ \level_2_sums[2][20] [6:0] }), .sum({ \level_3_sums[2][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[89] [4:0] }), .sum({ \level_1_sums[2][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[91] [4:0] }), .sum({ \level_1_sums[2][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[2][45] [5:0] }),
     .b({ \level_1_sums[2][44] [5:0] }), .sum({ \level_2_sums[2][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[93] [4:0] }), .sum({ \level_1_sums[2][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[95] [4:0] }), .sum({ \level_1_sums[2][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[2][47] [5:0] }),
     .b({ \level_1_sums[2][46] [5:0] }), .sum({ \level_2_sums[2][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[2][23] [6:0] }),
     .b({ \level_2_sums[2][22] [6:0] }), .sum({ \level_3_sums[2][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[2][11] [7:0] }),
     .b({ \level_3_sums[2][10] [7:0] }), .sum({ \level_4_sums[2][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[2][5] [8:0] }),
     .b({ \level_4_sums[2][4] [8:0] }), .sum({ \level_5_sums[2][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[97] [4:0] }), .sum({ \level_1_sums[2][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[99] [4:0] }), .sum({ \level_1_sums[2][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[2][49] [5:0] }),
     .b({ \level_1_sums[2][48] [5:0] }), .sum({ \level_2_sums[2][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[101] [4:0] }), .sum({ \level_1_sums[2][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[103] [4:0] }), .sum({ \level_1_sums[2][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[2][51] [5:0] }),
     .b({ \level_1_sums[2][50] [5:0] }), .sum({ \level_2_sums[2][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[2][25] [6:0] }),
     .b({ \level_2_sums[2][24] [6:0] }), .sum({ \level_3_sums[2][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[105] [4:0] }), .sum({ \level_1_sums[2][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[107] [4:0] }), .sum({ \level_1_sums[2][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[2][53] [5:0] }),
     .b({ \level_1_sums[2][52] [5:0] }), .sum({ \level_2_sums[2][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[109] [4:0] }), .sum({ \level_1_sums[2][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[111] [4:0] }), .sum({ \level_1_sums[2][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[2][55] [5:0] }),
     .b({ \level_1_sums[2][54] [5:0] }), .sum({ \level_2_sums[2][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[2][27] [6:0] }),
     .b({ \level_2_sums[2][26] [6:0] }), .sum({ \level_3_sums[2][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[2][13] [7:0] }),
     .b({ \level_3_sums[2][12] [7:0] }), .sum({ \level_4_sums[2][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[113] [4:0] }), .sum({ \level_1_sums[2][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[115] [4:0] }), .sum({ \level_1_sums[2][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[2][57] [5:0] }),
     .b({ \level_1_sums[2][56] [5:0] }), .sum({ \level_2_sums[2][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[117] [4:0] }), .sum({ \level_1_sums[2][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[119] [4:0] }), .sum({ \level_1_sums[2][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[2][59] [5:0] }),
     .b({ \level_1_sums[2][58] [5:0] }), .sum({ \level_2_sums[2][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[2][29] [6:0] }),
     .b({ \level_2_sums[2][28] [6:0] }), .sum({ \level_3_sums[2][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[121] [4:0] }), .sum({ \level_1_sums[2][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[123] [4:0] }), .sum({ \level_1_sums[2][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[2][61] [5:0] }),
     .b({ \level_1_sums[2][60] [5:0] }), .sum({ \level_2_sums[2][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[125] [4:0] }), .sum({ \level_1_sums[2][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[127] [4:0] }), .sum({ \level_1_sums[2][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[2][63] [5:0] }),
     .b({ \level_1_sums[2][62] [5:0] }), .sum({ \level_2_sums[2][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[2][31] [6:0] }),
     .b({ \level_2_sums[2][30] [6:0] }), .sum({ \level_3_sums[2][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[2][15] [7:0] }),
     .b({ \level_3_sums[2][14] [7:0] }), .sum({ \level_4_sums[2][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[2][7] [8:0] }),
     .b({ \level_4_sums[2][6] [8:0] }), .sum({ \level_5_sums[2][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[2][3] [9:0] }),
     .b({ \level_5_sums[2][2] [9:0] }), .sum({ \level_6_sums[2][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[2][1] [9:0] }),
     .b({ \level_6_sums[2][0] [9:0] }), .sum({ \level_7_sums[2][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[129] [4:0] }), .sum({ \level_1_sums[2][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[131] [4:0] }), .sum({ \level_1_sums[2][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[2][65] [5:0] }),
     .b({ \level_1_sums[2][64] [5:0] }), .sum({ \level_2_sums[2][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[133] [4:0] }), .sum({ \level_1_sums[2][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[135] [4:0] }), .sum({ \level_1_sums[2][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[2][67] [5:0] }),
     .b({ \level_1_sums[2][66] [5:0] }), .sum({ \level_2_sums[2][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[2][33] [6:0] }),
     .b({ \level_2_sums[2][32] [6:0] }), .sum({ \level_3_sums[2][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[137] [4:0] }), .sum({ \level_1_sums[2][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[139] [4:0] }), .sum({ \level_1_sums[2][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[2][69] [5:0] }),
     .b({ \level_1_sums[2][68] [5:0] }), .sum({ \level_2_sums[2][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[141] [4:0] }), .sum({ \level_1_sums[2][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[143] [4:0] }), .sum({ \level_1_sums[2][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[2][71] [5:0] }),
     .b({ \level_1_sums[2][70] [5:0] }), .sum({ \level_2_sums[2][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[2][35] [6:0] }),
     .b({ \level_2_sums[2][34] [6:0] }), .sum({ \level_3_sums[2][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[2][17] [7:0] }),
     .b({ \level_3_sums[2][16] [7:0] }), .sum({ \level_4_sums[2][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[145] [4:0] }), .sum({ \level_1_sums[2][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[147] [4:0] }), .sum({ \level_1_sums[2][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[2][73] [5:0] }),
     .b({ \level_1_sums[2][72] [5:0] }), .sum({ \level_2_sums[2][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[149] [4:0] }), .sum({ \level_1_sums[2][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[151] [4:0] }), .sum({ \level_1_sums[2][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[2][75] [5:0] }),
     .b({ \level_1_sums[2][74] [5:0] }), .sum({ \level_2_sums[2][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[2][37] [6:0] }),
     .b({ \level_2_sums[2][36] [6:0] }), .sum({ \level_3_sums[2][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[153] [4:0] }), .sum({ \level_1_sums[2][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[155] [4:0] }), .sum({ \level_1_sums[2][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[2][77] [5:0] }),
     .b({ \level_1_sums[2][76] [5:0] }), .sum({ \level_2_sums[2][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[157] [4:0] }), .sum({ \level_1_sums[2][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[159] [4:0] }), .sum({ \level_1_sums[2][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[2][79] [5:0] }),
     .b({ \level_1_sums[2][78] [5:0] }), .sum({ \level_2_sums[2][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[2][39] [6:0] }),
     .b({ \level_2_sums[2][38] [6:0] }), .sum({ \level_3_sums[2][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[2][19] [7:0] }),
     .b({ \level_3_sums[2][18] [7:0] }), .sum({ \level_4_sums[2][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[2][9] [8:0] }),
     .b({ \level_4_sums[2][8] [8:0] }), .sum({ \level_5_sums[2][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[161] [4:0] }), .sum({ \level_1_sums[2][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[163] [4:0] }), .sum({ \level_1_sums[2][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[2][81] [5:0] }),
     .b({ \level_1_sums[2][80] [5:0] }), .sum({ \level_2_sums[2][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[165] [4:0] }), .sum({ \level_1_sums[2][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[167] [4:0] }), .sum({ \level_1_sums[2][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[2][83] [5:0] }),
     .b({ \level_1_sums[2][82] [5:0] }), .sum({ \level_2_sums[2][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[2][41] [6:0] }),
     .b({ \level_2_sums[2][40] [6:0] }), .sum({ \level_3_sums[2][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[169] [4:0] }), .sum({ \level_1_sums[2][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[171] [4:0] }), .sum({ \level_1_sums[2][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[2][85] [5:0] }),
     .b({ \level_1_sums[2][84] [5:0] }), .sum({ \level_2_sums[2][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[173] [4:0] }), .sum({ \level_1_sums[2][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[175] [4:0] }), .sum({ \level_1_sums[2][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[2][87] [5:0] }),
     .b({ \level_1_sums[2][86] [5:0] }), .sum({ \level_2_sums[2][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[2][43] [6:0] }),
     .b({ \level_2_sums[2][42] [6:0] }), .sum({ \level_3_sums[2][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[2][21] [7:0] }),
     .b({ \level_3_sums[2][20] [7:0] }), .sum({ \level_4_sums[2][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[177] [4:0] }), .sum({ \level_1_sums[2][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[179] [4:0] }), .sum({ \level_1_sums[2][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[2][89] [5:0] }),
     .b({ \level_1_sums[2][88] [5:0] }), .sum({ \level_2_sums[2][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[181] [4:0] }), .sum({ \level_1_sums[2][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[183] [4:0] }), .sum({ \level_1_sums[2][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[2][91] [5:0] }),
     .b({ \level_1_sums[2][90] [5:0] }), .sum({ \level_2_sums[2][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[2][45] [6:0] }),
     .b({ \level_2_sums[2][44] [6:0] }), .sum({ \level_3_sums[2][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[185] [4:0] }), .sum({ \level_1_sums[2][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[187] [4:0] }), .sum({ \level_1_sums[2][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[2][93] [5:0] }),
     .b({ \level_1_sums[2][92] [5:0] }), .sum({ \level_2_sums[2][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[189] [4:0] }), .sum({ \level_1_sums[2][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[191] [4:0] }), .sum({ \level_1_sums[2][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[2][95] [5:0] }),
     .b({ \level_1_sums[2][94] [5:0] }), .sum({ \level_2_sums[2][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[2][47] [6:0] }),
     .b({ \level_2_sums[2][46] [6:0] }), .sum({ \level_3_sums[2][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[2][23] [7:0] }),
     .b({ \level_3_sums[2][22] [7:0] }), .sum({ \level_4_sums[2][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[2][11] [8:0] }),
     .b({ \level_4_sums[2][10] [8:0] }), .sum({ \level_5_sums[2][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[2][5] [9:0] }),
     .b({ \level_5_sums[2][4] [9:0] }), .sum({ \level_6_sums[2][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[193] [4:0] }), .sum({ \level_1_sums[2][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[195] [4:0] }), .sum({ \level_1_sums[2][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[2][97] [5:0] }),
     .b({ \level_1_sums[2][96] [5:0] }), .sum({ \level_2_sums[2][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[197] [4:0] }), .sum({ \level_1_sums[2][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[199] [4:0] }), .sum({ \level_1_sums[2][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[2][99] [5:0] }),
     .b({ \level_1_sums[2][98] [5:0] }), .sum({ \level_2_sums[2][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[2][49] [6:0] }),
     .b({ \level_2_sums[2][48] [6:0] }), .sum({ \level_3_sums[2][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[201] [4:0] }), .sum({ \level_1_sums[2][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[203] [4:0] }), .sum({ \level_1_sums[2][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[2][101] [5:0] }),
     .b({ \level_1_sums[2][100] [5:0] }), .sum({ \level_2_sums[2][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[205] [4:0] }), .sum({ \level_1_sums[2][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[207] [4:0] }), .sum({ \level_1_sums[2][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[2][103] [5:0] }),
     .b({ \level_1_sums[2][102] [5:0] }), .sum({ \level_2_sums[2][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[2][51] [6:0] }),
     .b({ \level_2_sums[2][50] [6:0] }), .sum({ \level_3_sums[2][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[2][25] [7:0] }),
     .b({ \level_3_sums[2][24] [7:0] }), .sum({ \level_4_sums[2][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[209] [4:0] }), .sum({ \level_1_sums[2][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[211] [4:0] }), .sum({ \level_1_sums[2][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[2][105] [5:0] }),
     .b({ \level_1_sums[2][104] [5:0] }), .sum({ \level_2_sums[2][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[213] [4:0] }), .sum({ \level_1_sums[2][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[215] [4:0] }), .sum({ \level_1_sums[2][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[2][107] [5:0] }),
     .b({ \level_1_sums[2][106] [5:0] }), .sum({ \level_2_sums[2][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[2][53] [6:0] }),
     .b({ \level_2_sums[2][52] [6:0] }), .sum({ \level_3_sums[2][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[217] [4:0] }), .sum({ \level_1_sums[2][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[219] [4:0] }), .sum({ \level_1_sums[2][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[2][109] [5:0] }),
     .b({ \level_1_sums[2][108] [5:0] }), .sum({ \level_2_sums[2][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[221] [4:0] }), .sum({ \level_1_sums[2][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[223] [4:0] }), .sum({ \level_1_sums[2][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[2][111] [5:0] }),
     .b({ \level_1_sums[2][110] [5:0] }), .sum({ \level_2_sums[2][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[2][55] [6:0] }),
     .b({ \level_2_sums[2][54] [6:0] }), .sum({ \level_3_sums[2][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[2][27] [7:0] }),
     .b({ \level_3_sums[2][26] [7:0] }), .sum({ \level_4_sums[2][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[2][13] [8:0] }),
     .b({ \level_4_sums[2][12] [8:0] }), .sum({ \level_5_sums[2][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[225] [4:0] }), .sum({ \level_1_sums[2][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[227] [4:0] }), .sum({ \level_1_sums[2][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[2][113] [5:0] }),
     .b({ \level_1_sums[2][112] [5:0] }), .sum({ \level_2_sums[2][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[229] [4:0] }), .sum({ \level_1_sums[2][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[231] [4:0] }), .sum({ \level_1_sums[2][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[2][115] [5:0] }),
     .b({ \level_1_sums[2][114] [5:0] }), .sum({ \level_2_sums[2][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[2][57] [6:0] }),
     .b({ \level_2_sums[2][56] [6:0] }), .sum({ \level_3_sums[2][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[233] [4:0] }), .sum({ \level_1_sums[2][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[235] [4:0] }), .sum({ \level_1_sums[2][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[2][117] [5:0] }),
     .b({ \level_1_sums[2][116] [5:0] }), .sum({ \level_2_sums[2][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[237] [4:0] }), .sum({ \level_1_sums[2][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[239] [4:0] }), .sum({ \level_1_sums[2][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[2][119] [5:0] }),
     .b({ \level_1_sums[2][118] [5:0] }), .sum({ \level_2_sums[2][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[2][59] [6:0] }),
     .b({ \level_2_sums[2][58] [6:0] }), .sum({ \level_3_sums[2][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[2][29] [7:0] }),
     .b({ \level_3_sums[2][28] [7:0] }), .sum({ \level_4_sums[2][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[241] [4:0] }), .sum({ \level_1_sums[2][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[243] [4:0] }), .sum({ \level_1_sums[2][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[2][121] [5:0] }),
     .b({ \level_1_sums[2][120] [5:0] }), .sum({ \level_2_sums[2][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[245] [4:0] }), .sum({ \level_1_sums[2][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[247] [4:0] }), .sum({ \level_1_sums[2][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[2][123] [5:0] }),
     .b({ \level_1_sums[2][122] [5:0] }), .sum({ \level_2_sums[2][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[2][61] [6:0] }),
     .b({ \level_2_sums[2][60] [6:0] }), .sum({ \level_3_sums[2][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[249] [4:0] }), .sum({ \level_1_sums[2][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[251] [4:0] }), .sum({ \level_1_sums[2][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[2][125] [5:0] }),
     .b({ \level_1_sums[2][124] [5:0] }), .sum({ \level_2_sums[2][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[253] [4:0] }), .sum({ \level_1_sums[2][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[2].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[2].product_terms[255] [4:0] }), .sum({ \level_1_sums[2][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[2][127] [5:0] }),
     .b({ \level_1_sums[2][126] [5:0] }), .sum({ \level_2_sums[2][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[2][63] [6:0] }),
     .b({ \level_2_sums[2][62] [6:0] }), .sum({ \level_3_sums[2][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[2][31] [7:0] }),
     .b({ \level_3_sums[2][30] [7:0] }), .sum({ \level_4_sums[2][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[2][15] [8:0] }),
     .b({ \level_4_sums[2][14] [8:0] }), .sum({ \level_5_sums[2][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[2][7] [9:0] }),
     .b({ \level_5_sums[2][6] [9:0] }), .sum({ \level_6_sums[2][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[2][3] [9:0] }),
     .b({ \level_6_sums[2][2] [9:0] }), .sum({ \level_7_sums[2][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[2].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[2][0] [9:0] }),
     .b({ \level_7_sums[2][1] [9:0] }), .sum({ \level_8_sums[2] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[3].relu_inst (.in_data({ \final_sums[3] [9:0] }), .out_data({ \out_sig[3] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[1] [4:0] }), .sum({ \level_1_sums[3][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[3] [4:0] }), .sum({ \level_1_sums[3][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[3][1] [5:0] }),
     .b({ \level_1_sums[3][0] [5:0] }), .sum({ \level_2_sums[3][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[5] [4:0] }), .sum({ \level_1_sums[3][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[7] [4:0] }), .sum({ \level_1_sums[3][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[3][3] [5:0] }),
     .b({ \level_1_sums[3][2] [5:0] }), .sum({ \level_2_sums[3][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[3][1] [6:0] }),
     .b({ \level_2_sums[3][0] [6:0] }), .sum({ \level_3_sums[3][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[9] [4:0] }), .sum({ \level_1_sums[3][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[11] [4:0] }), .sum({ \level_1_sums[3][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[3][5] [5:0] }),
     .b({ \level_1_sums[3][4] [5:0] }), .sum({ \level_2_sums[3][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[13] [4:0] }), .sum({ \level_1_sums[3][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[15] [4:0] }), .sum({ \level_1_sums[3][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[3][7] [5:0] }),
     .b({ \level_1_sums[3][6] [5:0] }), .sum({ \level_2_sums[3][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[3][3] [6:0] }),
     .b({ \level_2_sums[3][2] [6:0] }), .sum({ \level_3_sums[3][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[3][1] [7:0] }),
     .b({ \level_3_sums[3][0] [7:0] }), .sum({ \level_4_sums[3][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[17] [4:0] }), .sum({ \level_1_sums[3][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[19] [4:0] }), .sum({ \level_1_sums[3][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[3][9] [5:0] }),
     .b({ \level_1_sums[3][8] [5:0] }), .sum({ \level_2_sums[3][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[21] [4:0] }), .sum({ \level_1_sums[3][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[23] [4:0] }), .sum({ \level_1_sums[3][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[3][11] [5:0] }),
     .b({ \level_1_sums[3][10] [5:0] }), .sum({ \level_2_sums[3][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[3][5] [6:0] }),
     .b({ \level_2_sums[3][4] [6:0] }), .sum({ \level_3_sums[3][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[25] [4:0] }), .sum({ \level_1_sums[3][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[27] [4:0] }), .sum({ \level_1_sums[3][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[3][13] [5:0] }),
     .b({ \level_1_sums[3][12] [5:0] }), .sum({ \level_2_sums[3][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[29] [4:0] }), .sum({ \level_1_sums[3][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[31] [4:0] }), .sum({ \level_1_sums[3][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[3][15] [5:0] }),
     .b({ \level_1_sums[3][14] [5:0] }), .sum({ \level_2_sums[3][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[3][7] [6:0] }),
     .b({ \level_2_sums[3][6] [6:0] }), .sum({ \level_3_sums[3][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[3][3] [7:0] }),
     .b({ \level_3_sums[3][2] [7:0] }), .sum({ \level_4_sums[3][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[3][1] [8:0] }),
     .b({ \level_4_sums[3][0] [8:0] }), .sum({ \level_5_sums[3][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[33] [4:0] }), .sum({ \level_1_sums[3][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[35] [4:0] }), .sum({ \level_1_sums[3][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[3][17] [5:0] }),
     .b({ \level_1_sums[3][16] [5:0] }), .sum({ \level_2_sums[3][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[37] [4:0] }), .sum({ \level_1_sums[3][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[39] [4:0] }), .sum({ \level_1_sums[3][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[3][19] [5:0] }),
     .b({ \level_1_sums[3][18] [5:0] }), .sum({ \level_2_sums[3][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[3][9] [6:0] }),
     .b({ \level_2_sums[3][8] [6:0] }), .sum({ \level_3_sums[3][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[41] [4:0] }), .sum({ \level_1_sums[3][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[43] [4:0] }), .sum({ \level_1_sums[3][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[3][21] [5:0] }),
     .b({ \level_1_sums[3][20] [5:0] }), .sum({ \level_2_sums[3][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[45] [4:0] }), .sum({ \level_1_sums[3][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[47] [4:0] }), .sum({ \level_1_sums[3][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[3][23] [5:0] }),
     .b({ \level_1_sums[3][22] [5:0] }), .sum({ \level_2_sums[3][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[3][11] [6:0] }),
     .b({ \level_2_sums[3][10] [6:0] }), .sum({ \level_3_sums[3][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[3][5] [7:0] }),
     .b({ \level_3_sums[3][4] [7:0] }), .sum({ \level_4_sums[3][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[49] [4:0] }), .sum({ \level_1_sums[3][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[51] [4:0] }), .sum({ \level_1_sums[3][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[3][25] [5:0] }),
     .b({ \level_1_sums[3][24] [5:0] }), .sum({ \level_2_sums[3][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[53] [4:0] }), .sum({ \level_1_sums[3][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[55] [4:0] }), .sum({ \level_1_sums[3][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[3][27] [5:0] }),
     .b({ \level_1_sums[3][26] [5:0] }), .sum({ \level_2_sums[3][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[3][13] [6:0] }),
     .b({ \level_2_sums[3][12] [6:0] }), .sum({ \level_3_sums[3][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[57] [4:0] }), .sum({ \level_1_sums[3][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[59] [4:0] }), .sum({ \level_1_sums[3][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[3][29] [5:0] }),
     .b({ \level_1_sums[3][28] [5:0] }), .sum({ \level_2_sums[3][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[61] [4:0] }), .sum({ \level_1_sums[3][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[63] [4:0] }), .sum({ \level_1_sums[3][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[3][31] [5:0] }),
     .b({ \level_1_sums[3][30] [5:0] }), .sum({ \level_2_sums[3][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[3][15] [6:0] }),
     .b({ \level_2_sums[3][14] [6:0] }), .sum({ \level_3_sums[3][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[3][7] [7:0] }),
     .b({ \level_3_sums[3][6] [7:0] }), .sum({ \level_4_sums[3][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[3][3] [8:0] }),
     .b({ \level_4_sums[3][2] [8:0] }), .sum({ \level_5_sums[3][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[3][1] [9:0] }),
     .b({ \level_5_sums[3][0] [9:0] }), .sum({ \level_6_sums[3][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[65] [4:0] }), .sum({ \level_1_sums[3][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[67] [4:0] }), .sum({ \level_1_sums[3][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[3][33] [5:0] }),
     .b({ \level_1_sums[3][32] [5:0] }), .sum({ \level_2_sums[3][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[69] [4:0] }), .sum({ \level_1_sums[3][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[71] [4:0] }), .sum({ \level_1_sums[3][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[3][35] [5:0] }),
     .b({ \level_1_sums[3][34] [5:0] }), .sum({ \level_2_sums[3][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[3][17] [6:0] }),
     .b({ \level_2_sums[3][16] [6:0] }), .sum({ \level_3_sums[3][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[73] [4:0] }), .sum({ \level_1_sums[3][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[75] [4:0] }), .sum({ \level_1_sums[3][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[3][37] [5:0] }),
     .b({ \level_1_sums[3][36] [5:0] }), .sum({ \level_2_sums[3][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[77] [4:0] }), .sum({ \level_1_sums[3][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[79] [4:0] }), .sum({ \level_1_sums[3][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[3][39] [5:0] }),
     .b({ \level_1_sums[3][38] [5:0] }), .sum({ \level_2_sums[3][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[3][19] [6:0] }),
     .b({ \level_2_sums[3][18] [6:0] }), .sum({ \level_3_sums[3][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[3][9] [7:0] }),
     .b({ \level_3_sums[3][8] [7:0] }), .sum({ \level_4_sums[3][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[81] [4:0] }), .sum({ \level_1_sums[3][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[83] [4:0] }), .sum({ \level_1_sums[3][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[3][41] [5:0] }),
     .b({ \level_1_sums[3][40] [5:0] }), .sum({ \level_2_sums[3][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[85] [4:0] }), .sum({ \level_1_sums[3][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[87] [4:0] }), .sum({ \level_1_sums[3][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[3][43] [5:0] }),
     .b({ \level_1_sums[3][42] [5:0] }), .sum({ \level_2_sums[3][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[3][21] [6:0] }),
     .b({ \level_2_sums[3][20] [6:0] }), .sum({ \level_3_sums[3][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[89] [4:0] }), .sum({ \level_1_sums[3][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[91] [4:0] }), .sum({ \level_1_sums[3][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[3][45] [5:0] }),
     .b({ \level_1_sums[3][44] [5:0] }), .sum({ \level_2_sums[3][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[93] [4:0] }), .sum({ \level_1_sums[3][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[95] [4:0] }), .sum({ \level_1_sums[3][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[3][47] [5:0] }),
     .b({ \level_1_sums[3][46] [5:0] }), .sum({ \level_2_sums[3][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[3][23] [6:0] }),
     .b({ \level_2_sums[3][22] [6:0] }), .sum({ \level_3_sums[3][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[3][11] [7:0] }),
     .b({ \level_3_sums[3][10] [7:0] }), .sum({ \level_4_sums[3][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[3][5] [8:0] }),
     .b({ \level_4_sums[3][4] [8:0] }), .sum({ \level_5_sums[3][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[97] [4:0] }), .sum({ \level_1_sums[3][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[99] [4:0] }), .sum({ \level_1_sums[3][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[3][49] [5:0] }),
     .b({ \level_1_sums[3][48] [5:0] }), .sum({ \level_2_sums[3][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[101] [4:0] }), .sum({ \level_1_sums[3][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[103] [4:0] }), .sum({ \level_1_sums[3][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[3][51] [5:0] }),
     .b({ \level_1_sums[3][50] [5:0] }), .sum({ \level_2_sums[3][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[3][25] [6:0] }),
     .b({ \level_2_sums[3][24] [6:0] }), .sum({ \level_3_sums[3][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[105] [4:0] }), .sum({ \level_1_sums[3][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[107] [4:0] }), .sum({ \level_1_sums[3][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[3][53] [5:0] }),
     .b({ \level_1_sums[3][52] [5:0] }), .sum({ \level_2_sums[3][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[109] [4:0] }), .sum({ \level_1_sums[3][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[111] [4:0] }), .sum({ \level_1_sums[3][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[3][55] [5:0] }),
     .b({ \level_1_sums[3][54] [5:0] }), .sum({ \level_2_sums[3][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[3][27] [6:0] }),
     .b({ \level_2_sums[3][26] [6:0] }), .sum({ \level_3_sums[3][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[3][13] [7:0] }),
     .b({ \level_3_sums[3][12] [7:0] }), .sum({ \level_4_sums[3][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[113] [4:0] }), .sum({ \level_1_sums[3][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[115] [4:0] }), .sum({ \level_1_sums[3][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[3][57] [5:0] }),
     .b({ \level_1_sums[3][56] [5:0] }), .sum({ \level_2_sums[3][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[117] [4:0] }), .sum({ \level_1_sums[3][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[119] [4:0] }), .sum({ \level_1_sums[3][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[3][59] [5:0] }),
     .b({ \level_1_sums[3][58] [5:0] }), .sum({ \level_2_sums[3][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[3][29] [6:0] }),
     .b({ \level_2_sums[3][28] [6:0] }), .sum({ \level_3_sums[3][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[121] [4:0] }), .sum({ \level_1_sums[3][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[123] [4:0] }), .sum({ \level_1_sums[3][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[3][61] [5:0] }),
     .b({ \level_1_sums[3][60] [5:0] }), .sum({ \level_2_sums[3][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[125] [4:0] }), .sum({ \level_1_sums[3][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[127] [4:0] }), .sum({ \level_1_sums[3][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[3][63] [5:0] }),
     .b({ \level_1_sums[3][62] [5:0] }), .sum({ \level_2_sums[3][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[3][31] [6:0] }),
     .b({ \level_2_sums[3][30] [6:0] }), .sum({ \level_3_sums[3][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[3][15] [7:0] }),
     .b({ \level_3_sums[3][14] [7:0] }), .sum({ \level_4_sums[3][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[3][7] [8:0] }),
     .b({ \level_4_sums[3][6] [8:0] }), .sum({ \level_5_sums[3][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[3][3] [9:0] }),
     .b({ \level_5_sums[3][2] [9:0] }), .sum({ \level_6_sums[3][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[3][1] [9:0] }),
     .b({ \level_6_sums[3][0] [9:0] }), .sum({ \level_7_sums[3][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[129] [4:0] }), .sum({ \level_1_sums[3][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[131] [4:0] }), .sum({ \level_1_sums[3][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[3][65] [5:0] }),
     .b({ \level_1_sums[3][64] [5:0] }), .sum({ \level_2_sums[3][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[133] [4:0] }), .sum({ \level_1_sums[3][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[135] [4:0] }), .sum({ \level_1_sums[3][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[3][67] [5:0] }),
     .b({ \level_1_sums[3][66] [5:0] }), .sum({ \level_2_sums[3][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[3][33] [6:0] }),
     .b({ \level_2_sums[3][32] [6:0] }), .sum({ \level_3_sums[3][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[137] [4:0] }), .sum({ \level_1_sums[3][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[139] [4:0] }), .sum({ \level_1_sums[3][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[3][69] [5:0] }),
     .b({ \level_1_sums[3][68] [5:0] }), .sum({ \level_2_sums[3][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[141] [4:0] }), .sum({ \level_1_sums[3][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[143] [4:0] }), .sum({ \level_1_sums[3][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[3][71] [5:0] }),
     .b({ \level_1_sums[3][70] [5:0] }), .sum({ \level_2_sums[3][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[3][35] [6:0] }),
     .b({ \level_2_sums[3][34] [6:0] }), .sum({ \level_3_sums[3][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[3][17] [7:0] }),
     .b({ \level_3_sums[3][16] [7:0] }), .sum({ \level_4_sums[3][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[145] [4:0] }), .sum({ \level_1_sums[3][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[147] [4:0] }), .sum({ \level_1_sums[3][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[3][73] [5:0] }),
     .b({ \level_1_sums[3][72] [5:0] }), .sum({ \level_2_sums[3][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[149] [4:0] }), .sum({ \level_1_sums[3][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[151] [4:0] }), .sum({ \level_1_sums[3][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[3][75] [5:0] }),
     .b({ \level_1_sums[3][74] [5:0] }), .sum({ \level_2_sums[3][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[3][37] [6:0] }),
     .b({ \level_2_sums[3][36] [6:0] }), .sum({ \level_3_sums[3][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[153] [4:0] }), .sum({ \level_1_sums[3][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[155] [4:0] }), .sum({ \level_1_sums[3][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[3][77] [5:0] }),
     .b({ \level_1_sums[3][76] [5:0] }), .sum({ \level_2_sums[3][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[157] [4:0] }), .sum({ \level_1_sums[3][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[159] [4:0] }), .sum({ \level_1_sums[3][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[3][79] [5:0] }),
     .b({ \level_1_sums[3][78] [5:0] }), .sum({ \level_2_sums[3][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[3][39] [6:0] }),
     .b({ \level_2_sums[3][38] [6:0] }), .sum({ \level_3_sums[3][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[3][19] [7:0] }),
     .b({ \level_3_sums[3][18] [7:0] }), .sum({ \level_4_sums[3][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[3][9] [8:0] }),
     .b({ \level_4_sums[3][8] [8:0] }), .sum({ \level_5_sums[3][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[161] [4:0] }), .sum({ \level_1_sums[3][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[163] [4:0] }), .sum({ \level_1_sums[3][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[3][81] [5:0] }),
     .b({ \level_1_sums[3][80] [5:0] }), .sum({ \level_2_sums[3][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[165] [4:0] }), .sum({ \level_1_sums[3][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[167] [4:0] }), .sum({ \level_1_sums[3][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[3][83] [5:0] }),
     .b({ \level_1_sums[3][82] [5:0] }), .sum({ \level_2_sums[3][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[3][41] [6:0] }),
     .b({ \level_2_sums[3][40] [6:0] }), .sum({ \level_3_sums[3][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[169] [4:0] }), .sum({ \level_1_sums[3][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[171] [4:0] }), .sum({ \level_1_sums[3][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[3][85] [5:0] }),
     .b({ \level_1_sums[3][84] [5:0] }), .sum({ \level_2_sums[3][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[173] [4:0] }), .sum({ \level_1_sums[3][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[175] [4:0] }), .sum({ \level_1_sums[3][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[3][87] [5:0] }),
     .b({ \level_1_sums[3][86] [5:0] }), .sum({ \level_2_sums[3][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[3][43] [6:0] }),
     .b({ \level_2_sums[3][42] [6:0] }), .sum({ \level_3_sums[3][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[3][21] [7:0] }),
     .b({ \level_3_sums[3][20] [7:0] }), .sum({ \level_4_sums[3][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[177] [4:0] }), .sum({ \level_1_sums[3][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[179] [4:0] }), .sum({ \level_1_sums[3][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[3][89] [5:0] }),
     .b({ \level_1_sums[3][88] [5:0] }), .sum({ \level_2_sums[3][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[181] [4:0] }), .sum({ \level_1_sums[3][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[183] [4:0] }), .sum({ \level_1_sums[3][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[3][91] [5:0] }),
     .b({ \level_1_sums[3][90] [5:0] }), .sum({ \level_2_sums[3][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[3][45] [6:0] }),
     .b({ \level_2_sums[3][44] [6:0] }), .sum({ \level_3_sums[3][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[185] [4:0] }), .sum({ \level_1_sums[3][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[187] [4:0] }), .sum({ \level_1_sums[3][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[3][93] [5:0] }),
     .b({ \level_1_sums[3][92] [5:0] }), .sum({ \level_2_sums[3][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[189] [4:0] }), .sum({ \level_1_sums[3][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[191] [4:0] }), .sum({ \level_1_sums[3][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[3][95] [5:0] }),
     .b({ \level_1_sums[3][94] [5:0] }), .sum({ \level_2_sums[3][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[3][47] [6:0] }),
     .b({ \level_2_sums[3][46] [6:0] }), .sum({ \level_3_sums[3][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[3][23] [7:0] }),
     .b({ \level_3_sums[3][22] [7:0] }), .sum({ \level_4_sums[3][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[3][11] [8:0] }),
     .b({ \level_4_sums[3][10] [8:0] }), .sum({ \level_5_sums[3][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[3][5] [9:0] }),
     .b({ \level_5_sums[3][4] [9:0] }), .sum({ \level_6_sums[3][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[193] [4:0] }), .sum({ \level_1_sums[3][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[195] [4:0] }), .sum({ \level_1_sums[3][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[3][97] [5:0] }),
     .b({ \level_1_sums[3][96] [5:0] }), .sum({ \level_2_sums[3][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[197] [4:0] }), .sum({ \level_1_sums[3][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[199] [4:0] }), .sum({ \level_1_sums[3][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[3][99] [5:0] }),
     .b({ \level_1_sums[3][98] [5:0] }), .sum({ \level_2_sums[3][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[3][49] [6:0] }),
     .b({ \level_2_sums[3][48] [6:0] }), .sum({ \level_3_sums[3][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[201] [4:0] }), .sum({ \level_1_sums[3][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[203] [4:0] }), .sum({ \level_1_sums[3][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[3][101] [5:0] }),
     .b({ \level_1_sums[3][100] [5:0] }), .sum({ \level_2_sums[3][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[205] [4:0] }), .sum({ \level_1_sums[3][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[207] [4:0] }), .sum({ \level_1_sums[3][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[3][103] [5:0] }),
     .b({ \level_1_sums[3][102] [5:0] }), .sum({ \level_2_sums[3][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[3][51] [6:0] }),
     .b({ \level_2_sums[3][50] [6:0] }), .sum({ \level_3_sums[3][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[3][25] [7:0] }),
     .b({ \level_3_sums[3][24] [7:0] }), .sum({ \level_4_sums[3][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[209] [4:0] }), .sum({ \level_1_sums[3][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[211] [4:0] }), .sum({ \level_1_sums[3][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[3][105] [5:0] }),
     .b({ \level_1_sums[3][104] [5:0] }), .sum({ \level_2_sums[3][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[213] [4:0] }), .sum({ \level_1_sums[3][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[215] [4:0] }), .sum({ \level_1_sums[3][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[3][107] [5:0] }),
     .b({ \level_1_sums[3][106] [5:0] }), .sum({ \level_2_sums[3][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[3][53] [6:0] }),
     .b({ \level_2_sums[3][52] [6:0] }), .sum({ \level_3_sums[3][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[217] [4:0] }), .sum({ \level_1_sums[3][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[219] [4:0] }), .sum({ \level_1_sums[3][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[3][109] [5:0] }),
     .b({ \level_1_sums[3][108] [5:0] }), .sum({ \level_2_sums[3][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[221] [4:0] }), .sum({ \level_1_sums[3][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[223] [4:0] }), .sum({ \level_1_sums[3][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[3][111] [5:0] }),
     .b({ \level_1_sums[3][110] [5:0] }), .sum({ \level_2_sums[3][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[3][55] [6:0] }),
     .b({ \level_2_sums[3][54] [6:0] }), .sum({ \level_3_sums[3][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[3][27] [7:0] }),
     .b({ \level_3_sums[3][26] [7:0] }), .sum({ \level_4_sums[3][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[3][13] [8:0] }),
     .b({ \level_4_sums[3][12] [8:0] }), .sum({ \level_5_sums[3][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[225] [4:0] }), .sum({ \level_1_sums[3][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[227] [4:0] }), .sum({ \level_1_sums[3][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[3][113] [5:0] }),
     .b({ \level_1_sums[3][112] [5:0] }), .sum({ \level_2_sums[3][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[229] [4:0] }), .sum({ \level_1_sums[3][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[231] [4:0] }), .sum({ \level_1_sums[3][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[3][115] [5:0] }),
     .b({ \level_1_sums[3][114] [5:0] }), .sum({ \level_2_sums[3][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[3][57] [6:0] }),
     .b({ \level_2_sums[3][56] [6:0] }), .sum({ \level_3_sums[3][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[233] [4:0] }), .sum({ \level_1_sums[3][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[235] [4:0] }), .sum({ \level_1_sums[3][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[3][117] [5:0] }),
     .b({ \level_1_sums[3][116] [5:0] }), .sum({ \level_2_sums[3][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[237] [4:0] }), .sum({ \level_1_sums[3][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[239] [4:0] }), .sum({ \level_1_sums[3][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[3][119] [5:0] }),
     .b({ \level_1_sums[3][118] [5:0] }), .sum({ \level_2_sums[3][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[3][59] [6:0] }),
     .b({ \level_2_sums[3][58] [6:0] }), .sum({ \level_3_sums[3][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[3][29] [7:0] }),
     .b({ \level_3_sums[3][28] [7:0] }), .sum({ \level_4_sums[3][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[241] [4:0] }), .sum({ \level_1_sums[3][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[243] [4:0] }), .sum({ \level_1_sums[3][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[3][121] [5:0] }),
     .b({ \level_1_sums[3][120] [5:0] }), .sum({ \level_2_sums[3][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[245] [4:0] }), .sum({ \level_1_sums[3][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[247] [4:0] }), .sum({ \level_1_sums[3][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[3][123] [5:0] }),
     .b({ \level_1_sums[3][122] [5:0] }), .sum({ \level_2_sums[3][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[3][61] [6:0] }),
     .b({ \level_2_sums[3][60] [6:0] }), .sum({ \level_3_sums[3][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[249] [4:0] }), .sum({ \level_1_sums[3][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[251] [4:0] }), .sum({ \level_1_sums[3][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[3][125] [5:0] }),
     .b({ \level_1_sums[3][124] [5:0] }), .sum({ \level_2_sums[3][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[253] [4:0] }), .sum({ \level_1_sums[3][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[3].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[3].product_terms[255] [4:0] }), .sum({ \level_1_sums[3][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[3][127] [5:0] }),
     .b({ \level_1_sums[3][126] [5:0] }), .sum({ \level_2_sums[3][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[3][63] [6:0] }),
     .b({ \level_2_sums[3][62] [6:0] }), .sum({ \level_3_sums[3][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[3][31] [7:0] }),
     .b({ \level_3_sums[3][30] [7:0] }), .sum({ \level_4_sums[3][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[3][15] [8:0] }),
     .b({ \level_4_sums[3][14] [8:0] }), .sum({ \level_5_sums[3][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[3][7] [9:0] }),
     .b({ \level_5_sums[3][6] [9:0] }), .sum({ \level_6_sums[3][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[3][3] [9:0] }),
     .b({ \level_6_sums[3][2] [9:0] }), .sum({ \level_7_sums[3][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[3].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[3][0] [9:0] }),
     .b({ \level_7_sums[3][1] [9:0] }), .sum({ \level_8_sums[3] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[4].relu_inst (.in_data({ \final_sums[4] [9:0] }), .out_data({ \out_sig[4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[1] [4:0] }), .sum({ \level_1_sums[4][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[3] [4:0] }), .sum({ \level_1_sums[4][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[4][1] [5:0] }),
     .b({ \level_1_sums[4][0] [5:0] }), .sum({ \level_2_sums[4][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[5] [4:0] }), .sum({ \level_1_sums[4][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[7] [4:0] }), .sum({ \level_1_sums[4][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[4][3] [5:0] }),
     .b({ \level_1_sums[4][2] [5:0] }), .sum({ \level_2_sums[4][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[4][1] [6:0] }),
     .b({ \level_2_sums[4][0] [6:0] }), .sum({ \level_3_sums[4][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[9] [4:0] }), .sum({ \level_1_sums[4][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[11] [4:0] }), .sum({ \level_1_sums[4][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[4][5] [5:0] }),
     .b({ \level_1_sums[4][4] [5:0] }), .sum({ \level_2_sums[4][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[13] [4:0] }), .sum({ \level_1_sums[4][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[15] [4:0] }), .sum({ \level_1_sums[4][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[4][7] [5:0] }),
     .b({ \level_1_sums[4][6] [5:0] }), .sum({ \level_2_sums[4][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[4][3] [6:0] }),
     .b({ \level_2_sums[4][2] [6:0] }), .sum({ \level_3_sums[4][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[4][1] [7:0] }),
     .b({ \level_3_sums[4][0] [7:0] }), .sum({ \level_4_sums[4][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[17] [4:0] }), .sum({ \level_1_sums[4][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[19] [4:0] }), .sum({ \level_1_sums[4][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[4][9] [5:0] }),
     .b({ \level_1_sums[4][8] [5:0] }), .sum({ \level_2_sums[4][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[21] [4:0] }), .sum({ \level_1_sums[4][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[23] [4:0] }), .sum({ \level_1_sums[4][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[4][11] [5:0] }),
     .b({ \level_1_sums[4][10] [5:0] }), .sum({ \level_2_sums[4][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[4][5] [6:0] }),
     .b({ \level_2_sums[4][4] [6:0] }), .sum({ \level_3_sums[4][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[25] [4:0] }), .sum({ \level_1_sums[4][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[27] [4:0] }), .sum({ \level_1_sums[4][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[4][13] [5:0] }),
     .b({ \level_1_sums[4][12] [5:0] }), .sum({ \level_2_sums[4][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[29] [4:0] }), .sum({ \level_1_sums[4][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[31] [4:0] }), .sum({ \level_1_sums[4][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[4][15] [5:0] }),
     .b({ \level_1_sums[4][14] [5:0] }), .sum({ \level_2_sums[4][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[4][7] [6:0] }),
     .b({ \level_2_sums[4][6] [6:0] }), .sum({ \level_3_sums[4][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[4][3] [7:0] }),
     .b({ \level_3_sums[4][2] [7:0] }), .sum({ \level_4_sums[4][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[4][1] [8:0] }),
     .b({ \level_4_sums[4][0] [8:0] }), .sum({ \level_5_sums[4][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[33] [4:0] }), .sum({ \level_1_sums[4][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[35] [4:0] }), .sum({ \level_1_sums[4][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[4][17] [5:0] }),
     .b({ \level_1_sums[4][16] [5:0] }), .sum({ \level_2_sums[4][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[37] [4:0] }), .sum({ \level_1_sums[4][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[39] [4:0] }), .sum({ \level_1_sums[4][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[4][19] [5:0] }),
     .b({ \level_1_sums[4][18] [5:0] }), .sum({ \level_2_sums[4][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[4][9] [6:0] }),
     .b({ \level_2_sums[4][8] [6:0] }), .sum({ \level_3_sums[4][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[41] [4:0] }), .sum({ \level_1_sums[4][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[43] [4:0] }), .sum({ \level_1_sums[4][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[4][21] [5:0] }),
     .b({ \level_1_sums[4][20] [5:0] }), .sum({ \level_2_sums[4][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[45] [4:0] }), .sum({ \level_1_sums[4][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[47] [4:0] }), .sum({ \level_1_sums[4][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[4][23] [5:0] }),
     .b({ \level_1_sums[4][22] [5:0] }), .sum({ \level_2_sums[4][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[4][11] [6:0] }),
     .b({ \level_2_sums[4][10] [6:0] }), .sum({ \level_3_sums[4][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[4][5] [7:0] }),
     .b({ \level_3_sums[4][4] [7:0] }), .sum({ \level_4_sums[4][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[49] [4:0] }), .sum({ \level_1_sums[4][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[51] [4:0] }), .sum({ \level_1_sums[4][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[4][25] [5:0] }),
     .b({ \level_1_sums[4][24] [5:0] }), .sum({ \level_2_sums[4][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[53] [4:0] }), .sum({ \level_1_sums[4][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[55] [4:0] }), .sum({ \level_1_sums[4][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[4][27] [5:0] }),
     .b({ \level_1_sums[4][26] [5:0] }), .sum({ \level_2_sums[4][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[4][13] [6:0] }),
     .b({ \level_2_sums[4][12] [6:0] }), .sum({ \level_3_sums[4][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[57] [4:0] }), .sum({ \level_1_sums[4][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[59] [4:0] }), .sum({ \level_1_sums[4][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[4][29] [5:0] }),
     .b({ \level_1_sums[4][28] [5:0] }), .sum({ \level_2_sums[4][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[61] [4:0] }), .sum({ \level_1_sums[4][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[63] [4:0] }), .sum({ \level_1_sums[4][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[4][31] [5:0] }),
     .b({ \level_1_sums[4][30] [5:0] }), .sum({ \level_2_sums[4][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[4][15] [6:0] }),
     .b({ \level_2_sums[4][14] [6:0] }), .sum({ \level_3_sums[4][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[4][7] [7:0] }),
     .b({ \level_3_sums[4][6] [7:0] }), .sum({ \level_4_sums[4][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[4][3] [8:0] }),
     .b({ \level_4_sums[4][2] [8:0] }), .sum({ \level_5_sums[4][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[4][1] [9:0] }),
     .b({ \level_5_sums[4][0] [9:0] }), .sum({ \level_6_sums[4][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[65] [4:0] }), .sum({ \level_1_sums[4][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[67] [4:0] }), .sum({ \level_1_sums[4][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[4][33] [5:0] }),
     .b({ \level_1_sums[4][32] [5:0] }), .sum({ \level_2_sums[4][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[69] [4:0] }), .sum({ \level_1_sums[4][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[71] [4:0] }), .sum({ \level_1_sums[4][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[4][35] [5:0] }),
     .b({ \level_1_sums[4][34] [5:0] }), .sum({ \level_2_sums[4][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[4][17] [6:0] }),
     .b({ \level_2_sums[4][16] [6:0] }), .sum({ \level_3_sums[4][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[73] [4:0] }), .sum({ \level_1_sums[4][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[75] [4:0] }), .sum({ \level_1_sums[4][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[4][37] [5:0] }),
     .b({ \level_1_sums[4][36] [5:0] }), .sum({ \level_2_sums[4][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[77] [4:0] }), .sum({ \level_1_sums[4][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[79] [4:0] }), .sum({ \level_1_sums[4][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[4][39] [5:0] }),
     .b({ \level_1_sums[4][38] [5:0] }), .sum({ \level_2_sums[4][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[4][19] [6:0] }),
     .b({ \level_2_sums[4][18] [6:0] }), .sum({ \level_3_sums[4][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[4][9] [7:0] }),
     .b({ \level_3_sums[4][8] [7:0] }), .sum({ \level_4_sums[4][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[81] [4:0] }), .sum({ \level_1_sums[4][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[83] [4:0] }), .sum({ \level_1_sums[4][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[4][41] [5:0] }),
     .b({ \level_1_sums[4][40] [5:0] }), .sum({ \level_2_sums[4][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[85] [4:0] }), .sum({ \level_1_sums[4][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[87] [4:0] }), .sum({ \level_1_sums[4][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[4][43] [5:0] }),
     .b({ \level_1_sums[4][42] [5:0] }), .sum({ \level_2_sums[4][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[4][21] [6:0] }),
     .b({ \level_2_sums[4][20] [6:0] }), .sum({ \level_3_sums[4][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[89] [4:0] }), .sum({ \level_1_sums[4][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[91] [4:0] }), .sum({ \level_1_sums[4][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[4][45] [5:0] }),
     .b({ \level_1_sums[4][44] [5:0] }), .sum({ \level_2_sums[4][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[93] [4:0] }), .sum({ \level_1_sums[4][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[95] [4:0] }), .sum({ \level_1_sums[4][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[4][47] [5:0] }),
     .b({ \level_1_sums[4][46] [5:0] }), .sum({ \level_2_sums[4][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[4][23] [6:0] }),
     .b({ \level_2_sums[4][22] [6:0] }), .sum({ \level_3_sums[4][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[4][11] [7:0] }),
     .b({ \level_3_sums[4][10] [7:0] }), .sum({ \level_4_sums[4][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[4][5] [8:0] }),
     .b({ \level_4_sums[4][4] [8:0] }), .sum({ \level_5_sums[4][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[97] [4:0] }), .sum({ \level_1_sums[4][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[99] [4:0] }), .sum({ \level_1_sums[4][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[4][49] [5:0] }),
     .b({ \level_1_sums[4][48] [5:0] }), .sum({ \level_2_sums[4][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[101] [4:0] }), .sum({ \level_1_sums[4][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[103] [4:0] }), .sum({ \level_1_sums[4][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[4][51] [5:0] }),
     .b({ \level_1_sums[4][50] [5:0] }), .sum({ \level_2_sums[4][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[4][25] [6:0] }),
     .b({ \level_2_sums[4][24] [6:0] }), .sum({ \level_3_sums[4][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[105] [4:0] }), .sum({ \level_1_sums[4][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[107] [4:0] }), .sum({ \level_1_sums[4][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[4][53] [5:0] }),
     .b({ \level_1_sums[4][52] [5:0] }), .sum({ \level_2_sums[4][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[109] [4:0] }), .sum({ \level_1_sums[4][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[111] [4:0] }), .sum({ \level_1_sums[4][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[4][55] [5:0] }),
     .b({ \level_1_sums[4][54] [5:0] }), .sum({ \level_2_sums[4][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[4][27] [6:0] }),
     .b({ \level_2_sums[4][26] [6:0] }), .sum({ \level_3_sums[4][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[4][13] [7:0] }),
     .b({ \level_3_sums[4][12] [7:0] }), .sum({ \level_4_sums[4][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[113] [4:0] }), .sum({ \level_1_sums[4][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[115] [4:0] }), .sum({ \level_1_sums[4][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[4][57] [5:0] }),
     .b({ \level_1_sums[4][56] [5:0] }), .sum({ \level_2_sums[4][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[117] [4:0] }), .sum({ \level_1_sums[4][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[119] [4:0] }), .sum({ \level_1_sums[4][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[4][59] [5:0] }),
     .b({ \level_1_sums[4][58] [5:0] }), .sum({ \level_2_sums[4][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[4][29] [6:0] }),
     .b({ \level_2_sums[4][28] [6:0] }), .sum({ \level_3_sums[4][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[121] [4:0] }), .sum({ \level_1_sums[4][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[123] [4:0] }), .sum({ \level_1_sums[4][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[4][61] [5:0] }),
     .b({ \level_1_sums[4][60] [5:0] }), .sum({ \level_2_sums[4][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[125] [4:0] }), .sum({ \level_1_sums[4][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[127] [4:0] }), .sum({ \level_1_sums[4][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[4][63] [5:0] }),
     .b({ \level_1_sums[4][62] [5:0] }), .sum({ \level_2_sums[4][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[4][31] [6:0] }),
     .b({ \level_2_sums[4][30] [6:0] }), .sum({ \level_3_sums[4][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[4][15] [7:0] }),
     .b({ \level_3_sums[4][14] [7:0] }), .sum({ \level_4_sums[4][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[4][7] [8:0] }),
     .b({ \level_4_sums[4][6] [8:0] }), .sum({ \level_5_sums[4][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[4][3] [9:0] }),
     .b({ \level_5_sums[4][2] [9:0] }), .sum({ \level_6_sums[4][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[4][1] [9:0] }),
     .b({ \level_6_sums[4][0] [9:0] }), .sum({ \level_7_sums[4][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[129] [4:0] }), .sum({ \level_1_sums[4][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[131] [4:0] }), .sum({ \level_1_sums[4][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[4][65] [5:0] }),
     .b({ \level_1_sums[4][64] [5:0] }), .sum({ \level_2_sums[4][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[133] [4:0] }), .sum({ \level_1_sums[4][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[135] [4:0] }), .sum({ \level_1_sums[4][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[4][67] [5:0] }),
     .b({ \level_1_sums[4][66] [5:0] }), .sum({ \level_2_sums[4][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[4][33] [6:0] }),
     .b({ \level_2_sums[4][32] [6:0] }), .sum({ \level_3_sums[4][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[137] [4:0] }), .sum({ \level_1_sums[4][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[139] [4:0] }), .sum({ \level_1_sums[4][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[4][69] [5:0] }),
     .b({ \level_1_sums[4][68] [5:0] }), .sum({ \level_2_sums[4][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[141] [4:0] }), .sum({ \level_1_sums[4][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[143] [4:0] }), .sum({ \level_1_sums[4][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[4][71] [5:0] }),
     .b({ \level_1_sums[4][70] [5:0] }), .sum({ \level_2_sums[4][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[4][35] [6:0] }),
     .b({ \level_2_sums[4][34] [6:0] }), .sum({ \level_3_sums[4][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[4][17] [7:0] }),
     .b({ \level_3_sums[4][16] [7:0] }), .sum({ \level_4_sums[4][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[145] [4:0] }), .sum({ \level_1_sums[4][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[147] [4:0] }), .sum({ \level_1_sums[4][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[4][73] [5:0] }),
     .b({ \level_1_sums[4][72] [5:0] }), .sum({ \level_2_sums[4][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[149] [4:0] }), .sum({ \level_1_sums[4][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[151] [4:0] }), .sum({ \level_1_sums[4][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[4][75] [5:0] }),
     .b({ \level_1_sums[4][74] [5:0] }), .sum({ \level_2_sums[4][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[4][37] [6:0] }),
     .b({ \level_2_sums[4][36] [6:0] }), .sum({ \level_3_sums[4][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[153] [4:0] }), .sum({ \level_1_sums[4][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[155] [4:0] }), .sum({ \level_1_sums[4][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[4][77] [5:0] }),
     .b({ \level_1_sums[4][76] [5:0] }), .sum({ \level_2_sums[4][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[157] [4:0] }), .sum({ \level_1_sums[4][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[159] [4:0] }), .sum({ \level_1_sums[4][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[4][79] [5:0] }),
     .b({ \level_1_sums[4][78] [5:0] }), .sum({ \level_2_sums[4][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[4][39] [6:0] }),
     .b({ \level_2_sums[4][38] [6:0] }), .sum({ \level_3_sums[4][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[4][19] [7:0] }),
     .b({ \level_3_sums[4][18] [7:0] }), .sum({ \level_4_sums[4][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[4][9] [8:0] }),
     .b({ \level_4_sums[4][8] [8:0] }), .sum({ \level_5_sums[4][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[161] [4:0] }), .sum({ \level_1_sums[4][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[163] [4:0] }), .sum({ \level_1_sums[4][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[4][81] [5:0] }),
     .b({ \level_1_sums[4][80] [5:0] }), .sum({ \level_2_sums[4][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[165] [4:0] }), .sum({ \level_1_sums[4][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[167] [4:0] }), .sum({ \level_1_sums[4][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[4][83] [5:0] }),
     .b({ \level_1_sums[4][82] [5:0] }), .sum({ \level_2_sums[4][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[4][41] [6:0] }),
     .b({ \level_2_sums[4][40] [6:0] }), .sum({ \level_3_sums[4][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[169] [4:0] }), .sum({ \level_1_sums[4][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[171] [4:0] }), .sum({ \level_1_sums[4][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[4][85] [5:0] }),
     .b({ \level_1_sums[4][84] [5:0] }), .sum({ \level_2_sums[4][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[173] [4:0] }), .sum({ \level_1_sums[4][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[175] [4:0] }), .sum({ \level_1_sums[4][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[4][87] [5:0] }),
     .b({ \level_1_sums[4][86] [5:0] }), .sum({ \level_2_sums[4][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[4][43] [6:0] }),
     .b({ \level_2_sums[4][42] [6:0] }), .sum({ \level_3_sums[4][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[4][21] [7:0] }),
     .b({ \level_3_sums[4][20] [7:0] }), .sum({ \level_4_sums[4][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[177] [4:0] }), .sum({ \level_1_sums[4][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[179] [4:0] }), .sum({ \level_1_sums[4][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[4][89] [5:0] }),
     .b({ \level_1_sums[4][88] [5:0] }), .sum({ \level_2_sums[4][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[181] [4:0] }), .sum({ \level_1_sums[4][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[183] [4:0] }), .sum({ \level_1_sums[4][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[4][91] [5:0] }),
     .b({ \level_1_sums[4][90] [5:0] }), .sum({ \level_2_sums[4][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[4][45] [6:0] }),
     .b({ \level_2_sums[4][44] [6:0] }), .sum({ \level_3_sums[4][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[185] [4:0] }), .sum({ \level_1_sums[4][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[187] [4:0] }), .sum({ \level_1_sums[4][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[4][93] [5:0] }),
     .b({ \level_1_sums[4][92] [5:0] }), .sum({ \level_2_sums[4][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[189] [4:0] }), .sum({ \level_1_sums[4][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[191] [4:0] }), .sum({ \level_1_sums[4][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[4][95] [5:0] }),
     .b({ \level_1_sums[4][94] [5:0] }), .sum({ \level_2_sums[4][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[4][47] [6:0] }),
     .b({ \level_2_sums[4][46] [6:0] }), .sum({ \level_3_sums[4][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[4][23] [7:0] }),
     .b({ \level_3_sums[4][22] [7:0] }), .sum({ \level_4_sums[4][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[4][11] [8:0] }),
     .b({ \level_4_sums[4][10] [8:0] }), .sum({ \level_5_sums[4][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[4][5] [9:0] }),
     .b({ \level_5_sums[4][4] [9:0] }), .sum({ \level_6_sums[4][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[193] [4:0] }), .sum({ \level_1_sums[4][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[195] [4:0] }), .sum({ \level_1_sums[4][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[4][97] [5:0] }),
     .b({ \level_1_sums[4][96] [5:0] }), .sum({ \level_2_sums[4][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[197] [4:0] }), .sum({ \level_1_sums[4][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[199] [4:0] }), .sum({ \level_1_sums[4][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[4][99] [5:0] }),
     .b({ \level_1_sums[4][98] [5:0] }), .sum({ \level_2_sums[4][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[4][49] [6:0] }),
     .b({ \level_2_sums[4][48] [6:0] }), .sum({ \level_3_sums[4][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[201] [4:0] }), .sum({ \level_1_sums[4][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[203] [4:0] }), .sum({ \level_1_sums[4][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[4][101] [5:0] }),
     .b({ \level_1_sums[4][100] [5:0] }), .sum({ \level_2_sums[4][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[205] [4:0] }), .sum({ \level_1_sums[4][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[207] [4:0] }), .sum({ \level_1_sums[4][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[4][103] [5:0] }),
     .b({ \level_1_sums[4][102] [5:0] }), .sum({ \level_2_sums[4][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[4][51] [6:0] }),
     .b({ \level_2_sums[4][50] [6:0] }), .sum({ \level_3_sums[4][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[4][25] [7:0] }),
     .b({ \level_3_sums[4][24] [7:0] }), .sum({ \level_4_sums[4][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[209] [4:0] }), .sum({ \level_1_sums[4][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[211] [4:0] }), .sum({ \level_1_sums[4][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[4][105] [5:0] }),
     .b({ \level_1_sums[4][104] [5:0] }), .sum({ \level_2_sums[4][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[213] [4:0] }), .sum({ \level_1_sums[4][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[215] [4:0] }), .sum({ \level_1_sums[4][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[4][107] [5:0] }),
     .b({ \level_1_sums[4][106] [5:0] }), .sum({ \level_2_sums[4][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[4][53] [6:0] }),
     .b({ \level_2_sums[4][52] [6:0] }), .sum({ \level_3_sums[4][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[217] [4:0] }), .sum({ \level_1_sums[4][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[219] [4:0] }), .sum({ \level_1_sums[4][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[4][109] [5:0] }),
     .b({ \level_1_sums[4][108] [5:0] }), .sum({ \level_2_sums[4][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[221] [4:0] }), .sum({ \level_1_sums[4][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[223] [4:0] }), .sum({ \level_1_sums[4][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[4][111] [5:0] }),
     .b({ \level_1_sums[4][110] [5:0] }), .sum({ \level_2_sums[4][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[4][55] [6:0] }),
     .b({ \level_2_sums[4][54] [6:0] }), .sum({ \level_3_sums[4][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[4][27] [7:0] }),
     .b({ \level_3_sums[4][26] [7:0] }), .sum({ \level_4_sums[4][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[4][13] [8:0] }),
     .b({ \level_4_sums[4][12] [8:0] }), .sum({ \level_5_sums[4][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[225] [4:0] }), .sum({ \level_1_sums[4][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[227] [4:0] }), .sum({ \level_1_sums[4][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[4][113] [5:0] }),
     .b({ \level_1_sums[4][112] [5:0] }), .sum({ \level_2_sums[4][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[229] [4:0] }), .sum({ \level_1_sums[4][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[231] [4:0] }), .sum({ \level_1_sums[4][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[4][115] [5:0] }),
     .b({ \level_1_sums[4][114] [5:0] }), .sum({ \level_2_sums[4][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[4][57] [6:0] }),
     .b({ \level_2_sums[4][56] [6:0] }), .sum({ \level_3_sums[4][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[233] [4:0] }), .sum({ \level_1_sums[4][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[235] [4:0] }), .sum({ \level_1_sums[4][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[4][117] [5:0] }),
     .b({ \level_1_sums[4][116] [5:0] }), .sum({ \level_2_sums[4][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[237] [4:0] }), .sum({ \level_1_sums[4][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[239] [4:0] }), .sum({ \level_1_sums[4][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[4][119] [5:0] }),
     .b({ \level_1_sums[4][118] [5:0] }), .sum({ \level_2_sums[4][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[4][59] [6:0] }),
     .b({ \level_2_sums[4][58] [6:0] }), .sum({ \level_3_sums[4][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[4][29] [7:0] }),
     .b({ \level_3_sums[4][28] [7:0] }), .sum({ \level_4_sums[4][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[241] [4:0] }), .sum({ \level_1_sums[4][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[243] [4:0] }), .sum({ \level_1_sums[4][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[4][121] [5:0] }),
     .b({ \level_1_sums[4][120] [5:0] }), .sum({ \level_2_sums[4][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[245] [4:0] }), .sum({ \level_1_sums[4][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[247] [4:0] }), .sum({ \level_1_sums[4][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[4][123] [5:0] }),
     .b({ \level_1_sums[4][122] [5:0] }), .sum({ \level_2_sums[4][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[4][61] [6:0] }),
     .b({ \level_2_sums[4][60] [6:0] }), .sum({ \level_3_sums[4][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[249] [4:0] }), .sum({ \level_1_sums[4][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[251] [4:0] }), .sum({ \level_1_sums[4][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[4][125] [5:0] }),
     .b({ \level_1_sums[4][124] [5:0] }), .sum({ \level_2_sums[4][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[253] [4:0] }), .sum({ \level_1_sums[4][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[4].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[4].product_terms[255] [4:0] }), .sum({ \level_1_sums[4][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[4][127] [5:0] }),
     .b({ \level_1_sums[4][126] [5:0] }), .sum({ \level_2_sums[4][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[4][63] [6:0] }),
     .b({ \level_2_sums[4][62] [6:0] }), .sum({ \level_3_sums[4][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[4][31] [7:0] }),
     .b({ \level_3_sums[4][30] [7:0] }), .sum({ \level_4_sums[4][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[4][15] [8:0] }),
     .b({ \level_4_sums[4][14] [8:0] }), .sum({ \level_5_sums[4][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[4][7] [9:0] }),
     .b({ \level_5_sums[4][6] [9:0] }), .sum({ \level_6_sums[4][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[4][3] [9:0] }),
     .b({ \level_6_sums[4][2] [9:0] }), .sum({ \level_7_sums[4][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[4].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[4][0] [9:0] }),
     .b({ \level_7_sums[4][1] [9:0] }), .sum({ \level_8_sums[4] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[5].relu_inst (.in_data({ \final_sums[5] [9:0] }), .out_data({ \out_sig[5] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[1] [4:0] }), .sum({ \level_1_sums[5][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[3] [4:0] }), .sum({ \level_1_sums[5][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[5][1] [5:0] }),
     .b({ \level_1_sums[5][0] [5:0] }), .sum({ \level_2_sums[5][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[5] [4:0] }), .sum({ \level_1_sums[5][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[7] [4:0] }), .sum({ \level_1_sums[5][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[5][3] [5:0] }),
     .b({ \level_1_sums[5][2] [5:0] }), .sum({ \level_2_sums[5][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[5][1] [6:0] }),
     .b({ \level_2_sums[5][0] [6:0] }), .sum({ \level_3_sums[5][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[9] [4:0] }), .sum({ \level_1_sums[5][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[11] [4:0] }), .sum({ \level_1_sums[5][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[5][5] [5:0] }),
     .b({ \level_1_sums[5][4] [5:0] }), .sum({ \level_2_sums[5][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[13] [4:0] }), .sum({ \level_1_sums[5][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[15] [4:0] }), .sum({ \level_1_sums[5][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[5][7] [5:0] }),
     .b({ \level_1_sums[5][6] [5:0] }), .sum({ \level_2_sums[5][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[5][3] [6:0] }),
     .b({ \level_2_sums[5][2] [6:0] }), .sum({ \level_3_sums[5][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[5][1] [7:0] }),
     .b({ \level_3_sums[5][0] [7:0] }), .sum({ \level_4_sums[5][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[17] [4:0] }), .sum({ \level_1_sums[5][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[19] [4:0] }), .sum({ \level_1_sums[5][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[5][9] [5:0] }),
     .b({ \level_1_sums[5][8] [5:0] }), .sum({ \level_2_sums[5][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[21] [4:0] }), .sum({ \level_1_sums[5][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[23] [4:0] }), .sum({ \level_1_sums[5][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[5][11] [5:0] }),
     .b({ \level_1_sums[5][10] [5:0] }), .sum({ \level_2_sums[5][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[5][5] [6:0] }),
     .b({ \level_2_sums[5][4] [6:0] }), .sum({ \level_3_sums[5][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[25] [4:0] }), .sum({ \level_1_sums[5][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[27] [4:0] }), .sum({ \level_1_sums[5][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[5][13] [5:0] }),
     .b({ \level_1_sums[5][12] [5:0] }), .sum({ \level_2_sums[5][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[29] [4:0] }), .sum({ \level_1_sums[5][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[31] [4:0] }), .sum({ \level_1_sums[5][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[5][15] [5:0] }),
     .b({ \level_1_sums[5][14] [5:0] }), .sum({ \level_2_sums[5][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[5][7] [6:0] }),
     .b({ \level_2_sums[5][6] [6:0] }), .sum({ \level_3_sums[5][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[5][3] [7:0] }),
     .b({ \level_3_sums[5][2] [7:0] }), .sum({ \level_4_sums[5][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[5][1] [8:0] }),
     .b({ \level_4_sums[5][0] [8:0] }), .sum({ \level_5_sums[5][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[33] [4:0] }), .sum({ \level_1_sums[5][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[35] [4:0] }), .sum({ \level_1_sums[5][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[5][17] [5:0] }),
     .b({ \level_1_sums[5][16] [5:0] }), .sum({ \level_2_sums[5][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[37] [4:0] }), .sum({ \level_1_sums[5][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[39] [4:0] }), .sum({ \level_1_sums[5][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[5][19] [5:0] }),
     .b({ \level_1_sums[5][18] [5:0] }), .sum({ \level_2_sums[5][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[5][9] [6:0] }),
     .b({ \level_2_sums[5][8] [6:0] }), .sum({ \level_3_sums[5][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[41] [4:0] }), .sum({ \level_1_sums[5][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[43] [4:0] }), .sum({ \level_1_sums[5][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[5][21] [5:0] }),
     .b({ \level_1_sums[5][20] [5:0] }), .sum({ \level_2_sums[5][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[45] [4:0] }), .sum({ \level_1_sums[5][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[47] [4:0] }), .sum({ \level_1_sums[5][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[5][23] [5:0] }),
     .b({ \level_1_sums[5][22] [5:0] }), .sum({ \level_2_sums[5][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[5][11] [6:0] }),
     .b({ \level_2_sums[5][10] [6:0] }), .sum({ \level_3_sums[5][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[5][5] [7:0] }),
     .b({ \level_3_sums[5][4] [7:0] }), .sum({ \level_4_sums[5][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[49] [4:0] }), .sum({ \level_1_sums[5][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[51] [4:0] }), .sum({ \level_1_sums[5][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[5][25] [5:0] }),
     .b({ \level_1_sums[5][24] [5:0] }), .sum({ \level_2_sums[5][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[53] [4:0] }), .sum({ \level_1_sums[5][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[55] [4:0] }), .sum({ \level_1_sums[5][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[5][27] [5:0] }),
     .b({ \level_1_sums[5][26] [5:0] }), .sum({ \level_2_sums[5][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[5][13] [6:0] }),
     .b({ \level_2_sums[5][12] [6:0] }), .sum({ \level_3_sums[5][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[57] [4:0] }), .sum({ \level_1_sums[5][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[59] [4:0] }), .sum({ \level_1_sums[5][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[5][29] [5:0] }),
     .b({ \level_1_sums[5][28] [5:0] }), .sum({ \level_2_sums[5][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[61] [4:0] }), .sum({ \level_1_sums[5][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[63] [4:0] }), .sum({ \level_1_sums[5][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[5][31] [5:0] }),
     .b({ \level_1_sums[5][30] [5:0] }), .sum({ \level_2_sums[5][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[5][15] [6:0] }),
     .b({ \level_2_sums[5][14] [6:0] }), .sum({ \level_3_sums[5][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[5][7] [7:0] }),
     .b({ \level_3_sums[5][6] [7:0] }), .sum({ \level_4_sums[5][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[5][3] [8:0] }),
     .b({ \level_4_sums[5][2] [8:0] }), .sum({ \level_5_sums[5][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[5][1] [9:0] }),
     .b({ \level_5_sums[5][0] [9:0] }), .sum({ \level_6_sums[5][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[65] [4:0] }), .sum({ \level_1_sums[5][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[67] [4:0] }), .sum({ \level_1_sums[5][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[5][33] [5:0] }),
     .b({ \level_1_sums[5][32] [5:0] }), .sum({ \level_2_sums[5][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[69] [4:0] }), .sum({ \level_1_sums[5][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[71] [4:0] }), .sum({ \level_1_sums[5][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[5][35] [5:0] }),
     .b({ \level_1_sums[5][34] [5:0] }), .sum({ \level_2_sums[5][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[5][17] [6:0] }),
     .b({ \level_2_sums[5][16] [6:0] }), .sum({ \level_3_sums[5][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[73] [4:0] }), .sum({ \level_1_sums[5][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[75] [4:0] }), .sum({ \level_1_sums[5][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[5][37] [5:0] }),
     .b({ \level_1_sums[5][36] [5:0] }), .sum({ \level_2_sums[5][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[77] [4:0] }), .sum({ \level_1_sums[5][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[79] [4:0] }), .sum({ \level_1_sums[5][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[5][39] [5:0] }),
     .b({ \level_1_sums[5][38] [5:0] }), .sum({ \level_2_sums[5][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[5][19] [6:0] }),
     .b({ \level_2_sums[5][18] [6:0] }), .sum({ \level_3_sums[5][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[5][9] [7:0] }),
     .b({ \level_3_sums[5][8] [7:0] }), .sum({ \level_4_sums[5][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[81] [4:0] }), .sum({ \level_1_sums[5][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[83] [4:0] }), .sum({ \level_1_sums[5][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[5][41] [5:0] }),
     .b({ \level_1_sums[5][40] [5:0] }), .sum({ \level_2_sums[5][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[85] [4:0] }), .sum({ \level_1_sums[5][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[87] [4:0] }), .sum({ \level_1_sums[5][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[5][43] [5:0] }),
     .b({ \level_1_sums[5][42] [5:0] }), .sum({ \level_2_sums[5][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[5][21] [6:0] }),
     .b({ \level_2_sums[5][20] [6:0] }), .sum({ \level_3_sums[5][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[89] [4:0] }), .sum({ \level_1_sums[5][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[91] [4:0] }), .sum({ \level_1_sums[5][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[5][45] [5:0] }),
     .b({ \level_1_sums[5][44] [5:0] }), .sum({ \level_2_sums[5][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[93] [4:0] }), .sum({ \level_1_sums[5][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[95] [4:0] }), .sum({ \level_1_sums[5][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[5][47] [5:0] }),
     .b({ \level_1_sums[5][46] [5:0] }), .sum({ \level_2_sums[5][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[5][23] [6:0] }),
     .b({ \level_2_sums[5][22] [6:0] }), .sum({ \level_3_sums[5][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[5][11] [7:0] }),
     .b({ \level_3_sums[5][10] [7:0] }), .sum({ \level_4_sums[5][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[5][5] [8:0] }),
     .b({ \level_4_sums[5][4] [8:0] }), .sum({ \level_5_sums[5][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[97] [4:0] }), .sum({ \level_1_sums[5][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[99] [4:0] }), .sum({ \level_1_sums[5][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[5][49] [5:0] }),
     .b({ \level_1_sums[5][48] [5:0] }), .sum({ \level_2_sums[5][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[101] [4:0] }), .sum({ \level_1_sums[5][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[103] [4:0] }), .sum({ \level_1_sums[5][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[5][51] [5:0] }),
     .b({ \level_1_sums[5][50] [5:0] }), .sum({ \level_2_sums[5][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[5][25] [6:0] }),
     .b({ \level_2_sums[5][24] [6:0] }), .sum({ \level_3_sums[5][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[105] [4:0] }), .sum({ \level_1_sums[5][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[107] [4:0] }), .sum({ \level_1_sums[5][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[5][53] [5:0] }),
     .b({ \level_1_sums[5][52] [5:0] }), .sum({ \level_2_sums[5][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[109] [4:0] }), .sum({ \level_1_sums[5][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[111] [4:0] }), .sum({ \level_1_sums[5][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[5][55] [5:0] }),
     .b({ \level_1_sums[5][54] [5:0] }), .sum({ \level_2_sums[5][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[5][27] [6:0] }),
     .b({ \level_2_sums[5][26] [6:0] }), .sum({ \level_3_sums[5][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[5][13] [7:0] }),
     .b({ \level_3_sums[5][12] [7:0] }), .sum({ \level_4_sums[5][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[113] [4:0] }), .sum({ \level_1_sums[5][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[115] [4:0] }), .sum({ \level_1_sums[5][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[5][57] [5:0] }),
     .b({ \level_1_sums[5][56] [5:0] }), .sum({ \level_2_sums[5][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[117] [4:0] }), .sum({ \level_1_sums[5][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[119] [4:0] }), .sum({ \level_1_sums[5][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[5][59] [5:0] }),
     .b({ \level_1_sums[5][58] [5:0] }), .sum({ \level_2_sums[5][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[5][29] [6:0] }),
     .b({ \level_2_sums[5][28] [6:0] }), .sum({ \level_3_sums[5][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[121] [4:0] }), .sum({ \level_1_sums[5][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[123] [4:0] }), .sum({ \level_1_sums[5][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[5][61] [5:0] }),
     .b({ \level_1_sums[5][60] [5:0] }), .sum({ \level_2_sums[5][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[125] [4:0] }), .sum({ \level_1_sums[5][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[127] [4:0] }), .sum({ \level_1_sums[5][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[5][63] [5:0] }),
     .b({ \level_1_sums[5][62] [5:0] }), .sum({ \level_2_sums[5][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[5][31] [6:0] }),
     .b({ \level_2_sums[5][30] [6:0] }), .sum({ \level_3_sums[5][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[5][15] [7:0] }),
     .b({ \level_3_sums[5][14] [7:0] }), .sum({ \level_4_sums[5][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[5][7] [8:0] }),
     .b({ \level_4_sums[5][6] [8:0] }), .sum({ \level_5_sums[5][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[5][3] [9:0] }),
     .b({ \level_5_sums[5][2] [9:0] }), .sum({ \level_6_sums[5][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[5][1] [9:0] }),
     .b({ \level_6_sums[5][0] [9:0] }), .sum({ \level_7_sums[5][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[129] [4:0] }), .sum({ \level_1_sums[5][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[131] [4:0] }), .sum({ \level_1_sums[5][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[5][65] [5:0] }),
     .b({ \level_1_sums[5][64] [5:0] }), .sum({ \level_2_sums[5][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[133] [4:0] }), .sum({ \level_1_sums[5][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[135] [4:0] }), .sum({ \level_1_sums[5][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[5][67] [5:0] }),
     .b({ \level_1_sums[5][66] [5:0] }), .sum({ \level_2_sums[5][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[5][33] [6:0] }),
     .b({ \level_2_sums[5][32] [6:0] }), .sum({ \level_3_sums[5][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[137] [4:0] }), .sum({ \level_1_sums[5][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[139] [4:0] }), .sum({ \level_1_sums[5][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[5][69] [5:0] }),
     .b({ \level_1_sums[5][68] [5:0] }), .sum({ \level_2_sums[5][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[141] [4:0] }), .sum({ \level_1_sums[5][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[143] [4:0] }), .sum({ \level_1_sums[5][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[5][71] [5:0] }),
     .b({ \level_1_sums[5][70] [5:0] }), .sum({ \level_2_sums[5][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[5][35] [6:0] }),
     .b({ \level_2_sums[5][34] [6:0] }), .sum({ \level_3_sums[5][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[5][17] [7:0] }),
     .b({ \level_3_sums[5][16] [7:0] }), .sum({ \level_4_sums[5][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[145] [4:0] }), .sum({ \level_1_sums[5][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[147] [4:0] }), .sum({ \level_1_sums[5][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[5][73] [5:0] }),
     .b({ \level_1_sums[5][72] [5:0] }), .sum({ \level_2_sums[5][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[149] [4:0] }), .sum({ \level_1_sums[5][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[151] [4:0] }), .sum({ \level_1_sums[5][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[5][75] [5:0] }),
     .b({ \level_1_sums[5][74] [5:0] }), .sum({ \level_2_sums[5][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[5][37] [6:0] }),
     .b({ \level_2_sums[5][36] [6:0] }), .sum({ \level_3_sums[5][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[153] [4:0] }), .sum({ \level_1_sums[5][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[155] [4:0] }), .sum({ \level_1_sums[5][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[5][77] [5:0] }),
     .b({ \level_1_sums[5][76] [5:0] }), .sum({ \level_2_sums[5][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[157] [4:0] }), .sum({ \level_1_sums[5][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[159] [4:0] }), .sum({ \level_1_sums[5][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[5][79] [5:0] }),
     .b({ \level_1_sums[5][78] [5:0] }), .sum({ \level_2_sums[5][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[5][39] [6:0] }),
     .b({ \level_2_sums[5][38] [6:0] }), .sum({ \level_3_sums[5][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[5][19] [7:0] }),
     .b({ \level_3_sums[5][18] [7:0] }), .sum({ \level_4_sums[5][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[5][9] [8:0] }),
     .b({ \level_4_sums[5][8] [8:0] }), .sum({ \level_5_sums[5][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[161] [4:0] }), .sum({ \level_1_sums[5][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[163] [4:0] }), .sum({ \level_1_sums[5][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[5][81] [5:0] }),
     .b({ \level_1_sums[5][80] [5:0] }), .sum({ \level_2_sums[5][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[165] [4:0] }), .sum({ \level_1_sums[5][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[167] [4:0] }), .sum({ \level_1_sums[5][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[5][83] [5:0] }),
     .b({ \level_1_sums[5][82] [5:0] }), .sum({ \level_2_sums[5][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[5][41] [6:0] }),
     .b({ \level_2_sums[5][40] [6:0] }), .sum({ \level_3_sums[5][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[169] [4:0] }), .sum({ \level_1_sums[5][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[171] [4:0] }), .sum({ \level_1_sums[5][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[5][85] [5:0] }),
     .b({ \level_1_sums[5][84] [5:0] }), .sum({ \level_2_sums[5][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[173] [4:0] }), .sum({ \level_1_sums[5][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[175] [4:0] }), .sum({ \level_1_sums[5][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[5][87] [5:0] }),
     .b({ \level_1_sums[5][86] [5:0] }), .sum({ \level_2_sums[5][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[5][43] [6:0] }),
     .b({ \level_2_sums[5][42] [6:0] }), .sum({ \level_3_sums[5][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[5][21] [7:0] }),
     .b({ \level_3_sums[5][20] [7:0] }), .sum({ \level_4_sums[5][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[177] [4:0] }), .sum({ \level_1_sums[5][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[179] [4:0] }), .sum({ \level_1_sums[5][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[5][89] [5:0] }),
     .b({ \level_1_sums[5][88] [5:0] }), .sum({ \level_2_sums[5][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[181] [4:0] }), .sum({ \level_1_sums[5][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[183] [4:0] }), .sum({ \level_1_sums[5][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[5][91] [5:0] }),
     .b({ \level_1_sums[5][90] [5:0] }), .sum({ \level_2_sums[5][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[5][45] [6:0] }),
     .b({ \level_2_sums[5][44] [6:0] }), .sum({ \level_3_sums[5][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[185] [4:0] }), .sum({ \level_1_sums[5][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[187] [4:0] }), .sum({ \level_1_sums[5][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[5][93] [5:0] }),
     .b({ \level_1_sums[5][92] [5:0] }), .sum({ \level_2_sums[5][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[189] [4:0] }), .sum({ \level_1_sums[5][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[191] [4:0] }), .sum({ \level_1_sums[5][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[5][95] [5:0] }),
     .b({ \level_1_sums[5][94] [5:0] }), .sum({ \level_2_sums[5][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[5][47] [6:0] }),
     .b({ \level_2_sums[5][46] [6:0] }), .sum({ \level_3_sums[5][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[5][23] [7:0] }),
     .b({ \level_3_sums[5][22] [7:0] }), .sum({ \level_4_sums[5][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[5][11] [8:0] }),
     .b({ \level_4_sums[5][10] [8:0] }), .sum({ \level_5_sums[5][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[5][5] [9:0] }),
     .b({ \level_5_sums[5][4] [9:0] }), .sum({ \level_6_sums[5][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[193] [4:0] }), .sum({ \level_1_sums[5][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[195] [4:0] }), .sum({ \level_1_sums[5][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[5][97] [5:0] }),
     .b({ \level_1_sums[5][96] [5:0] }), .sum({ \level_2_sums[5][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[197] [4:0] }), .sum({ \level_1_sums[5][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[199] [4:0] }), .sum({ \level_1_sums[5][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[5][99] [5:0] }),
     .b({ \level_1_sums[5][98] [5:0] }), .sum({ \level_2_sums[5][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[5][49] [6:0] }),
     .b({ \level_2_sums[5][48] [6:0] }), .sum({ \level_3_sums[5][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[201] [4:0] }), .sum({ \level_1_sums[5][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[203] [4:0] }), .sum({ \level_1_sums[5][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[5][101] [5:0] }),
     .b({ \level_1_sums[5][100] [5:0] }), .sum({ \level_2_sums[5][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[205] [4:0] }), .sum({ \level_1_sums[5][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[207] [4:0] }), .sum({ \level_1_sums[5][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[5][103] [5:0] }),
     .b({ \level_1_sums[5][102] [5:0] }), .sum({ \level_2_sums[5][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[5][51] [6:0] }),
     .b({ \level_2_sums[5][50] [6:0] }), .sum({ \level_3_sums[5][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[5][25] [7:0] }),
     .b({ \level_3_sums[5][24] [7:0] }), .sum({ \level_4_sums[5][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[209] [4:0] }), .sum({ \level_1_sums[5][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[211] [4:0] }), .sum({ \level_1_sums[5][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[5][105] [5:0] }),
     .b({ \level_1_sums[5][104] [5:0] }), .sum({ \level_2_sums[5][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[213] [4:0] }), .sum({ \level_1_sums[5][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[215] [4:0] }), .sum({ \level_1_sums[5][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[5][107] [5:0] }),
     .b({ \level_1_sums[5][106] [5:0] }), .sum({ \level_2_sums[5][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[5][53] [6:0] }),
     .b({ \level_2_sums[5][52] [6:0] }), .sum({ \level_3_sums[5][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[217] [4:0] }), .sum({ \level_1_sums[5][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[219] [4:0] }), .sum({ \level_1_sums[5][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[5][109] [5:0] }),
     .b({ \level_1_sums[5][108] [5:0] }), .sum({ \level_2_sums[5][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[221] [4:0] }), .sum({ \level_1_sums[5][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[223] [4:0] }), .sum({ \level_1_sums[5][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[5][111] [5:0] }),
     .b({ \level_1_sums[5][110] [5:0] }), .sum({ \level_2_sums[5][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[5][55] [6:0] }),
     .b({ \level_2_sums[5][54] [6:0] }), .sum({ \level_3_sums[5][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[5][27] [7:0] }),
     .b({ \level_3_sums[5][26] [7:0] }), .sum({ \level_4_sums[5][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[5][13] [8:0] }),
     .b({ \level_4_sums[5][12] [8:0] }), .sum({ \level_5_sums[5][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[225] [4:0] }), .sum({ \level_1_sums[5][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[227] [4:0] }), .sum({ \level_1_sums[5][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[5][113] [5:0] }),
     .b({ \level_1_sums[5][112] [5:0] }), .sum({ \level_2_sums[5][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[229] [4:0] }), .sum({ \level_1_sums[5][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[231] [4:0] }), .sum({ \level_1_sums[5][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[5][115] [5:0] }),
     .b({ \level_1_sums[5][114] [5:0] }), .sum({ \level_2_sums[5][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[5][57] [6:0] }),
     .b({ \level_2_sums[5][56] [6:0] }), .sum({ \level_3_sums[5][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[233] [4:0] }), .sum({ \level_1_sums[5][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[235] [4:0] }), .sum({ \level_1_sums[5][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[5][117] [5:0] }),
     .b({ \level_1_sums[5][116] [5:0] }), .sum({ \level_2_sums[5][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[237] [4:0] }), .sum({ \level_1_sums[5][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[239] [4:0] }), .sum({ \level_1_sums[5][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[5][119] [5:0] }),
     .b({ \level_1_sums[5][118] [5:0] }), .sum({ \level_2_sums[5][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[5][59] [6:0] }),
     .b({ \level_2_sums[5][58] [6:0] }), .sum({ \level_3_sums[5][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[5][29] [7:0] }),
     .b({ \level_3_sums[5][28] [7:0] }), .sum({ \level_4_sums[5][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[241] [4:0] }), .sum({ \level_1_sums[5][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[243] [4:0] }), .sum({ \level_1_sums[5][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[5][121] [5:0] }),
     .b({ \level_1_sums[5][120] [5:0] }), .sum({ \level_2_sums[5][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[245] [4:0] }), .sum({ \level_1_sums[5][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[247] [4:0] }), .sum({ \level_1_sums[5][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[5][123] [5:0] }),
     .b({ \level_1_sums[5][122] [5:0] }), .sum({ \level_2_sums[5][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[5][61] [6:0] }),
     .b({ \level_2_sums[5][60] [6:0] }), .sum({ \level_3_sums[5][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[249] [4:0] }), .sum({ \level_1_sums[5][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[251] [4:0] }), .sum({ \level_1_sums[5][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[5][125] [5:0] }),
     .b({ \level_1_sums[5][124] [5:0] }), .sum({ \level_2_sums[5][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[253] [4:0] }), .sum({ \level_1_sums[5][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[5].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[5].product_terms[255] [4:0] }), .sum({ \level_1_sums[5][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[5][127] [5:0] }),
     .b({ \level_1_sums[5][126] [5:0] }), .sum({ \level_2_sums[5][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[5][63] [6:0] }),
     .b({ \level_2_sums[5][62] [6:0] }), .sum({ \level_3_sums[5][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[5][31] [7:0] }),
     .b({ \level_3_sums[5][30] [7:0] }), .sum({ \level_4_sums[5][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[5][15] [8:0] }),
     .b({ \level_4_sums[5][14] [8:0] }), .sum({ \level_5_sums[5][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[5][7] [9:0] }),
     .b({ \level_5_sums[5][6] [9:0] }), .sum({ \level_6_sums[5][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[5][3] [9:0] }),
     .b({ \level_6_sums[5][2] [9:0] }), .sum({ \level_7_sums[5][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[5].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[5][0] [9:0] }),
     .b({ \level_7_sums[5][1] [9:0] }), .sum({ \level_8_sums[5] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[6].relu_inst (.in_data({ \final_sums[6] [9:0] }), .out_data({ \out_sig[6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[1] [4:0] }), .sum({ \level_1_sums[6][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[3] [4:0] }), .sum({ \level_1_sums[6][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[6][1] [5:0] }),
     .b({ \level_1_sums[6][0] [5:0] }), .sum({ \level_2_sums[6][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[5] [4:0] }), .sum({ \level_1_sums[6][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[7] [4:0] }), .sum({ \level_1_sums[6][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[6][3] [5:0] }),
     .b({ \level_1_sums[6][2] [5:0] }), .sum({ \level_2_sums[6][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[6][1] [6:0] }),
     .b({ \level_2_sums[6][0] [6:0] }), .sum({ \level_3_sums[6][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[9] [4:0] }), .sum({ \level_1_sums[6][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[11] [4:0] }), .sum({ \level_1_sums[6][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[6][5] [5:0] }),
     .b({ \level_1_sums[6][4] [5:0] }), .sum({ \level_2_sums[6][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[13] [4:0] }), .sum({ \level_1_sums[6][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[15] [4:0] }), .sum({ \level_1_sums[6][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[6][7] [5:0] }),
     .b({ \level_1_sums[6][6] [5:0] }), .sum({ \level_2_sums[6][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[6][3] [6:0] }),
     .b({ \level_2_sums[6][2] [6:0] }), .sum({ \level_3_sums[6][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[6][1] [7:0] }),
     .b({ \level_3_sums[6][0] [7:0] }), .sum({ \level_4_sums[6][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[17] [4:0] }), .sum({ \level_1_sums[6][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[19] [4:0] }), .sum({ \level_1_sums[6][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[6][9] [5:0] }),
     .b({ \level_1_sums[6][8] [5:0] }), .sum({ \level_2_sums[6][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[21] [4:0] }), .sum({ \level_1_sums[6][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[23] [4:0] }), .sum({ \level_1_sums[6][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[6][11] [5:0] }),
     .b({ \level_1_sums[6][10] [5:0] }), .sum({ \level_2_sums[6][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[6][5] [6:0] }),
     .b({ \level_2_sums[6][4] [6:0] }), .sum({ \level_3_sums[6][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[25] [4:0] }), .sum({ \level_1_sums[6][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[27] [4:0] }), .sum({ \level_1_sums[6][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[6][13] [5:0] }),
     .b({ \level_1_sums[6][12] [5:0] }), .sum({ \level_2_sums[6][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[29] [4:0] }), .sum({ \level_1_sums[6][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[31] [4:0] }), .sum({ \level_1_sums[6][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[6][15] [5:0] }),
     .b({ \level_1_sums[6][14] [5:0] }), .sum({ \level_2_sums[6][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[6][7] [6:0] }),
     .b({ \level_2_sums[6][6] [6:0] }), .sum({ \level_3_sums[6][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[6][3] [7:0] }),
     .b({ \level_3_sums[6][2] [7:0] }), .sum({ \level_4_sums[6][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[6][1] [8:0] }),
     .b({ \level_4_sums[6][0] [8:0] }), .sum({ \level_5_sums[6][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[33] [4:0] }), .sum({ \level_1_sums[6][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[35] [4:0] }), .sum({ \level_1_sums[6][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[6][17] [5:0] }),
     .b({ \level_1_sums[6][16] [5:0] }), .sum({ \level_2_sums[6][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[37] [4:0] }), .sum({ \level_1_sums[6][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[39] [4:0] }), .sum({ \level_1_sums[6][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[6][19] [5:0] }),
     .b({ \level_1_sums[6][18] [5:0] }), .sum({ \level_2_sums[6][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[6][9] [6:0] }),
     .b({ \level_2_sums[6][8] [6:0] }), .sum({ \level_3_sums[6][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[41] [4:0] }), .sum({ \level_1_sums[6][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[43] [4:0] }), .sum({ \level_1_sums[6][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[6][21] [5:0] }),
     .b({ \level_1_sums[6][20] [5:0] }), .sum({ \level_2_sums[6][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[45] [4:0] }), .sum({ \level_1_sums[6][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[47] [4:0] }), .sum({ \level_1_sums[6][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[6][23] [5:0] }),
     .b({ \level_1_sums[6][22] [5:0] }), .sum({ \level_2_sums[6][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[6][11] [6:0] }),
     .b({ \level_2_sums[6][10] [6:0] }), .sum({ \level_3_sums[6][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[6][5] [7:0] }),
     .b({ \level_3_sums[6][4] [7:0] }), .sum({ \level_4_sums[6][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[49] [4:0] }), .sum({ \level_1_sums[6][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[51] [4:0] }), .sum({ \level_1_sums[6][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[6][25] [5:0] }),
     .b({ \level_1_sums[6][24] [5:0] }), .sum({ \level_2_sums[6][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[53] [4:0] }), .sum({ \level_1_sums[6][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[55] [4:0] }), .sum({ \level_1_sums[6][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[6][27] [5:0] }),
     .b({ \level_1_sums[6][26] [5:0] }), .sum({ \level_2_sums[6][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[6][13] [6:0] }),
     .b({ \level_2_sums[6][12] [6:0] }), .sum({ \level_3_sums[6][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[57] [4:0] }), .sum({ \level_1_sums[6][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[59] [4:0] }), .sum({ \level_1_sums[6][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[6][29] [5:0] }),
     .b({ \level_1_sums[6][28] [5:0] }), .sum({ \level_2_sums[6][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[61] [4:0] }), .sum({ \level_1_sums[6][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[63] [4:0] }), .sum({ \level_1_sums[6][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[6][31] [5:0] }),
     .b({ \level_1_sums[6][30] [5:0] }), .sum({ \level_2_sums[6][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[6][15] [6:0] }),
     .b({ \level_2_sums[6][14] [6:0] }), .sum({ \level_3_sums[6][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[6][7] [7:0] }),
     .b({ \level_3_sums[6][6] [7:0] }), .sum({ \level_4_sums[6][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[6][3] [8:0] }),
     .b({ \level_4_sums[6][2] [8:0] }), .sum({ \level_5_sums[6][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[6][1] [9:0] }),
     .b({ \level_5_sums[6][0] [9:0] }), .sum({ \level_6_sums[6][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[65] [4:0] }), .sum({ \level_1_sums[6][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[67] [4:0] }), .sum({ \level_1_sums[6][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[6][33] [5:0] }),
     .b({ \level_1_sums[6][32] [5:0] }), .sum({ \level_2_sums[6][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[69] [4:0] }), .sum({ \level_1_sums[6][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[71] [4:0] }), .sum({ \level_1_sums[6][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[6][35] [5:0] }),
     .b({ \level_1_sums[6][34] [5:0] }), .sum({ \level_2_sums[6][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[6][17] [6:0] }),
     .b({ \level_2_sums[6][16] [6:0] }), .sum({ \level_3_sums[6][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[73] [4:0] }), .sum({ \level_1_sums[6][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[75] [4:0] }), .sum({ \level_1_sums[6][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[6][37] [5:0] }),
     .b({ \level_1_sums[6][36] [5:0] }), .sum({ \level_2_sums[6][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[77] [4:0] }), .sum({ \level_1_sums[6][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[79] [4:0] }), .sum({ \level_1_sums[6][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[6][39] [5:0] }),
     .b({ \level_1_sums[6][38] [5:0] }), .sum({ \level_2_sums[6][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[6][19] [6:0] }),
     .b({ \level_2_sums[6][18] [6:0] }), .sum({ \level_3_sums[6][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[6][9] [7:0] }),
     .b({ \level_3_sums[6][8] [7:0] }), .sum({ \level_4_sums[6][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[81] [4:0] }), .sum({ \level_1_sums[6][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[83] [4:0] }), .sum({ \level_1_sums[6][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[6][41] [5:0] }),
     .b({ \level_1_sums[6][40] [5:0] }), .sum({ \level_2_sums[6][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[85] [4:0] }), .sum({ \level_1_sums[6][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[87] [4:0] }), .sum({ \level_1_sums[6][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[6][43] [5:0] }),
     .b({ \level_1_sums[6][42] [5:0] }), .sum({ \level_2_sums[6][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[6][21] [6:0] }),
     .b({ \level_2_sums[6][20] [6:0] }), .sum({ \level_3_sums[6][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[89] [4:0] }), .sum({ \level_1_sums[6][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[91] [4:0] }), .sum({ \level_1_sums[6][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[6][45] [5:0] }),
     .b({ \level_1_sums[6][44] [5:0] }), .sum({ \level_2_sums[6][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[93] [4:0] }), .sum({ \level_1_sums[6][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[95] [4:0] }), .sum({ \level_1_sums[6][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[6][47] [5:0] }),
     .b({ \level_1_sums[6][46] [5:0] }), .sum({ \level_2_sums[6][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[6][23] [6:0] }),
     .b({ \level_2_sums[6][22] [6:0] }), .sum({ \level_3_sums[6][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[6][11] [7:0] }),
     .b({ \level_3_sums[6][10] [7:0] }), .sum({ \level_4_sums[6][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[6][5] [8:0] }),
     .b({ \level_4_sums[6][4] [8:0] }), .sum({ \level_5_sums[6][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[97] [4:0] }), .sum({ \level_1_sums[6][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[99] [4:0] }), .sum({ \level_1_sums[6][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[6][49] [5:0] }),
     .b({ \level_1_sums[6][48] [5:0] }), .sum({ \level_2_sums[6][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[101] [4:0] }), .sum({ \level_1_sums[6][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[103] [4:0] }), .sum({ \level_1_sums[6][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[6][51] [5:0] }),
     .b({ \level_1_sums[6][50] [5:0] }), .sum({ \level_2_sums[6][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[6][25] [6:0] }),
     .b({ \level_2_sums[6][24] [6:0] }), .sum({ \level_3_sums[6][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[105] [4:0] }), .sum({ \level_1_sums[6][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[107] [4:0] }), .sum({ \level_1_sums[6][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[6][53] [5:0] }),
     .b({ \level_1_sums[6][52] [5:0] }), .sum({ \level_2_sums[6][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[109] [4:0] }), .sum({ \level_1_sums[6][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[111] [4:0] }), .sum({ \level_1_sums[6][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[6][55] [5:0] }),
     .b({ \level_1_sums[6][54] [5:0] }), .sum({ \level_2_sums[6][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[6][27] [6:0] }),
     .b({ \level_2_sums[6][26] [6:0] }), .sum({ \level_3_sums[6][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[6][13] [7:0] }),
     .b({ \level_3_sums[6][12] [7:0] }), .sum({ \level_4_sums[6][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[113] [4:0] }), .sum({ \level_1_sums[6][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[115] [4:0] }), .sum({ \level_1_sums[6][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[6][57] [5:0] }),
     .b({ \level_1_sums[6][56] [5:0] }), .sum({ \level_2_sums[6][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[117] [4:0] }), .sum({ \level_1_sums[6][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[119] [4:0] }), .sum({ \level_1_sums[6][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[6][59] [5:0] }),
     .b({ \level_1_sums[6][58] [5:0] }), .sum({ \level_2_sums[6][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[6][29] [6:0] }),
     .b({ \level_2_sums[6][28] [6:0] }), .sum({ \level_3_sums[6][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[121] [4:0] }), .sum({ \level_1_sums[6][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[123] [4:0] }), .sum({ \level_1_sums[6][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[6][61] [5:0] }),
     .b({ \level_1_sums[6][60] [5:0] }), .sum({ \level_2_sums[6][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[125] [4:0] }), .sum({ \level_1_sums[6][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[127] [4:0] }), .sum({ \level_1_sums[6][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[6][63] [5:0] }),
     .b({ \level_1_sums[6][62] [5:0] }), .sum({ \level_2_sums[6][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[6][31] [6:0] }),
     .b({ \level_2_sums[6][30] [6:0] }), .sum({ \level_3_sums[6][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[6][15] [7:0] }),
     .b({ \level_3_sums[6][14] [7:0] }), .sum({ \level_4_sums[6][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[6][7] [8:0] }),
     .b({ \level_4_sums[6][6] [8:0] }), .sum({ \level_5_sums[6][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[6][3] [9:0] }),
     .b({ \level_5_sums[6][2] [9:0] }), .sum({ \level_6_sums[6][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[6][1] [9:0] }),
     .b({ \level_6_sums[6][0] [9:0] }), .sum({ \level_7_sums[6][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[129] [4:0] }), .sum({ \level_1_sums[6][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[131] [4:0] }), .sum({ \level_1_sums[6][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[6][65] [5:0] }),
     .b({ \level_1_sums[6][64] [5:0] }), .sum({ \level_2_sums[6][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[133] [4:0] }), .sum({ \level_1_sums[6][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[135] [4:0] }), .sum({ \level_1_sums[6][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[6][67] [5:0] }),
     .b({ \level_1_sums[6][66] [5:0] }), .sum({ \level_2_sums[6][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[6][33] [6:0] }),
     .b({ \level_2_sums[6][32] [6:0] }), .sum({ \level_3_sums[6][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[137] [4:0] }), .sum({ \level_1_sums[6][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[139] [4:0] }), .sum({ \level_1_sums[6][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[6][69] [5:0] }),
     .b({ \level_1_sums[6][68] [5:0] }), .sum({ \level_2_sums[6][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[141] [4:0] }), .sum({ \level_1_sums[6][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[143] [4:0] }), .sum({ \level_1_sums[6][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[6][71] [5:0] }),
     .b({ \level_1_sums[6][70] [5:0] }), .sum({ \level_2_sums[6][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[6][35] [6:0] }),
     .b({ \level_2_sums[6][34] [6:0] }), .sum({ \level_3_sums[6][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[6][17] [7:0] }),
     .b({ \level_3_sums[6][16] [7:0] }), .sum({ \level_4_sums[6][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[145] [4:0] }), .sum({ \level_1_sums[6][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[147] [4:0] }), .sum({ \level_1_sums[6][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[6][73] [5:0] }),
     .b({ \level_1_sums[6][72] [5:0] }), .sum({ \level_2_sums[6][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[149] [4:0] }), .sum({ \level_1_sums[6][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[151] [4:0] }), .sum({ \level_1_sums[6][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[6][75] [5:0] }),
     .b({ \level_1_sums[6][74] [5:0] }), .sum({ \level_2_sums[6][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[6][37] [6:0] }),
     .b({ \level_2_sums[6][36] [6:0] }), .sum({ \level_3_sums[6][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[153] [4:0] }), .sum({ \level_1_sums[6][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[155] [4:0] }), .sum({ \level_1_sums[6][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[6][77] [5:0] }),
     .b({ \level_1_sums[6][76] [5:0] }), .sum({ \level_2_sums[6][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[157] [4:0] }), .sum({ \level_1_sums[6][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[159] [4:0] }), .sum({ \level_1_sums[6][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[6][79] [5:0] }),
     .b({ \level_1_sums[6][78] [5:0] }), .sum({ \level_2_sums[6][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[6][39] [6:0] }),
     .b({ \level_2_sums[6][38] [6:0] }), .sum({ \level_3_sums[6][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[6][19] [7:0] }),
     .b({ \level_3_sums[6][18] [7:0] }), .sum({ \level_4_sums[6][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[6][9] [8:0] }),
     .b({ \level_4_sums[6][8] [8:0] }), .sum({ \level_5_sums[6][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[161] [4:0] }), .sum({ \level_1_sums[6][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[163] [4:0] }), .sum({ \level_1_sums[6][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[6][81] [5:0] }),
     .b({ \level_1_sums[6][80] [5:0] }), .sum({ \level_2_sums[6][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[165] [4:0] }), .sum({ \level_1_sums[6][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[167] [4:0] }), .sum({ \level_1_sums[6][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[6][83] [5:0] }),
     .b({ \level_1_sums[6][82] [5:0] }), .sum({ \level_2_sums[6][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[6][41] [6:0] }),
     .b({ \level_2_sums[6][40] [6:0] }), .sum({ \level_3_sums[6][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[169] [4:0] }), .sum({ \level_1_sums[6][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[171] [4:0] }), .sum({ \level_1_sums[6][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[6][85] [5:0] }),
     .b({ \level_1_sums[6][84] [5:0] }), .sum({ \level_2_sums[6][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[173] [4:0] }), .sum({ \level_1_sums[6][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[175] [4:0] }), .sum({ \level_1_sums[6][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[6][87] [5:0] }),
     .b({ \level_1_sums[6][86] [5:0] }), .sum({ \level_2_sums[6][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[6][43] [6:0] }),
     .b({ \level_2_sums[6][42] [6:0] }), .sum({ \level_3_sums[6][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[6][21] [7:0] }),
     .b({ \level_3_sums[6][20] [7:0] }), .sum({ \level_4_sums[6][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[177] [4:0] }), .sum({ \level_1_sums[6][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[179] [4:0] }), .sum({ \level_1_sums[6][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[6][89] [5:0] }),
     .b({ \level_1_sums[6][88] [5:0] }), .sum({ \level_2_sums[6][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[181] [4:0] }), .sum({ \level_1_sums[6][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[183] [4:0] }), .sum({ \level_1_sums[6][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[6][91] [5:0] }),
     .b({ \level_1_sums[6][90] [5:0] }), .sum({ \level_2_sums[6][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[6][45] [6:0] }),
     .b({ \level_2_sums[6][44] [6:0] }), .sum({ \level_3_sums[6][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[185] [4:0] }), .sum({ \level_1_sums[6][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[187] [4:0] }), .sum({ \level_1_sums[6][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[6][93] [5:0] }),
     .b({ \level_1_sums[6][92] [5:0] }), .sum({ \level_2_sums[6][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[189] [4:0] }), .sum({ \level_1_sums[6][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[191] [4:0] }), .sum({ \level_1_sums[6][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[6][95] [5:0] }),
     .b({ \level_1_sums[6][94] [5:0] }), .sum({ \level_2_sums[6][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[6][47] [6:0] }),
     .b({ \level_2_sums[6][46] [6:0] }), .sum({ \level_3_sums[6][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[6][23] [7:0] }),
     .b({ \level_3_sums[6][22] [7:0] }), .sum({ \level_4_sums[6][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[6][11] [8:0] }),
     .b({ \level_4_sums[6][10] [8:0] }), .sum({ \level_5_sums[6][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[6][5] [9:0] }),
     .b({ \level_5_sums[6][4] [9:0] }), .sum({ \level_6_sums[6][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[193] [4:0] }), .sum({ \level_1_sums[6][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[195] [4:0] }), .sum({ \level_1_sums[6][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[6][97] [5:0] }),
     .b({ \level_1_sums[6][96] [5:0] }), .sum({ \level_2_sums[6][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[197] [4:0] }), .sum({ \level_1_sums[6][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[199] [4:0] }), .sum({ \level_1_sums[6][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[6][99] [5:0] }),
     .b({ \level_1_sums[6][98] [5:0] }), .sum({ \level_2_sums[6][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[6][49] [6:0] }),
     .b({ \level_2_sums[6][48] [6:0] }), .sum({ \level_3_sums[6][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[201] [4:0] }), .sum({ \level_1_sums[6][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[203] [4:0] }), .sum({ \level_1_sums[6][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[6][101] [5:0] }),
     .b({ \level_1_sums[6][100] [5:0] }), .sum({ \level_2_sums[6][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[205] [4:0] }), .sum({ \level_1_sums[6][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[207] [4:0] }), .sum({ \level_1_sums[6][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[6][103] [5:0] }),
     .b({ \level_1_sums[6][102] [5:0] }), .sum({ \level_2_sums[6][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[6][51] [6:0] }),
     .b({ \level_2_sums[6][50] [6:0] }), .sum({ \level_3_sums[6][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[6][25] [7:0] }),
     .b({ \level_3_sums[6][24] [7:0] }), .sum({ \level_4_sums[6][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[209] [4:0] }), .sum({ \level_1_sums[6][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[211] [4:0] }), .sum({ \level_1_sums[6][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[6][105] [5:0] }),
     .b({ \level_1_sums[6][104] [5:0] }), .sum({ \level_2_sums[6][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[213] [4:0] }), .sum({ \level_1_sums[6][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[215] [4:0] }), .sum({ \level_1_sums[6][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[6][107] [5:0] }),
     .b({ \level_1_sums[6][106] [5:0] }), .sum({ \level_2_sums[6][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[6][53] [6:0] }),
     .b({ \level_2_sums[6][52] [6:0] }), .sum({ \level_3_sums[6][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[217] [4:0] }), .sum({ \level_1_sums[6][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[219] [4:0] }), .sum({ \level_1_sums[6][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[6][109] [5:0] }),
     .b({ \level_1_sums[6][108] [5:0] }), .sum({ \level_2_sums[6][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[221] [4:0] }), .sum({ \level_1_sums[6][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[223] [4:0] }), .sum({ \level_1_sums[6][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[6][111] [5:0] }),
     .b({ \level_1_sums[6][110] [5:0] }), .sum({ \level_2_sums[6][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[6][55] [6:0] }),
     .b({ \level_2_sums[6][54] [6:0] }), .sum({ \level_3_sums[6][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[6][27] [7:0] }),
     .b({ \level_3_sums[6][26] [7:0] }), .sum({ \level_4_sums[6][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[6][13] [8:0] }),
     .b({ \level_4_sums[6][12] [8:0] }), .sum({ \level_5_sums[6][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[225] [4:0] }), .sum({ \level_1_sums[6][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[227] [4:0] }), .sum({ \level_1_sums[6][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[6][113] [5:0] }),
     .b({ \level_1_sums[6][112] [5:0] }), .sum({ \level_2_sums[6][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[229] [4:0] }), .sum({ \level_1_sums[6][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[231] [4:0] }), .sum({ \level_1_sums[6][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[6][115] [5:0] }),
     .b({ \level_1_sums[6][114] [5:0] }), .sum({ \level_2_sums[6][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[6][57] [6:0] }),
     .b({ \level_2_sums[6][56] [6:0] }), .sum({ \level_3_sums[6][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[233] [4:0] }), .sum({ \level_1_sums[6][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[235] [4:0] }), .sum({ \level_1_sums[6][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[6][117] [5:0] }),
     .b({ \level_1_sums[6][116] [5:0] }), .sum({ \level_2_sums[6][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[237] [4:0] }), .sum({ \level_1_sums[6][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[239] [4:0] }), .sum({ \level_1_sums[6][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[6][119] [5:0] }),
     .b({ \level_1_sums[6][118] [5:0] }), .sum({ \level_2_sums[6][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[6][59] [6:0] }),
     .b({ \level_2_sums[6][58] [6:0] }), .sum({ \level_3_sums[6][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[6][29] [7:0] }),
     .b({ \level_3_sums[6][28] [7:0] }), .sum({ \level_4_sums[6][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[241] [4:0] }), .sum({ \level_1_sums[6][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[243] [4:0] }), .sum({ \level_1_sums[6][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[6][121] [5:0] }),
     .b({ \level_1_sums[6][120] [5:0] }), .sum({ \level_2_sums[6][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[245] [4:0] }), .sum({ \level_1_sums[6][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[247] [4:0] }), .sum({ \level_1_sums[6][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[6][123] [5:0] }),
     .b({ \level_1_sums[6][122] [5:0] }), .sum({ \level_2_sums[6][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[6][61] [6:0] }),
     .b({ \level_2_sums[6][60] [6:0] }), .sum({ \level_3_sums[6][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[249] [4:0] }), .sum({ \level_1_sums[6][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[251] [4:0] }), .sum({ \level_1_sums[6][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[6][125] [5:0] }),
     .b({ \level_1_sums[6][124] [5:0] }), .sum({ \level_2_sums[6][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[253] [4:0] }), .sum({ \level_1_sums[6][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[6].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[6].product_terms[255] [4:0] }), .sum({ \level_1_sums[6][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[6][127] [5:0] }),
     .b({ \level_1_sums[6][126] [5:0] }), .sum({ \level_2_sums[6][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[6][63] [6:0] }),
     .b({ \level_2_sums[6][62] [6:0] }), .sum({ \level_3_sums[6][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[6][31] [7:0] }),
     .b({ \level_3_sums[6][30] [7:0] }), .sum({ \level_4_sums[6][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[6][15] [8:0] }),
     .b({ \level_4_sums[6][14] [8:0] }), .sum({ \level_5_sums[6][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[6][7] [9:0] }),
     .b({ \level_5_sums[6][6] [9:0] }), .sum({ \level_6_sums[6][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[6][3] [9:0] }),
     .b({ \level_6_sums[6][2] [9:0] }), .sum({ \level_7_sums[6][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[6].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[6][0] [9:0] }),
     .b({ \level_7_sums[6][1] [9:0] }), .sum({ \level_8_sums[6] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[7].relu_inst (.in_data({ \final_sums[7] [9:0] }), .out_data({ \out_sig[7] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[1] [4:0] }), .sum({ \level_1_sums[7][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[3] [4:0] }), .sum({ \level_1_sums[7][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[7][1] [5:0] }),
     .b({ \level_1_sums[7][0] [5:0] }), .sum({ \level_2_sums[7][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[5] [4:0] }), .sum({ \level_1_sums[7][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[7] [4:0] }), .sum({ \level_1_sums[7][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[7][3] [5:0] }),
     .b({ \level_1_sums[7][2] [5:0] }), .sum({ \level_2_sums[7][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[7][1] [6:0] }),
     .b({ \level_2_sums[7][0] [6:0] }), .sum({ \level_3_sums[7][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[9] [4:0] }), .sum({ \level_1_sums[7][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[11] [4:0] }), .sum({ \level_1_sums[7][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[7][5] [5:0] }),
     .b({ \level_1_sums[7][4] [5:0] }), .sum({ \level_2_sums[7][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[13] [4:0] }), .sum({ \level_1_sums[7][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[15] [4:0] }), .sum({ \level_1_sums[7][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[7][7] [5:0] }),
     .b({ \level_1_sums[7][6] [5:0] }), .sum({ \level_2_sums[7][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[7][3] [6:0] }),
     .b({ \level_2_sums[7][2] [6:0] }), .sum({ \level_3_sums[7][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[7][1] [7:0] }),
     .b({ \level_3_sums[7][0] [7:0] }), .sum({ \level_4_sums[7][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[17] [4:0] }), .sum({ \level_1_sums[7][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[19] [4:0] }), .sum({ \level_1_sums[7][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[7][9] [5:0] }),
     .b({ \level_1_sums[7][8] [5:0] }), .sum({ \level_2_sums[7][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[21] [4:0] }), .sum({ \level_1_sums[7][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[23] [4:0] }), .sum({ \level_1_sums[7][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[7][11] [5:0] }),
     .b({ \level_1_sums[7][10] [5:0] }), .sum({ \level_2_sums[7][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[7][5] [6:0] }),
     .b({ \level_2_sums[7][4] [6:0] }), .sum({ \level_3_sums[7][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[25] [4:0] }), .sum({ \level_1_sums[7][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[27] [4:0] }), .sum({ \level_1_sums[7][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[7][13] [5:0] }),
     .b({ \level_1_sums[7][12] [5:0] }), .sum({ \level_2_sums[7][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[29] [4:0] }), .sum({ \level_1_sums[7][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[31] [4:0] }), .sum({ \level_1_sums[7][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[7][15] [5:0] }),
     .b({ \level_1_sums[7][14] [5:0] }), .sum({ \level_2_sums[7][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[7][7] [6:0] }),
     .b({ \level_2_sums[7][6] [6:0] }), .sum({ \level_3_sums[7][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[7][3] [7:0] }),
     .b({ \level_3_sums[7][2] [7:0] }), .sum({ \level_4_sums[7][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[7][1] [8:0] }),
     .b({ \level_4_sums[7][0] [8:0] }), .sum({ \level_5_sums[7][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[33] [4:0] }), .sum({ \level_1_sums[7][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[35] [4:0] }), .sum({ \level_1_sums[7][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[7][17] [5:0] }),
     .b({ \level_1_sums[7][16] [5:0] }), .sum({ \level_2_sums[7][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[37] [4:0] }), .sum({ \level_1_sums[7][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[39] [4:0] }), .sum({ \level_1_sums[7][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[7][19] [5:0] }),
     .b({ \level_1_sums[7][18] [5:0] }), .sum({ \level_2_sums[7][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[7][9] [6:0] }),
     .b({ \level_2_sums[7][8] [6:0] }), .sum({ \level_3_sums[7][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[41] [4:0] }), .sum({ \level_1_sums[7][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[43] [4:0] }), .sum({ \level_1_sums[7][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[7][21] [5:0] }),
     .b({ \level_1_sums[7][20] [5:0] }), .sum({ \level_2_sums[7][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[45] [4:0] }), .sum({ \level_1_sums[7][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[47] [4:0] }), .sum({ \level_1_sums[7][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[7][23] [5:0] }),
     .b({ \level_1_sums[7][22] [5:0] }), .sum({ \level_2_sums[7][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[7][11] [6:0] }),
     .b({ \level_2_sums[7][10] [6:0] }), .sum({ \level_3_sums[7][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[7][5] [7:0] }),
     .b({ \level_3_sums[7][4] [7:0] }), .sum({ \level_4_sums[7][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[49] [4:0] }), .sum({ \level_1_sums[7][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[51] [4:0] }), .sum({ \level_1_sums[7][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[7][25] [5:0] }),
     .b({ \level_1_sums[7][24] [5:0] }), .sum({ \level_2_sums[7][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[53] [4:0] }), .sum({ \level_1_sums[7][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[55] [4:0] }), .sum({ \level_1_sums[7][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[7][27] [5:0] }),
     .b({ \level_1_sums[7][26] [5:0] }), .sum({ \level_2_sums[7][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[7][13] [6:0] }),
     .b({ \level_2_sums[7][12] [6:0] }), .sum({ \level_3_sums[7][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[57] [4:0] }), .sum({ \level_1_sums[7][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[59] [4:0] }), .sum({ \level_1_sums[7][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[7][29] [5:0] }),
     .b({ \level_1_sums[7][28] [5:0] }), .sum({ \level_2_sums[7][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[61] [4:0] }), .sum({ \level_1_sums[7][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[63] [4:0] }), .sum({ \level_1_sums[7][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[7][31] [5:0] }),
     .b({ \level_1_sums[7][30] [5:0] }), .sum({ \level_2_sums[7][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[7][15] [6:0] }),
     .b({ \level_2_sums[7][14] [6:0] }), .sum({ \level_3_sums[7][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[7][7] [7:0] }),
     .b({ \level_3_sums[7][6] [7:0] }), .sum({ \level_4_sums[7][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[7][3] [8:0] }),
     .b({ \level_4_sums[7][2] [8:0] }), .sum({ \level_5_sums[7][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[7][1] [9:0] }),
     .b({ \level_5_sums[7][0] [9:0] }), .sum({ \level_6_sums[7][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[65] [4:0] }), .sum({ \level_1_sums[7][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[67] [4:0] }), .sum({ \level_1_sums[7][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[7][33] [5:0] }),
     .b({ \level_1_sums[7][32] [5:0] }), .sum({ \level_2_sums[7][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[69] [4:0] }), .sum({ \level_1_sums[7][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[71] [4:0] }), .sum({ \level_1_sums[7][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[7][35] [5:0] }),
     .b({ \level_1_sums[7][34] [5:0] }), .sum({ \level_2_sums[7][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[7][17] [6:0] }),
     .b({ \level_2_sums[7][16] [6:0] }), .sum({ \level_3_sums[7][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[73] [4:0] }), .sum({ \level_1_sums[7][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[75] [4:0] }), .sum({ \level_1_sums[7][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[7][37] [5:0] }),
     .b({ \level_1_sums[7][36] [5:0] }), .sum({ \level_2_sums[7][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[77] [4:0] }), .sum({ \level_1_sums[7][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[79] [4:0] }), .sum({ \level_1_sums[7][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[7][39] [5:0] }),
     .b({ \level_1_sums[7][38] [5:0] }), .sum({ \level_2_sums[7][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[7][19] [6:0] }),
     .b({ \level_2_sums[7][18] [6:0] }), .sum({ \level_3_sums[7][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[7][9] [7:0] }),
     .b({ \level_3_sums[7][8] [7:0] }), .sum({ \level_4_sums[7][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[81] [4:0] }), .sum({ \level_1_sums[7][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[83] [4:0] }), .sum({ \level_1_sums[7][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[7][41] [5:0] }),
     .b({ \level_1_sums[7][40] [5:0] }), .sum({ \level_2_sums[7][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[85] [4:0] }), .sum({ \level_1_sums[7][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[87] [4:0] }), .sum({ \level_1_sums[7][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[7][43] [5:0] }),
     .b({ \level_1_sums[7][42] [5:0] }), .sum({ \level_2_sums[7][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[7][21] [6:0] }),
     .b({ \level_2_sums[7][20] [6:0] }), .sum({ \level_3_sums[7][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[89] [4:0] }), .sum({ \level_1_sums[7][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[91] [4:0] }), .sum({ \level_1_sums[7][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[7][45] [5:0] }),
     .b({ \level_1_sums[7][44] [5:0] }), .sum({ \level_2_sums[7][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[93] [4:0] }), .sum({ \level_1_sums[7][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[95] [4:0] }), .sum({ \level_1_sums[7][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[7][47] [5:0] }),
     .b({ \level_1_sums[7][46] [5:0] }), .sum({ \level_2_sums[7][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[7][23] [6:0] }),
     .b({ \level_2_sums[7][22] [6:0] }), .sum({ \level_3_sums[7][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[7][11] [7:0] }),
     .b({ \level_3_sums[7][10] [7:0] }), .sum({ \level_4_sums[7][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[7][5] [8:0] }),
     .b({ \level_4_sums[7][4] [8:0] }), .sum({ \level_5_sums[7][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[97] [4:0] }), .sum({ \level_1_sums[7][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[99] [4:0] }), .sum({ \level_1_sums[7][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[7][49] [5:0] }),
     .b({ \level_1_sums[7][48] [5:0] }), .sum({ \level_2_sums[7][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[101] [4:0] }), .sum({ \level_1_sums[7][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[103] [4:0] }), .sum({ \level_1_sums[7][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[7][51] [5:0] }),
     .b({ \level_1_sums[7][50] [5:0] }), .sum({ \level_2_sums[7][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[7][25] [6:0] }),
     .b({ \level_2_sums[7][24] [6:0] }), .sum({ \level_3_sums[7][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[105] [4:0] }), .sum({ \level_1_sums[7][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[107] [4:0] }), .sum({ \level_1_sums[7][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[7][53] [5:0] }),
     .b({ \level_1_sums[7][52] [5:0] }), .sum({ \level_2_sums[7][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[109] [4:0] }), .sum({ \level_1_sums[7][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[111] [4:0] }), .sum({ \level_1_sums[7][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[7][55] [5:0] }),
     .b({ \level_1_sums[7][54] [5:0] }), .sum({ \level_2_sums[7][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[7][27] [6:0] }),
     .b({ \level_2_sums[7][26] [6:0] }), .sum({ \level_3_sums[7][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[7][13] [7:0] }),
     .b({ \level_3_sums[7][12] [7:0] }), .sum({ \level_4_sums[7][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[113] [4:0] }), .sum({ \level_1_sums[7][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[115] [4:0] }), .sum({ \level_1_sums[7][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[7][57] [5:0] }),
     .b({ \level_1_sums[7][56] [5:0] }), .sum({ \level_2_sums[7][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[117] [4:0] }), .sum({ \level_1_sums[7][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[119] [4:0] }), .sum({ \level_1_sums[7][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[7][59] [5:0] }),
     .b({ \level_1_sums[7][58] [5:0] }), .sum({ \level_2_sums[7][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[7][29] [6:0] }),
     .b({ \level_2_sums[7][28] [6:0] }), .sum({ \level_3_sums[7][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[121] [4:0] }), .sum({ \level_1_sums[7][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[123] [4:0] }), .sum({ \level_1_sums[7][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[7][61] [5:0] }),
     .b({ \level_1_sums[7][60] [5:0] }), .sum({ \level_2_sums[7][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[125] [4:0] }), .sum({ \level_1_sums[7][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[127] [4:0] }), .sum({ \level_1_sums[7][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[7][63] [5:0] }),
     .b({ \level_1_sums[7][62] [5:0] }), .sum({ \level_2_sums[7][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[7][31] [6:0] }),
     .b({ \level_2_sums[7][30] [6:0] }), .sum({ \level_3_sums[7][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[7][15] [7:0] }),
     .b({ \level_3_sums[7][14] [7:0] }), .sum({ \level_4_sums[7][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[7][7] [8:0] }),
     .b({ \level_4_sums[7][6] [8:0] }), .sum({ \level_5_sums[7][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[7][3] [9:0] }),
     .b({ \level_5_sums[7][2] [9:0] }), .sum({ \level_6_sums[7][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[7][1] [9:0] }),
     .b({ \level_6_sums[7][0] [9:0] }), .sum({ \level_7_sums[7][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[129] [4:0] }), .sum({ \level_1_sums[7][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[131] [4:0] }), .sum({ \level_1_sums[7][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[7][65] [5:0] }),
     .b({ \level_1_sums[7][64] [5:0] }), .sum({ \level_2_sums[7][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[133] [4:0] }), .sum({ \level_1_sums[7][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[135] [4:0] }), .sum({ \level_1_sums[7][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[7][67] [5:0] }),
     .b({ \level_1_sums[7][66] [5:0] }), .sum({ \level_2_sums[7][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[7][33] [6:0] }),
     .b({ \level_2_sums[7][32] [6:0] }), .sum({ \level_3_sums[7][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[137] [4:0] }), .sum({ \level_1_sums[7][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[139] [4:0] }), .sum({ \level_1_sums[7][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[7][69] [5:0] }),
     .b({ \level_1_sums[7][68] [5:0] }), .sum({ \level_2_sums[7][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[141] [4:0] }), .sum({ \level_1_sums[7][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[143] [4:0] }), .sum({ \level_1_sums[7][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[7][71] [5:0] }),
     .b({ \level_1_sums[7][70] [5:0] }), .sum({ \level_2_sums[7][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[7][35] [6:0] }),
     .b({ \level_2_sums[7][34] [6:0] }), .sum({ \level_3_sums[7][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[7][17] [7:0] }),
     .b({ \level_3_sums[7][16] [7:0] }), .sum({ \level_4_sums[7][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[145] [4:0] }), .sum({ \level_1_sums[7][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[147] [4:0] }), .sum({ \level_1_sums[7][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[7][73] [5:0] }),
     .b({ \level_1_sums[7][72] [5:0] }), .sum({ \level_2_sums[7][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[149] [4:0] }), .sum({ \level_1_sums[7][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[151] [4:0] }), .sum({ \level_1_sums[7][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[7][75] [5:0] }),
     .b({ \level_1_sums[7][74] [5:0] }), .sum({ \level_2_sums[7][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[7][37] [6:0] }),
     .b({ \level_2_sums[7][36] [6:0] }), .sum({ \level_3_sums[7][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[153] [4:0] }), .sum({ \level_1_sums[7][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[155] [4:0] }), .sum({ \level_1_sums[7][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[7][77] [5:0] }),
     .b({ \level_1_sums[7][76] [5:0] }), .sum({ \level_2_sums[7][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[157] [4:0] }), .sum({ \level_1_sums[7][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[159] [4:0] }), .sum({ \level_1_sums[7][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[7][79] [5:0] }),
     .b({ \level_1_sums[7][78] [5:0] }), .sum({ \level_2_sums[7][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[7][39] [6:0] }),
     .b({ \level_2_sums[7][38] [6:0] }), .sum({ \level_3_sums[7][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[7][19] [7:0] }),
     .b({ \level_3_sums[7][18] [7:0] }), .sum({ \level_4_sums[7][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[7][9] [8:0] }),
     .b({ \level_4_sums[7][8] [8:0] }), .sum({ \level_5_sums[7][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[161] [4:0] }), .sum({ \level_1_sums[7][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[163] [4:0] }), .sum({ \level_1_sums[7][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[7][81] [5:0] }),
     .b({ \level_1_sums[7][80] [5:0] }), .sum({ \level_2_sums[7][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[165] [4:0] }), .sum({ \level_1_sums[7][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[167] [4:0] }), .sum({ \level_1_sums[7][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[7][83] [5:0] }),
     .b({ \level_1_sums[7][82] [5:0] }), .sum({ \level_2_sums[7][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[7][41] [6:0] }),
     .b({ \level_2_sums[7][40] [6:0] }), .sum({ \level_3_sums[7][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[169] [4:0] }), .sum({ \level_1_sums[7][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[171] [4:0] }), .sum({ \level_1_sums[7][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[7][85] [5:0] }),
     .b({ \level_1_sums[7][84] [5:0] }), .sum({ \level_2_sums[7][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[173] [4:0] }), .sum({ \level_1_sums[7][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[175] [4:0] }), .sum({ \level_1_sums[7][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[7][87] [5:0] }),
     .b({ \level_1_sums[7][86] [5:0] }), .sum({ \level_2_sums[7][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[7][43] [6:0] }),
     .b({ \level_2_sums[7][42] [6:0] }), .sum({ \level_3_sums[7][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[7][21] [7:0] }),
     .b({ \level_3_sums[7][20] [7:0] }), .sum({ \level_4_sums[7][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[177] [4:0] }), .sum({ \level_1_sums[7][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[179] [4:0] }), .sum({ \level_1_sums[7][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[7][89] [5:0] }),
     .b({ \level_1_sums[7][88] [5:0] }), .sum({ \level_2_sums[7][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[181] [4:0] }), .sum({ \level_1_sums[7][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[183] [4:0] }), .sum({ \level_1_sums[7][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[7][91] [5:0] }),
     .b({ \level_1_sums[7][90] [5:0] }), .sum({ \level_2_sums[7][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[7][45] [6:0] }),
     .b({ \level_2_sums[7][44] [6:0] }), .sum({ \level_3_sums[7][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[185] [4:0] }), .sum({ \level_1_sums[7][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[187] [4:0] }), .sum({ \level_1_sums[7][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[7][93] [5:0] }),
     .b({ \level_1_sums[7][92] [5:0] }), .sum({ \level_2_sums[7][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[189] [4:0] }), .sum({ \level_1_sums[7][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[191] [4:0] }), .sum({ \level_1_sums[7][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[7][95] [5:0] }),
     .b({ \level_1_sums[7][94] [5:0] }), .sum({ \level_2_sums[7][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[7][47] [6:0] }),
     .b({ \level_2_sums[7][46] [6:0] }), .sum({ \level_3_sums[7][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[7][23] [7:0] }),
     .b({ \level_3_sums[7][22] [7:0] }), .sum({ \level_4_sums[7][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[7][11] [8:0] }),
     .b({ \level_4_sums[7][10] [8:0] }), .sum({ \level_5_sums[7][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[7][5] [9:0] }),
     .b({ \level_5_sums[7][4] [9:0] }), .sum({ \level_6_sums[7][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[193] [4:0] }), .sum({ \level_1_sums[7][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[195] [4:0] }), .sum({ \level_1_sums[7][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[7][97] [5:0] }),
     .b({ \level_1_sums[7][96] [5:0] }), .sum({ \level_2_sums[7][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[197] [4:0] }), .sum({ \level_1_sums[7][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[199] [4:0] }), .sum({ \level_1_sums[7][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[7][99] [5:0] }),
     .b({ \level_1_sums[7][98] [5:0] }), .sum({ \level_2_sums[7][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[7][49] [6:0] }),
     .b({ \level_2_sums[7][48] [6:0] }), .sum({ \level_3_sums[7][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[201] [4:0] }), .sum({ \level_1_sums[7][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[203] [4:0] }), .sum({ \level_1_sums[7][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[7][101] [5:0] }),
     .b({ \level_1_sums[7][100] [5:0] }), .sum({ \level_2_sums[7][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[205] [4:0] }), .sum({ \level_1_sums[7][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[207] [4:0] }), .sum({ \level_1_sums[7][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[7][103] [5:0] }),
     .b({ \level_1_sums[7][102] [5:0] }), .sum({ \level_2_sums[7][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[7][51] [6:0] }),
     .b({ \level_2_sums[7][50] [6:0] }), .sum({ \level_3_sums[7][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[7][25] [7:0] }),
     .b({ \level_3_sums[7][24] [7:0] }), .sum({ \level_4_sums[7][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[209] [4:0] }), .sum({ \level_1_sums[7][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[211] [4:0] }), .sum({ \level_1_sums[7][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[7][105] [5:0] }),
     .b({ \level_1_sums[7][104] [5:0] }), .sum({ \level_2_sums[7][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[213] [4:0] }), .sum({ \level_1_sums[7][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[215] [4:0] }), .sum({ \level_1_sums[7][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[7][107] [5:0] }),
     .b({ \level_1_sums[7][106] [5:0] }), .sum({ \level_2_sums[7][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[7][53] [6:0] }),
     .b({ \level_2_sums[7][52] [6:0] }), .sum({ \level_3_sums[7][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[217] [4:0] }), .sum({ \level_1_sums[7][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[219] [4:0] }), .sum({ \level_1_sums[7][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[7][109] [5:0] }),
     .b({ \level_1_sums[7][108] [5:0] }), .sum({ \level_2_sums[7][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[221] [4:0] }), .sum({ \level_1_sums[7][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[223] [4:0] }), .sum({ \level_1_sums[7][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[7][111] [5:0] }),
     .b({ \level_1_sums[7][110] [5:0] }), .sum({ \level_2_sums[7][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[7][55] [6:0] }),
     .b({ \level_2_sums[7][54] [6:0] }), .sum({ \level_3_sums[7][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[7][27] [7:0] }),
     .b({ \level_3_sums[7][26] [7:0] }), .sum({ \level_4_sums[7][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[7][13] [8:0] }),
     .b({ \level_4_sums[7][12] [8:0] }), .sum({ \level_5_sums[7][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[225] [4:0] }), .sum({ \level_1_sums[7][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[227] [4:0] }), .sum({ \level_1_sums[7][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[7][113] [5:0] }),
     .b({ \level_1_sums[7][112] [5:0] }), .sum({ \level_2_sums[7][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[229] [4:0] }), .sum({ \level_1_sums[7][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[231] [4:0] }), .sum({ \level_1_sums[7][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[7][115] [5:0] }),
     .b({ \level_1_sums[7][114] [5:0] }), .sum({ \level_2_sums[7][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[7][57] [6:0] }),
     .b({ \level_2_sums[7][56] [6:0] }), .sum({ \level_3_sums[7][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[233] [4:0] }), .sum({ \level_1_sums[7][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[235] [4:0] }), .sum({ \level_1_sums[7][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[7][117] [5:0] }),
     .b({ \level_1_sums[7][116] [5:0] }), .sum({ \level_2_sums[7][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[237] [4:0] }), .sum({ \level_1_sums[7][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[239] [4:0] }), .sum({ \level_1_sums[7][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[7][119] [5:0] }),
     .b({ \level_1_sums[7][118] [5:0] }), .sum({ \level_2_sums[7][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[7][59] [6:0] }),
     .b({ \level_2_sums[7][58] [6:0] }), .sum({ \level_3_sums[7][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[7][29] [7:0] }),
     .b({ \level_3_sums[7][28] [7:0] }), .sum({ \level_4_sums[7][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[241] [4:0] }), .sum({ \level_1_sums[7][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[243] [4:0] }), .sum({ \level_1_sums[7][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[7][121] [5:0] }),
     .b({ \level_1_sums[7][120] [5:0] }), .sum({ \level_2_sums[7][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[245] [4:0] }), .sum({ \level_1_sums[7][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[247] [4:0] }), .sum({ \level_1_sums[7][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[7][123] [5:0] }),
     .b({ \level_1_sums[7][122] [5:0] }), .sum({ \level_2_sums[7][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[7][61] [6:0] }),
     .b({ \level_2_sums[7][60] [6:0] }), .sum({ \level_3_sums[7][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[249] [4:0] }), .sum({ \level_1_sums[7][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[251] [4:0] }), .sum({ \level_1_sums[7][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[7][125] [5:0] }),
     .b({ \level_1_sums[7][124] [5:0] }), .sum({ \level_2_sums[7][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[253] [4:0] }), .sum({ \level_1_sums[7][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[7].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[7].product_terms[255] [4:0] }), .sum({ \level_1_sums[7][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[7][127] [5:0] }),
     .b({ \level_1_sums[7][126] [5:0] }), .sum({ \level_2_sums[7][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[7][63] [6:0] }),
     .b({ \level_2_sums[7][62] [6:0] }), .sum({ \level_3_sums[7][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[7][31] [7:0] }),
     .b({ \level_3_sums[7][30] [7:0] }), .sum({ \level_4_sums[7][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[7][15] [8:0] }),
     .b({ \level_4_sums[7][14] [8:0] }), .sum({ \level_5_sums[7][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[7][7] [9:0] }),
     .b({ \level_5_sums[7][6] [9:0] }), .sum({ \level_6_sums[7][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[7][3] [9:0] }),
     .b({ \level_6_sums[7][2] [9:0] }), .sum({ \level_7_sums[7][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[7].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[7][0] [9:0] }),
     .b({ \level_7_sums[7][1] [9:0] }), .sum({ \level_8_sums[7] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[8].relu_inst (.in_data({ \final_sums[8] [9:0] }), .out_data({ \out_sig[8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[1] [4:0] }), .sum({ \level_1_sums[8][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[3] [4:0] }), .sum({ \level_1_sums[8][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[8][1] [5:0] }),
     .b({ \level_1_sums[8][0] [5:0] }), .sum({ \level_2_sums[8][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[5] [4:0] }), .sum({ \level_1_sums[8][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[7] [4:0] }), .sum({ \level_1_sums[8][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[8][3] [5:0] }),
     .b({ \level_1_sums[8][2] [5:0] }), .sum({ \level_2_sums[8][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[8][1] [6:0] }),
     .b({ \level_2_sums[8][0] [6:0] }), .sum({ \level_3_sums[8][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[9] [4:0] }), .sum({ \level_1_sums[8][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[11] [4:0] }), .sum({ \level_1_sums[8][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[8][5] [5:0] }),
     .b({ \level_1_sums[8][4] [5:0] }), .sum({ \level_2_sums[8][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[13] [4:0] }), .sum({ \level_1_sums[8][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[15] [4:0] }), .sum({ \level_1_sums[8][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[8][7] [5:0] }),
     .b({ \level_1_sums[8][6] [5:0] }), .sum({ \level_2_sums[8][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[8][3] [6:0] }),
     .b({ \level_2_sums[8][2] [6:0] }), .sum({ \level_3_sums[8][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[8][1] [7:0] }),
     .b({ \level_3_sums[8][0] [7:0] }), .sum({ \level_4_sums[8][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[17] [4:0] }), .sum({ \level_1_sums[8][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[19] [4:0] }), .sum({ \level_1_sums[8][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[8][9] [5:0] }),
     .b({ \level_1_sums[8][8] [5:0] }), .sum({ \level_2_sums[8][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[21] [4:0] }), .sum({ \level_1_sums[8][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[23] [4:0] }), .sum({ \level_1_sums[8][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[8][11] [5:0] }),
     .b({ \level_1_sums[8][10] [5:0] }), .sum({ \level_2_sums[8][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[8][5] [6:0] }),
     .b({ \level_2_sums[8][4] [6:0] }), .sum({ \level_3_sums[8][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[25] [4:0] }), .sum({ \level_1_sums[8][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[27] [4:0] }), .sum({ \level_1_sums[8][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[8][13] [5:0] }),
     .b({ \level_1_sums[8][12] [5:0] }), .sum({ \level_2_sums[8][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[29] [4:0] }), .sum({ \level_1_sums[8][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[31] [4:0] }), .sum({ \level_1_sums[8][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[8][15] [5:0] }),
     .b({ \level_1_sums[8][14] [5:0] }), .sum({ \level_2_sums[8][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[8][7] [6:0] }),
     .b({ \level_2_sums[8][6] [6:0] }), .sum({ \level_3_sums[8][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[8][3] [7:0] }),
     .b({ \level_3_sums[8][2] [7:0] }), .sum({ \level_4_sums[8][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[8][1] [8:0] }),
     .b({ \level_4_sums[8][0] [8:0] }), .sum({ \level_5_sums[8][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[33] [4:0] }), .sum({ \level_1_sums[8][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[35] [4:0] }), .sum({ \level_1_sums[8][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[8][17] [5:0] }),
     .b({ \level_1_sums[8][16] [5:0] }), .sum({ \level_2_sums[8][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[37] [4:0] }), .sum({ \level_1_sums[8][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[39] [4:0] }), .sum({ \level_1_sums[8][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[8][19] [5:0] }),
     .b({ \level_1_sums[8][18] [5:0] }), .sum({ \level_2_sums[8][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[8][9] [6:0] }),
     .b({ \level_2_sums[8][8] [6:0] }), .sum({ \level_3_sums[8][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[41] [4:0] }), .sum({ \level_1_sums[8][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[43] [4:0] }), .sum({ \level_1_sums[8][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[8][21] [5:0] }),
     .b({ \level_1_sums[8][20] [5:0] }), .sum({ \level_2_sums[8][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[45] [4:0] }), .sum({ \level_1_sums[8][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[47] [4:0] }), .sum({ \level_1_sums[8][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[8][23] [5:0] }),
     .b({ \level_1_sums[8][22] [5:0] }), .sum({ \level_2_sums[8][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[8][11] [6:0] }),
     .b({ \level_2_sums[8][10] [6:0] }), .sum({ \level_3_sums[8][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[8][5] [7:0] }),
     .b({ \level_3_sums[8][4] [7:0] }), .sum({ \level_4_sums[8][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[49] [4:0] }), .sum({ \level_1_sums[8][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[51] [4:0] }), .sum({ \level_1_sums[8][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[8][25] [5:0] }),
     .b({ \level_1_sums[8][24] [5:0] }), .sum({ \level_2_sums[8][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[53] [4:0] }), .sum({ \level_1_sums[8][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[55] [4:0] }), .sum({ \level_1_sums[8][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[8][27] [5:0] }),
     .b({ \level_1_sums[8][26] [5:0] }), .sum({ \level_2_sums[8][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[8][13] [6:0] }),
     .b({ \level_2_sums[8][12] [6:0] }), .sum({ \level_3_sums[8][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[57] [4:0] }), .sum({ \level_1_sums[8][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[59] [4:0] }), .sum({ \level_1_sums[8][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[8][29] [5:0] }),
     .b({ \level_1_sums[8][28] [5:0] }), .sum({ \level_2_sums[8][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[61] [4:0] }), .sum({ \level_1_sums[8][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[63] [4:0] }), .sum({ \level_1_sums[8][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[8][31] [5:0] }),
     .b({ \level_1_sums[8][30] [5:0] }), .sum({ \level_2_sums[8][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[8][15] [6:0] }),
     .b({ \level_2_sums[8][14] [6:0] }), .sum({ \level_3_sums[8][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[8][7] [7:0] }),
     .b({ \level_3_sums[8][6] [7:0] }), .sum({ \level_4_sums[8][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[8][3] [8:0] }),
     .b({ \level_4_sums[8][2] [8:0] }), .sum({ \level_5_sums[8][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[8][1] [9:0] }),
     .b({ \level_5_sums[8][0] [9:0] }), .sum({ \level_6_sums[8][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[65] [4:0] }), .sum({ \level_1_sums[8][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[67] [4:0] }), .sum({ \level_1_sums[8][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[8][33] [5:0] }),
     .b({ \level_1_sums[8][32] [5:0] }), .sum({ \level_2_sums[8][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[69] [4:0] }), .sum({ \level_1_sums[8][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[71] [4:0] }), .sum({ \level_1_sums[8][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[8][35] [5:0] }),
     .b({ \level_1_sums[8][34] [5:0] }), .sum({ \level_2_sums[8][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[8][17] [6:0] }),
     .b({ \level_2_sums[8][16] [6:0] }), .sum({ \level_3_sums[8][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[73] [4:0] }), .sum({ \level_1_sums[8][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[75] [4:0] }), .sum({ \level_1_sums[8][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[8][37] [5:0] }),
     .b({ \level_1_sums[8][36] [5:0] }), .sum({ \level_2_sums[8][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[77] [4:0] }), .sum({ \level_1_sums[8][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[79] [4:0] }), .sum({ \level_1_sums[8][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[8][39] [5:0] }),
     .b({ \level_1_sums[8][38] [5:0] }), .sum({ \level_2_sums[8][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[8][19] [6:0] }),
     .b({ \level_2_sums[8][18] [6:0] }), .sum({ \level_3_sums[8][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[8][9] [7:0] }),
     .b({ \level_3_sums[8][8] [7:0] }), .sum({ \level_4_sums[8][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[81] [4:0] }), .sum({ \level_1_sums[8][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[83] [4:0] }), .sum({ \level_1_sums[8][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[8][41] [5:0] }),
     .b({ \level_1_sums[8][40] [5:0] }), .sum({ \level_2_sums[8][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[85] [4:0] }), .sum({ \level_1_sums[8][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[87] [4:0] }), .sum({ \level_1_sums[8][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[8][43] [5:0] }),
     .b({ \level_1_sums[8][42] [5:0] }), .sum({ \level_2_sums[8][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[8][21] [6:0] }),
     .b({ \level_2_sums[8][20] [6:0] }), .sum({ \level_3_sums[8][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[89] [4:0] }), .sum({ \level_1_sums[8][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[91] [4:0] }), .sum({ \level_1_sums[8][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[8][45] [5:0] }),
     .b({ \level_1_sums[8][44] [5:0] }), .sum({ \level_2_sums[8][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[93] [4:0] }), .sum({ \level_1_sums[8][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[95] [4:0] }), .sum({ \level_1_sums[8][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[8][47] [5:0] }),
     .b({ \level_1_sums[8][46] [5:0] }), .sum({ \level_2_sums[8][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[8][23] [6:0] }),
     .b({ \level_2_sums[8][22] [6:0] }), .sum({ \level_3_sums[8][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[8][11] [7:0] }),
     .b({ \level_3_sums[8][10] [7:0] }), .sum({ \level_4_sums[8][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[8][5] [8:0] }),
     .b({ \level_4_sums[8][4] [8:0] }), .sum({ \level_5_sums[8][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[97] [4:0] }), .sum({ \level_1_sums[8][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[99] [4:0] }), .sum({ \level_1_sums[8][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[8][49] [5:0] }),
     .b({ \level_1_sums[8][48] [5:0] }), .sum({ \level_2_sums[8][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[101] [4:0] }), .sum({ \level_1_sums[8][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[103] [4:0] }), .sum({ \level_1_sums[8][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[8][51] [5:0] }),
     .b({ \level_1_sums[8][50] [5:0] }), .sum({ \level_2_sums[8][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[8][25] [6:0] }),
     .b({ \level_2_sums[8][24] [6:0] }), .sum({ \level_3_sums[8][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[105] [4:0] }), .sum({ \level_1_sums[8][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[107] [4:0] }), .sum({ \level_1_sums[8][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[8][53] [5:0] }),
     .b({ \level_1_sums[8][52] [5:0] }), .sum({ \level_2_sums[8][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[109] [4:0] }), .sum({ \level_1_sums[8][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[111] [4:0] }), .sum({ \level_1_sums[8][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[8][55] [5:0] }),
     .b({ \level_1_sums[8][54] [5:0] }), .sum({ \level_2_sums[8][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[8][27] [6:0] }),
     .b({ \level_2_sums[8][26] [6:0] }), .sum({ \level_3_sums[8][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[8][13] [7:0] }),
     .b({ \level_3_sums[8][12] [7:0] }), .sum({ \level_4_sums[8][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[113] [4:0] }), .sum({ \level_1_sums[8][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[115] [4:0] }), .sum({ \level_1_sums[8][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[8][57] [5:0] }),
     .b({ \level_1_sums[8][56] [5:0] }), .sum({ \level_2_sums[8][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[117] [4:0] }), .sum({ \level_1_sums[8][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[119] [4:0] }), .sum({ \level_1_sums[8][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[8][59] [5:0] }),
     .b({ \level_1_sums[8][58] [5:0] }), .sum({ \level_2_sums[8][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[8][29] [6:0] }),
     .b({ \level_2_sums[8][28] [6:0] }), .sum({ \level_3_sums[8][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[121] [4:0] }), .sum({ \level_1_sums[8][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[123] [4:0] }), .sum({ \level_1_sums[8][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[8][61] [5:0] }),
     .b({ \level_1_sums[8][60] [5:0] }), .sum({ \level_2_sums[8][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[125] [4:0] }), .sum({ \level_1_sums[8][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[127] [4:0] }), .sum({ \level_1_sums[8][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[8][63] [5:0] }),
     .b({ \level_1_sums[8][62] [5:0] }), .sum({ \level_2_sums[8][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[8][31] [6:0] }),
     .b({ \level_2_sums[8][30] [6:0] }), .sum({ \level_3_sums[8][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[8][15] [7:0] }),
     .b({ \level_3_sums[8][14] [7:0] }), .sum({ \level_4_sums[8][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[8][7] [8:0] }),
     .b({ \level_4_sums[8][6] [8:0] }), .sum({ \level_5_sums[8][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[8][3] [9:0] }),
     .b({ \level_5_sums[8][2] [9:0] }), .sum({ \level_6_sums[8][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[8][1] [9:0] }),
     .b({ \level_6_sums[8][0] [9:0] }), .sum({ \level_7_sums[8][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[129] [4:0] }), .sum({ \level_1_sums[8][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[131] [4:0] }), .sum({ \level_1_sums[8][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[8][65] [5:0] }),
     .b({ \level_1_sums[8][64] [5:0] }), .sum({ \level_2_sums[8][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[133] [4:0] }), .sum({ \level_1_sums[8][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[135] [4:0] }), .sum({ \level_1_sums[8][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[8][67] [5:0] }),
     .b({ \level_1_sums[8][66] [5:0] }), .sum({ \level_2_sums[8][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[8][33] [6:0] }),
     .b({ \level_2_sums[8][32] [6:0] }), .sum({ \level_3_sums[8][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[137] [4:0] }), .sum({ \level_1_sums[8][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[139] [4:0] }), .sum({ \level_1_sums[8][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[8][69] [5:0] }),
     .b({ \level_1_sums[8][68] [5:0] }), .sum({ \level_2_sums[8][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[141] [4:0] }), .sum({ \level_1_sums[8][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[143] [4:0] }), .sum({ \level_1_sums[8][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[8][71] [5:0] }),
     .b({ \level_1_sums[8][70] [5:0] }), .sum({ \level_2_sums[8][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[8][35] [6:0] }),
     .b({ \level_2_sums[8][34] [6:0] }), .sum({ \level_3_sums[8][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[8][17] [7:0] }),
     .b({ \level_3_sums[8][16] [7:0] }), .sum({ \level_4_sums[8][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[145] [4:0] }), .sum({ \level_1_sums[8][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[147] [4:0] }), .sum({ \level_1_sums[8][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[8][73] [5:0] }),
     .b({ \level_1_sums[8][72] [5:0] }), .sum({ \level_2_sums[8][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[149] [4:0] }), .sum({ \level_1_sums[8][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[151] [4:0] }), .sum({ \level_1_sums[8][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[8][75] [5:0] }),
     .b({ \level_1_sums[8][74] [5:0] }), .sum({ \level_2_sums[8][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[8][37] [6:0] }),
     .b({ \level_2_sums[8][36] [6:0] }), .sum({ \level_3_sums[8][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[153] [4:0] }), .sum({ \level_1_sums[8][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[155] [4:0] }), .sum({ \level_1_sums[8][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[8][77] [5:0] }),
     .b({ \level_1_sums[8][76] [5:0] }), .sum({ \level_2_sums[8][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[157] [4:0] }), .sum({ \level_1_sums[8][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[159] [4:0] }), .sum({ \level_1_sums[8][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[8][79] [5:0] }),
     .b({ \level_1_sums[8][78] [5:0] }), .sum({ \level_2_sums[8][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[8][39] [6:0] }),
     .b({ \level_2_sums[8][38] [6:0] }), .sum({ \level_3_sums[8][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[8][19] [7:0] }),
     .b({ \level_3_sums[8][18] [7:0] }), .sum({ \level_4_sums[8][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[8][9] [8:0] }),
     .b({ \level_4_sums[8][8] [8:0] }), .sum({ \level_5_sums[8][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[161] [4:0] }), .sum({ \level_1_sums[8][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[163] [4:0] }), .sum({ \level_1_sums[8][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[8][81] [5:0] }),
     .b({ \level_1_sums[8][80] [5:0] }), .sum({ \level_2_sums[8][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[165] [4:0] }), .sum({ \level_1_sums[8][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[167] [4:0] }), .sum({ \level_1_sums[8][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[8][83] [5:0] }),
     .b({ \level_1_sums[8][82] [5:0] }), .sum({ \level_2_sums[8][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[8][41] [6:0] }),
     .b({ \level_2_sums[8][40] [6:0] }), .sum({ \level_3_sums[8][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[169] [4:0] }), .sum({ \level_1_sums[8][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[171] [4:0] }), .sum({ \level_1_sums[8][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[8][85] [5:0] }),
     .b({ \level_1_sums[8][84] [5:0] }), .sum({ \level_2_sums[8][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[173] [4:0] }), .sum({ \level_1_sums[8][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[175] [4:0] }), .sum({ \level_1_sums[8][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[8][87] [5:0] }),
     .b({ \level_1_sums[8][86] [5:0] }), .sum({ \level_2_sums[8][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[8][43] [6:0] }),
     .b({ \level_2_sums[8][42] [6:0] }), .sum({ \level_3_sums[8][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[8][21] [7:0] }),
     .b({ \level_3_sums[8][20] [7:0] }), .sum({ \level_4_sums[8][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[177] [4:0] }), .sum({ \level_1_sums[8][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[179] [4:0] }), .sum({ \level_1_sums[8][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[8][89] [5:0] }),
     .b({ \level_1_sums[8][88] [5:0] }), .sum({ \level_2_sums[8][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[181] [4:0] }), .sum({ \level_1_sums[8][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[183] [4:0] }), .sum({ \level_1_sums[8][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[8][91] [5:0] }),
     .b({ \level_1_sums[8][90] [5:0] }), .sum({ \level_2_sums[8][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[8][45] [6:0] }),
     .b({ \level_2_sums[8][44] [6:0] }), .sum({ \level_3_sums[8][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[185] [4:0] }), .sum({ \level_1_sums[8][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[187] [4:0] }), .sum({ \level_1_sums[8][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[8][93] [5:0] }),
     .b({ \level_1_sums[8][92] [5:0] }), .sum({ \level_2_sums[8][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[189] [4:0] }), .sum({ \level_1_sums[8][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[191] [4:0] }), .sum({ \level_1_sums[8][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[8][95] [5:0] }),
     .b({ \level_1_sums[8][94] [5:0] }), .sum({ \level_2_sums[8][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[8][47] [6:0] }),
     .b({ \level_2_sums[8][46] [6:0] }), .sum({ \level_3_sums[8][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[8][23] [7:0] }),
     .b({ \level_3_sums[8][22] [7:0] }), .sum({ \level_4_sums[8][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[8][11] [8:0] }),
     .b({ \level_4_sums[8][10] [8:0] }), .sum({ \level_5_sums[8][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[8][5] [9:0] }),
     .b({ \level_5_sums[8][4] [9:0] }), .sum({ \level_6_sums[8][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[193] [4:0] }), .sum({ \level_1_sums[8][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[195] [4:0] }), .sum({ \level_1_sums[8][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[8][97] [5:0] }),
     .b({ \level_1_sums[8][96] [5:0] }), .sum({ \level_2_sums[8][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[197] [4:0] }), .sum({ \level_1_sums[8][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[199] [4:0] }), .sum({ \level_1_sums[8][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[8][99] [5:0] }),
     .b({ \level_1_sums[8][98] [5:0] }), .sum({ \level_2_sums[8][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[8][49] [6:0] }),
     .b({ \level_2_sums[8][48] [6:0] }), .sum({ \level_3_sums[8][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[201] [4:0] }), .sum({ \level_1_sums[8][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[203] [4:0] }), .sum({ \level_1_sums[8][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[8][101] [5:0] }),
     .b({ \level_1_sums[8][100] [5:0] }), .sum({ \level_2_sums[8][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[205] [4:0] }), .sum({ \level_1_sums[8][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[207] [4:0] }), .sum({ \level_1_sums[8][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[8][103] [5:0] }),
     .b({ \level_1_sums[8][102] [5:0] }), .sum({ \level_2_sums[8][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[8][51] [6:0] }),
     .b({ \level_2_sums[8][50] [6:0] }), .sum({ \level_3_sums[8][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[8][25] [7:0] }),
     .b({ \level_3_sums[8][24] [7:0] }), .sum({ \level_4_sums[8][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[209] [4:0] }), .sum({ \level_1_sums[8][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[211] [4:0] }), .sum({ \level_1_sums[8][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[8][105] [5:0] }),
     .b({ \level_1_sums[8][104] [5:0] }), .sum({ \level_2_sums[8][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[213] [4:0] }), .sum({ \level_1_sums[8][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[215] [4:0] }), .sum({ \level_1_sums[8][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[8][107] [5:0] }),
     .b({ \level_1_sums[8][106] [5:0] }), .sum({ \level_2_sums[8][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[8][53] [6:0] }),
     .b({ \level_2_sums[8][52] [6:0] }), .sum({ \level_3_sums[8][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[217] [4:0] }), .sum({ \level_1_sums[8][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[219] [4:0] }), .sum({ \level_1_sums[8][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[8][109] [5:0] }),
     .b({ \level_1_sums[8][108] [5:0] }), .sum({ \level_2_sums[8][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[221] [4:0] }), .sum({ \level_1_sums[8][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[223] [4:0] }), .sum({ \level_1_sums[8][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[8][111] [5:0] }),
     .b({ \level_1_sums[8][110] [5:0] }), .sum({ \level_2_sums[8][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[8][55] [6:0] }),
     .b({ \level_2_sums[8][54] [6:0] }), .sum({ \level_3_sums[8][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[8][27] [7:0] }),
     .b({ \level_3_sums[8][26] [7:0] }), .sum({ \level_4_sums[8][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[8][13] [8:0] }),
     .b({ \level_4_sums[8][12] [8:0] }), .sum({ \level_5_sums[8][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[225] [4:0] }), .sum({ \level_1_sums[8][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[227] [4:0] }), .sum({ \level_1_sums[8][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[8][113] [5:0] }),
     .b({ \level_1_sums[8][112] [5:0] }), .sum({ \level_2_sums[8][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[229] [4:0] }), .sum({ \level_1_sums[8][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[231] [4:0] }), .sum({ \level_1_sums[8][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[8][115] [5:0] }),
     .b({ \level_1_sums[8][114] [5:0] }), .sum({ \level_2_sums[8][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[8][57] [6:0] }),
     .b({ \level_2_sums[8][56] [6:0] }), .sum({ \level_3_sums[8][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[233] [4:0] }), .sum({ \level_1_sums[8][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[235] [4:0] }), .sum({ \level_1_sums[8][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[8][117] [5:0] }),
     .b({ \level_1_sums[8][116] [5:0] }), .sum({ \level_2_sums[8][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[237] [4:0] }), .sum({ \level_1_sums[8][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[239] [4:0] }), .sum({ \level_1_sums[8][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[8][119] [5:0] }),
     .b({ \level_1_sums[8][118] [5:0] }), .sum({ \level_2_sums[8][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[8][59] [6:0] }),
     .b({ \level_2_sums[8][58] [6:0] }), .sum({ \level_3_sums[8][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[8][29] [7:0] }),
     .b({ \level_3_sums[8][28] [7:0] }), .sum({ \level_4_sums[8][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[241] [4:0] }), .sum({ \level_1_sums[8][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[243] [4:0] }), .sum({ \level_1_sums[8][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[8][121] [5:0] }),
     .b({ \level_1_sums[8][120] [5:0] }), .sum({ \level_2_sums[8][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[245] [4:0] }), .sum({ \level_1_sums[8][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[247] [4:0] }), .sum({ \level_1_sums[8][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[8][123] [5:0] }),
     .b({ \level_1_sums[8][122] [5:0] }), .sum({ \level_2_sums[8][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[8][61] [6:0] }),
     .b({ \level_2_sums[8][60] [6:0] }), .sum({ \level_3_sums[8][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[249] [4:0] }), .sum({ \level_1_sums[8][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[251] [4:0] }), .sum({ \level_1_sums[8][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[8][125] [5:0] }),
     .b({ \level_1_sums[8][124] [5:0] }), .sum({ \level_2_sums[8][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[253] [4:0] }), .sum({ \level_1_sums[8][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[8].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[8].product_terms[255] [4:0] }), .sum({ \level_1_sums[8][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[8][127] [5:0] }),
     .b({ \level_1_sums[8][126] [5:0] }), .sum({ \level_2_sums[8][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[8][63] [6:0] }),
     .b({ \level_2_sums[8][62] [6:0] }), .sum({ \level_3_sums[8][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[8][31] [7:0] }),
     .b({ \level_3_sums[8][30] [7:0] }), .sum({ \level_4_sums[8][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[8][15] [8:0] }),
     .b({ \level_4_sums[8][14] [8:0] }), .sum({ \level_5_sums[8][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[8][7] [9:0] }),
     .b({ \level_5_sums[8][6] [9:0] }), .sum({ \level_6_sums[8][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[8][3] [9:0] }),
     .b({ \level_6_sums[8][2] [9:0] }), .sum({ \level_7_sums[8][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[8].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[8][0] [9:0] }),
     .b({ \level_7_sums[8][1] [9:0] }), .sum({ \level_8_sums[8] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[9].relu_inst (.in_data({ \final_sums[9] [9:0] }), .out_data({ \out_sig[9] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[1] [4:0] }), .sum({ \level_1_sums[9][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[3] [4:0] }), .sum({ \level_1_sums[9][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[9][1] [5:0] }),
     .b({ \level_1_sums[9][0] [5:0] }), .sum({ \level_2_sums[9][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[5] [4:0] }), .sum({ \level_1_sums[9][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[7] [4:0] }), .sum({ \level_1_sums[9][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[9][3] [5:0] }),
     .b({ \level_1_sums[9][2] [5:0] }), .sum({ \level_2_sums[9][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[9][1] [6:0] }),
     .b({ \level_2_sums[9][0] [6:0] }), .sum({ \level_3_sums[9][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[9] [4:0] }), .sum({ \level_1_sums[9][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[11] [4:0] }), .sum({ \level_1_sums[9][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[9][5] [5:0] }),
     .b({ \level_1_sums[9][4] [5:0] }), .sum({ \level_2_sums[9][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[13] [4:0] }), .sum({ \level_1_sums[9][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[15] [4:0] }), .sum({ \level_1_sums[9][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[9][7] [5:0] }),
     .b({ \level_1_sums[9][6] [5:0] }), .sum({ \level_2_sums[9][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[9][3] [6:0] }),
     .b({ \level_2_sums[9][2] [6:0] }), .sum({ \level_3_sums[9][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[9][1] [7:0] }),
     .b({ \level_3_sums[9][0] [7:0] }), .sum({ \level_4_sums[9][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[17] [4:0] }), .sum({ \level_1_sums[9][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[19] [4:0] }), .sum({ \level_1_sums[9][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[9][9] [5:0] }),
     .b({ \level_1_sums[9][8] [5:0] }), .sum({ \level_2_sums[9][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[21] [4:0] }), .sum({ \level_1_sums[9][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[23] [4:0] }), .sum({ \level_1_sums[9][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[9][11] [5:0] }),
     .b({ \level_1_sums[9][10] [5:0] }), .sum({ \level_2_sums[9][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[9][5] [6:0] }),
     .b({ \level_2_sums[9][4] [6:0] }), .sum({ \level_3_sums[9][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[25] [4:0] }), .sum({ \level_1_sums[9][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[27] [4:0] }), .sum({ \level_1_sums[9][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[9][13] [5:0] }),
     .b({ \level_1_sums[9][12] [5:0] }), .sum({ \level_2_sums[9][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[29] [4:0] }), .sum({ \level_1_sums[9][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[31] [4:0] }), .sum({ \level_1_sums[9][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[9][15] [5:0] }),
     .b({ \level_1_sums[9][14] [5:0] }), .sum({ \level_2_sums[9][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[9][7] [6:0] }),
     .b({ \level_2_sums[9][6] [6:0] }), .sum({ \level_3_sums[9][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[9][3] [7:0] }),
     .b({ \level_3_sums[9][2] [7:0] }), .sum({ \level_4_sums[9][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[9][1] [8:0] }),
     .b({ \level_4_sums[9][0] [8:0] }), .sum({ \level_5_sums[9][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[33] [4:0] }), .sum({ \level_1_sums[9][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[35] [4:0] }), .sum({ \level_1_sums[9][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[9][17] [5:0] }),
     .b({ \level_1_sums[9][16] [5:0] }), .sum({ \level_2_sums[9][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[37] [4:0] }), .sum({ \level_1_sums[9][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[39] [4:0] }), .sum({ \level_1_sums[9][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[9][19] [5:0] }),
     .b({ \level_1_sums[9][18] [5:0] }), .sum({ \level_2_sums[9][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[9][9] [6:0] }),
     .b({ \level_2_sums[9][8] [6:0] }), .sum({ \level_3_sums[9][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[41] [4:0] }), .sum({ \level_1_sums[9][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[43] [4:0] }), .sum({ \level_1_sums[9][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[9][21] [5:0] }),
     .b({ \level_1_sums[9][20] [5:0] }), .sum({ \level_2_sums[9][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[45] [4:0] }), .sum({ \level_1_sums[9][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[47] [4:0] }), .sum({ \level_1_sums[9][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[9][23] [5:0] }),
     .b({ \level_1_sums[9][22] [5:0] }), .sum({ \level_2_sums[9][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[9][11] [6:0] }),
     .b({ \level_2_sums[9][10] [6:0] }), .sum({ \level_3_sums[9][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[9][5] [7:0] }),
     .b({ \level_3_sums[9][4] [7:0] }), .sum({ \level_4_sums[9][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[49] [4:0] }), .sum({ \level_1_sums[9][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[51] [4:0] }), .sum({ \level_1_sums[9][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[9][25] [5:0] }),
     .b({ \level_1_sums[9][24] [5:0] }), .sum({ \level_2_sums[9][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[53] [4:0] }), .sum({ \level_1_sums[9][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[55] [4:0] }), .sum({ \level_1_sums[9][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[9][27] [5:0] }),
     .b({ \level_1_sums[9][26] [5:0] }), .sum({ \level_2_sums[9][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[9][13] [6:0] }),
     .b({ \level_2_sums[9][12] [6:0] }), .sum({ \level_3_sums[9][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[57] [4:0] }), .sum({ \level_1_sums[9][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[59] [4:0] }), .sum({ \level_1_sums[9][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[9][29] [5:0] }),
     .b({ \level_1_sums[9][28] [5:0] }), .sum({ \level_2_sums[9][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[61] [4:0] }), .sum({ \level_1_sums[9][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[63] [4:0] }), .sum({ \level_1_sums[9][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[9][31] [5:0] }),
     .b({ \level_1_sums[9][30] [5:0] }), .sum({ \level_2_sums[9][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[9][15] [6:0] }),
     .b({ \level_2_sums[9][14] [6:0] }), .sum({ \level_3_sums[9][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[9][7] [7:0] }),
     .b({ \level_3_sums[9][6] [7:0] }), .sum({ \level_4_sums[9][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[9][3] [8:0] }),
     .b({ \level_4_sums[9][2] [8:0] }), .sum({ \level_5_sums[9][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[9][1] [9:0] }),
     .b({ \level_5_sums[9][0] [9:0] }), .sum({ \level_6_sums[9][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[65] [4:0] }), .sum({ \level_1_sums[9][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[67] [4:0] }), .sum({ \level_1_sums[9][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[9][33] [5:0] }),
     .b({ \level_1_sums[9][32] [5:0] }), .sum({ \level_2_sums[9][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[69] [4:0] }), .sum({ \level_1_sums[9][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[71] [4:0] }), .sum({ \level_1_sums[9][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[9][35] [5:0] }),
     .b({ \level_1_sums[9][34] [5:0] }), .sum({ \level_2_sums[9][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[9][17] [6:0] }),
     .b({ \level_2_sums[9][16] [6:0] }), .sum({ \level_3_sums[9][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[73] [4:0] }), .sum({ \level_1_sums[9][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[75] [4:0] }), .sum({ \level_1_sums[9][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[9][37] [5:0] }),
     .b({ \level_1_sums[9][36] [5:0] }), .sum({ \level_2_sums[9][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[77] [4:0] }), .sum({ \level_1_sums[9][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[79] [4:0] }), .sum({ \level_1_sums[9][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[9][39] [5:0] }),
     .b({ \level_1_sums[9][38] [5:0] }), .sum({ \level_2_sums[9][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[9][19] [6:0] }),
     .b({ \level_2_sums[9][18] [6:0] }), .sum({ \level_3_sums[9][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[9][9] [7:0] }),
     .b({ \level_3_sums[9][8] [7:0] }), .sum({ \level_4_sums[9][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[81] [4:0] }), .sum({ \level_1_sums[9][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[83] [4:0] }), .sum({ \level_1_sums[9][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[9][41] [5:0] }),
     .b({ \level_1_sums[9][40] [5:0] }), .sum({ \level_2_sums[9][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[85] [4:0] }), .sum({ \level_1_sums[9][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[87] [4:0] }), .sum({ \level_1_sums[9][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[9][43] [5:0] }),
     .b({ \level_1_sums[9][42] [5:0] }), .sum({ \level_2_sums[9][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[9][21] [6:0] }),
     .b({ \level_2_sums[9][20] [6:0] }), .sum({ \level_3_sums[9][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[89] [4:0] }), .sum({ \level_1_sums[9][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[91] [4:0] }), .sum({ \level_1_sums[9][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[9][45] [5:0] }),
     .b({ \level_1_sums[9][44] [5:0] }), .sum({ \level_2_sums[9][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[93] [4:0] }), .sum({ \level_1_sums[9][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[95] [4:0] }), .sum({ \level_1_sums[9][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[9][47] [5:0] }),
     .b({ \level_1_sums[9][46] [5:0] }), .sum({ \level_2_sums[9][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[9][23] [6:0] }),
     .b({ \level_2_sums[9][22] [6:0] }), .sum({ \level_3_sums[9][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[9][11] [7:0] }),
     .b({ \level_3_sums[9][10] [7:0] }), .sum({ \level_4_sums[9][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[9][5] [8:0] }),
     .b({ \level_4_sums[9][4] [8:0] }), .sum({ \level_5_sums[9][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[97] [4:0] }), .sum({ \level_1_sums[9][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[99] [4:0] }), .sum({ \level_1_sums[9][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[9][49] [5:0] }),
     .b({ \level_1_sums[9][48] [5:0] }), .sum({ \level_2_sums[9][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[101] [4:0] }), .sum({ \level_1_sums[9][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[103] [4:0] }), .sum({ \level_1_sums[9][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[9][51] [5:0] }),
     .b({ \level_1_sums[9][50] [5:0] }), .sum({ \level_2_sums[9][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[103].adder_octets.adder_inst (.a({ \level_2_sums[9][25] [6:0] }),
     .b({ \level_2_sums[9][24] [6:0] }), .sum({ \level_3_sums[9][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[105] [4:0] }), .sum({ \level_1_sums[9][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[107] [4:0] }), .sum({ \level_1_sums[9][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[9][53] [5:0] }),
     .b({ \level_1_sums[9][52] [5:0] }), .sum({ \level_2_sums[9][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[109] [4:0] }), .sum({ \level_1_sums[9][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[111] [4:0] }), .sum({ \level_1_sums[9][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[9][55] [5:0] }),
     .b({ \level_1_sums[9][54] [5:0] }), .sum({ \level_2_sums[9][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[111].adder_octets.adder_inst (.a({ \level_2_sums[9][27] [6:0] }),
     .b({ \level_2_sums[9][26] [6:0] }), .sum({ \level_3_sums[9][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[9][13] [7:0] }),
     .b({ \level_3_sums[9][12] [7:0] }), .sum({ \level_4_sums[9][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[113] [4:0] }), .sum({ \level_1_sums[9][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[115] [4:0] }), .sum({ \level_1_sums[9][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[9][57] [5:0] }),
     .b({ \level_1_sums[9][56] [5:0] }), .sum({ \level_2_sums[9][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[117] [4:0] }), .sum({ \level_1_sums[9][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[119] [4:0] }), .sum({ \level_1_sums[9][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[9][59] [5:0] }),
     .b({ \level_1_sums[9][58] [5:0] }), .sum({ \level_2_sums[9][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[119].adder_octets.adder_inst (.a({ \level_2_sums[9][29] [6:0] }),
     .b({ \level_2_sums[9][28] [6:0] }), .sum({ \level_3_sums[9][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[121] [4:0] }), .sum({ \level_1_sums[9][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[123] [4:0] }), .sum({ \level_1_sums[9][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[9][61] [5:0] }),
     .b({ \level_1_sums[9][60] [5:0] }), .sum({ \level_2_sums[9][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[125] [4:0] }), .sum({ \level_1_sums[9][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[127] [4:0] }), .sum({ \level_1_sums[9][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[9][63] [5:0] }),
     .b({ \level_1_sums[9][62] [5:0] }), .sum({ \level_2_sums[9][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_octets.adder_inst (.a({ \level_2_sums[9][31] [6:0] }),
     .b({ \level_2_sums[9][30] [6:0] }), .sum({ \level_3_sums[9][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[9][15] [7:0] }),
     .b({ \level_3_sums[9][14] [7:0] }), .sum({ \level_4_sums[9][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[9][7] [8:0] }),
     .b({ \level_4_sums[9][6] [8:0] }), .sum({ \level_5_sums[9][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[9][3] [9:0] }),
     .b({ \level_5_sums[9][2] [9:0] }), .sum({ \level_6_sums[9][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[9][1] [9:0] }),
     .b({ \level_6_sums[9][0] [9:0] }), .sum({ \level_7_sums[9][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[129] [4:0] }), .sum({ \level_1_sums[9][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[131] [4:0] }), .sum({ \level_1_sums[9][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[9][65] [5:0] }),
     .b({ \level_1_sums[9][64] [5:0] }), .sum({ \level_2_sums[9][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[133] [4:0] }), .sum({ \level_1_sums[9][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[135] [4:0] }), .sum({ \level_1_sums[9][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[9][67] [5:0] }),
     .b({ \level_1_sums[9][66] [5:0] }), .sum({ \level_2_sums[9][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[135].adder_octets.adder_inst (.a({ \level_2_sums[9][33] [6:0] }),
     .b({ \level_2_sums[9][32] [6:0] }), .sum({ \level_3_sums[9][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[137] [4:0] }), .sum({ \level_1_sums[9][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[139] [4:0] }), .sum({ \level_1_sums[9][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[9][69] [5:0] }),
     .b({ \level_1_sums[9][68] [5:0] }), .sum({ \level_2_sums[9][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[141] [4:0] }), .sum({ \level_1_sums[9][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[143] [4:0] }), .sum({ \level_1_sums[9][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[9][71] [5:0] }),
     .b({ \level_1_sums[9][70] [5:0] }), .sum({ \level_2_sums[9][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[143].adder_octets.adder_inst (.a({ \level_2_sums[9][35] [6:0] }),
     .b({ \level_2_sums[9][34] [6:0] }), .sum({ \level_3_sums[9][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[9][17] [7:0] }),
     .b({ \level_3_sums[9][16] [7:0] }), .sum({ \level_4_sums[9][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[145] [4:0] }), .sum({ \level_1_sums[9][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[147] [4:0] }), .sum({ \level_1_sums[9][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[9][73] [5:0] }),
     .b({ \level_1_sums[9][72] [5:0] }), .sum({ \level_2_sums[9][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[149] [4:0] }), .sum({ \level_1_sums[9][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[151] [4:0] }), .sum({ \level_1_sums[9][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[9][75] [5:0] }),
     .b({ \level_1_sums[9][74] [5:0] }), .sum({ \level_2_sums[9][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[151].adder_octets.adder_inst (.a({ \level_2_sums[9][37] [6:0] }),
     .b({ \level_2_sums[9][36] [6:0] }), .sum({ \level_3_sums[9][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[153] [4:0] }), .sum({ \level_1_sums[9][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[155] [4:0] }), .sum({ \level_1_sums[9][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[9][77] [5:0] }),
     .b({ \level_1_sums[9][76] [5:0] }), .sum({ \level_2_sums[9][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[157] [4:0] }), .sum({ \level_1_sums[9][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[159] [4:0] }), .sum({ \level_1_sums[9][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[9][79] [5:0] }),
     .b({ \level_1_sums[9][78] [5:0] }), .sum({ \level_2_sums[9][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[159].adder_octets.adder_inst (.a({ \level_2_sums[9][39] [6:0] }),
     .b({ \level_2_sums[9][38] [6:0] }), .sum({ \level_3_sums[9][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[9][19] [7:0] }),
     .b({ \level_3_sums[9][18] [7:0] }), .sum({ \level_4_sums[9][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[9][9] [8:0] }),
     .b({ \level_4_sums[9][8] [8:0] }), .sum({ \level_5_sums[9][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[161] [4:0] }), .sum({ \level_1_sums[9][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[163] [4:0] }), .sum({ \level_1_sums[9][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[9][81] [5:0] }),
     .b({ \level_1_sums[9][80] [5:0] }), .sum({ \level_2_sums[9][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[165] [4:0] }), .sum({ \level_1_sums[9][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[167] [4:0] }), .sum({ \level_1_sums[9][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[9][83] [5:0] }),
     .b({ \level_1_sums[9][82] [5:0] }), .sum({ \level_2_sums[9][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[167].adder_octets.adder_inst (.a({ \level_2_sums[9][41] [6:0] }),
     .b({ \level_2_sums[9][40] [6:0] }), .sum({ \level_3_sums[9][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[169] [4:0] }), .sum({ \level_1_sums[9][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[171] [4:0] }), .sum({ \level_1_sums[9][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[9][85] [5:0] }),
     .b({ \level_1_sums[9][84] [5:0] }), .sum({ \level_2_sums[9][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[173] [4:0] }), .sum({ \level_1_sums[9][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[175] [4:0] }), .sum({ \level_1_sums[9][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[9][87] [5:0] }),
     .b({ \level_1_sums[9][86] [5:0] }), .sum({ \level_2_sums[9][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[175].adder_octets.adder_inst (.a({ \level_2_sums[9][43] [6:0] }),
     .b({ \level_2_sums[9][42] [6:0] }), .sum({ \level_3_sums[9][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[9][21] [7:0] }),
     .b({ \level_3_sums[9][20] [7:0] }), .sum({ \level_4_sums[9][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[177] [4:0] }), .sum({ \level_1_sums[9][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[179] [4:0] }), .sum({ \level_1_sums[9][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[9][89] [5:0] }),
     .b({ \level_1_sums[9][88] [5:0] }), .sum({ \level_2_sums[9][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[181] [4:0] }), .sum({ \level_1_sums[9][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[183] [4:0] }), .sum({ \level_1_sums[9][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[9][91] [5:0] }),
     .b({ \level_1_sums[9][90] [5:0] }), .sum({ \level_2_sums[9][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[183].adder_octets.adder_inst (.a({ \level_2_sums[9][45] [6:0] }),
     .b({ \level_2_sums[9][44] [6:0] }), .sum({ \level_3_sums[9][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[185] [4:0] }), .sum({ \level_1_sums[9][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[187] [4:0] }), .sum({ \level_1_sums[9][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[9][93] [5:0] }),
     .b({ \level_1_sums[9][92] [5:0] }), .sum({ \level_2_sums[9][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[189] [4:0] }), .sum({ \level_1_sums[9][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[191] [4:0] }), .sum({ \level_1_sums[9][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[9][95] [5:0] }),
     .b({ \level_1_sums[9][94] [5:0] }), .sum({ \level_2_sums[9][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_octets.adder_inst (.a({ \level_2_sums[9][47] [6:0] }),
     .b({ \level_2_sums[9][46] [6:0] }), .sum({ \level_3_sums[9][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[9][23] [7:0] }),
     .b({ \level_3_sums[9][22] [7:0] }), .sum({ \level_4_sums[9][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[9][11] [8:0] }),
     .b({ \level_4_sums[9][10] [8:0] }), .sum({ \level_5_sums[9][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[9][5] [9:0] }),
     .b({ \level_5_sums[9][4] [9:0] }), .sum({ \level_6_sums[9][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[193] [4:0] }), .sum({ \level_1_sums[9][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[195] [4:0] }), .sum({ \level_1_sums[9][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[9][97] [5:0] }),
     .b({ \level_1_sums[9][96] [5:0] }), .sum({ \level_2_sums[9][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[197] [4:0] }), .sum({ \level_1_sums[9][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[199] [4:0] }), .sum({ \level_1_sums[9][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[9][99] [5:0] }),
     .b({ \level_1_sums[9][98] [5:0] }), .sum({ \level_2_sums[9][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[199].adder_octets.adder_inst (.a({ \level_2_sums[9][49] [6:0] }),
     .b({ \level_2_sums[9][48] [6:0] }), .sum({ \level_3_sums[9][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[201] [4:0] }), .sum({ \level_1_sums[9][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[203] [4:0] }), .sum({ \level_1_sums[9][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[9][101] [5:0] }),
     .b({ \level_1_sums[9][100] [5:0] }), .sum({ \level_2_sums[9][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[205] [4:0] }), .sum({ \level_1_sums[9][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[207] [4:0] }), .sum({ \level_1_sums[9][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[9][103] [5:0] }),
     .b({ \level_1_sums[9][102] [5:0] }), .sum({ \level_2_sums[9][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[207].adder_octets.adder_inst (.a({ \level_2_sums[9][51] [6:0] }),
     .b({ \level_2_sums[9][50] [6:0] }), .sum({ \level_3_sums[9][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[9][25] [7:0] }),
     .b({ \level_3_sums[9][24] [7:0] }), .sum({ \level_4_sums[9][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[209] [4:0] }), .sum({ \level_1_sums[9][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[211] [4:0] }), .sum({ \level_1_sums[9][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[9][105] [5:0] }),
     .b({ \level_1_sums[9][104] [5:0] }), .sum({ \level_2_sums[9][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[213] [4:0] }), .sum({ \level_1_sums[9][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[215] [4:0] }), .sum({ \level_1_sums[9][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[9][107] [5:0] }),
     .b({ \level_1_sums[9][106] [5:0] }), .sum({ \level_2_sums[9][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[215].adder_octets.adder_inst (.a({ \level_2_sums[9][53] [6:0] }),
     .b({ \level_2_sums[9][52] [6:0] }), .sum({ \level_3_sums[9][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[217] [4:0] }), .sum({ \level_1_sums[9][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[219] [4:0] }), .sum({ \level_1_sums[9][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[9][109] [5:0] }),
     .b({ \level_1_sums[9][108] [5:0] }), .sum({ \level_2_sums[9][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[221] [4:0] }), .sum({ \level_1_sums[9][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[223] [4:0] }), .sum({ \level_1_sums[9][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[9][111] [5:0] }),
     .b({ \level_1_sums[9][110] [5:0] }), .sum({ \level_2_sums[9][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[223].adder_octets.adder_inst (.a({ \level_2_sums[9][55] [6:0] }),
     .b({ \level_2_sums[9][54] [6:0] }), .sum({ \level_3_sums[9][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[9][27] [7:0] }),
     .b({ \level_3_sums[9][26] [7:0] }), .sum({ \level_4_sums[9][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[9][13] [8:0] }),
     .b({ \level_4_sums[9][12] [8:0] }), .sum({ \level_5_sums[9][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[225] [4:0] }), .sum({ \level_1_sums[9][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[227] [4:0] }), .sum({ \level_1_sums[9][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[9][113] [5:0] }),
     .b({ \level_1_sums[9][112] [5:0] }), .sum({ \level_2_sums[9][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[229] [4:0] }), .sum({ \level_1_sums[9][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[231] [4:0] }), .sum({ \level_1_sums[9][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[9][115] [5:0] }),
     .b({ \level_1_sums[9][114] [5:0] }), .sum({ \level_2_sums[9][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[231].adder_octets.adder_inst (.a({ \level_2_sums[9][57] [6:0] }),
     .b({ \level_2_sums[9][56] [6:0] }), .sum({ \level_3_sums[9][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[233] [4:0] }), .sum({ \level_1_sums[9][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[235] [4:0] }), .sum({ \level_1_sums[9][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[9][117] [5:0] }),
     .b({ \level_1_sums[9][116] [5:0] }), .sum({ \level_2_sums[9][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[237] [4:0] }), .sum({ \level_1_sums[9][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[239] [4:0] }), .sum({ \level_1_sums[9][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[9][119] [5:0] }),
     .b({ \level_1_sums[9][118] [5:0] }), .sum({ \level_2_sums[9][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[239].adder_octets.adder_inst (.a({ \level_2_sums[9][59] [6:0] }),
     .b({ \level_2_sums[9][58] [6:0] }), .sum({ \level_3_sums[9][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[9][29] [7:0] }),
     .b({ \level_3_sums[9][28] [7:0] }), .sum({ \level_4_sums[9][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[241] [4:0] }), .sum({ \level_1_sums[9][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[243] [4:0] }), .sum({ \level_1_sums[9][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[9][121] [5:0] }),
     .b({ \level_1_sums[9][120] [5:0] }), .sum({ \level_2_sums[9][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[245] [4:0] }), .sum({ \level_1_sums[9][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[247] [4:0] }), .sum({ \level_1_sums[9][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[9][123] [5:0] }),
     .b({ \level_1_sums[9][122] [5:0] }), .sum({ \level_2_sums[9][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[247].adder_octets.adder_inst (.a({ \level_2_sums[9][61] [6:0] }),
     .b({ \level_2_sums[9][60] [6:0] }), .sum({ \level_3_sums[9][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[249] [4:0] }), .sum({ \level_1_sums[9][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[251] [4:0] }), .sum({ \level_1_sums[9][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[9][125] [5:0] }),
     .b({ \level_1_sums[9][124] [5:0] }), .sum({ \level_2_sums[9][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[253] [4:0] }), .sum({ \level_1_sums[9][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[9].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[9].product_terms[255] [4:0] }), .sum({ \level_1_sums[9][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[9][127] [5:0] }),
     .b({ \level_1_sums[9][126] [5:0] }), .sum({ \level_2_sums[9][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_octets.adder_inst (.a({ \level_2_sums[9][63] [6:0] }),
     .b({ \level_2_sums[9][62] [6:0] }), .sum({ \level_3_sums[9][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[9][31] [7:0] }),
     .b({ \level_3_sums[9][30] [7:0] }), .sum({ \level_4_sums[9][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[9][15] [8:0] }),
     .b({ \level_4_sums[9][14] [8:0] }), .sum({ \level_5_sums[9][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[9][7] [9:0] }),
     .b({ \level_5_sums[9][6] [9:0] }), .sum({ \level_6_sums[9][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[9][3] [9:0] }),
     .b({ \level_6_sums[9][2] [9:0] }), .sum({ \level_7_sums[9][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[9].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[9][0] [9:0] }),
     .b({ \level_7_sums[9][1] [9:0] }), .sum({ \level_8_sums[9] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[10].relu_inst (.in_data({ \final_sums[10] [9:0] }), .out_data({ \out_sig[10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[1] [4:0] }), .sum({ \level_1_sums[10][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[3] [4:0] }), .sum({ \level_1_sums[10][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[10][1] [5:0] }),
     .b({ \level_1_sums[10][0] [5:0] }), .sum({ \level_2_sums[10][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[5] [4:0] }), .sum({ \level_1_sums[10][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[7] [4:0] }), .sum({ \level_1_sums[10][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[10][3] [5:0] }),
     .b({ \level_1_sums[10][2] [5:0] }), .sum({ \level_2_sums[10][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[10][1] [6:0] }),
     .b({ \level_2_sums[10][0] [6:0] }), .sum({ \level_3_sums[10][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[9] [4:0] }), .sum({ \level_1_sums[10][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[11] [4:0] }), .sum({ \level_1_sums[10][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[10][5] [5:0] }),
     .b({ \level_1_sums[10][4] [5:0] }), .sum({ \level_2_sums[10][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[13] [4:0] }), .sum({ \level_1_sums[10][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[15] [4:0] }), .sum({ \level_1_sums[10][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[10][7] [5:0] }),
     .b({ \level_1_sums[10][6] [5:0] }), .sum({ \level_2_sums[10][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[10][3] [6:0] }),
     .b({ \level_2_sums[10][2] [6:0] }), .sum({ \level_3_sums[10][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[10][1] [7:0] }),
     .b({ \level_3_sums[10][0] [7:0] }), .sum({ \level_4_sums[10][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[17] [4:0] }), .sum({ \level_1_sums[10][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[19] [4:0] }), .sum({ \level_1_sums[10][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[10][9] [5:0] }),
     .b({ \level_1_sums[10][8] [5:0] }), .sum({ \level_2_sums[10][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[21] [4:0] }), .sum({ \level_1_sums[10][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[23] [4:0] }), .sum({ \level_1_sums[10][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[10][11] [5:0] }),
     .b({ \level_1_sums[10][10] [5:0] }), .sum({ \level_2_sums[10][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[10][5] [6:0] }),
     .b({ \level_2_sums[10][4] [6:0] }), .sum({ \level_3_sums[10][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[25] [4:0] }), .sum({ \level_1_sums[10][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[27] [4:0] }), .sum({ \level_1_sums[10][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[10][13] [5:0] }),
     .b({ \level_1_sums[10][12] [5:0] }), .sum({ \level_2_sums[10][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[29] [4:0] }), .sum({ \level_1_sums[10][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[31] [4:0] }), .sum({ \level_1_sums[10][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[10][15] [5:0] }),
     .b({ \level_1_sums[10][14] [5:0] }), .sum({ \level_2_sums[10][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[10][7] [6:0] }),
     .b({ \level_2_sums[10][6] [6:0] }), .sum({ \level_3_sums[10][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[10][3] [7:0] }),
     .b({ \level_3_sums[10][2] [7:0] }), .sum({ \level_4_sums[10][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[10][1] [8:0] }),
     .b({ \level_4_sums[10][0] [8:0] }), .sum({ \level_5_sums[10][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[33] [4:0] }), .sum({ \level_1_sums[10][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[35] [4:0] }), .sum({ \level_1_sums[10][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[10][17] [5:0] }),
     .b({ \level_1_sums[10][16] [5:0] }), .sum({ \level_2_sums[10][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[37] [4:0] }), .sum({ \level_1_sums[10][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[39] [4:0] }), .sum({ \level_1_sums[10][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[10][19] [5:0] }),
     .b({ \level_1_sums[10][18] [5:0] }), .sum({ \level_2_sums[10][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[10][9] [6:0] }),
     .b({ \level_2_sums[10][8] [6:0] }), .sum({ \level_3_sums[10][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[41] [4:0] }), .sum({ \level_1_sums[10][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[43] [4:0] }), .sum({ \level_1_sums[10][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[10][21] [5:0] }),
     .b({ \level_1_sums[10][20] [5:0] }), .sum({ \level_2_sums[10][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[45] [4:0] }), .sum({ \level_1_sums[10][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[47] [4:0] }), .sum({ \level_1_sums[10][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[10][23] [5:0] }),
     .b({ \level_1_sums[10][22] [5:0] }), .sum({ \level_2_sums[10][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[10][11] [6:0] }),
     .b({ \level_2_sums[10][10] [6:0] }), .sum({ \level_3_sums[10][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[10][5] [7:0] }),
     .b({ \level_3_sums[10][4] [7:0] }), .sum({ \level_4_sums[10][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[49] [4:0] }), .sum({ \level_1_sums[10][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[51] [4:0] }), .sum({ \level_1_sums[10][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[10][25] [5:0] }),
     .b({ \level_1_sums[10][24] [5:0] }), .sum({ \level_2_sums[10][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[53] [4:0] }), .sum({ \level_1_sums[10][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[55] [4:0] }), .sum({ \level_1_sums[10][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[10][27] [5:0] }),
     .b({ \level_1_sums[10][26] [5:0] }), .sum({ \level_2_sums[10][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[10][13] [6:0] }),
     .b({ \level_2_sums[10][12] [6:0] }), .sum({ \level_3_sums[10][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[57] [4:0] }), .sum({ \level_1_sums[10][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[59] [4:0] }), .sum({ \level_1_sums[10][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[10][29] [5:0] }),
     .b({ \level_1_sums[10][28] [5:0] }), .sum({ \level_2_sums[10][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[61] [4:0] }), .sum({ \level_1_sums[10][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[63] [4:0] }), .sum({ \level_1_sums[10][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[10][31] [5:0] }),
     .b({ \level_1_sums[10][30] [5:0] }), .sum({ \level_2_sums[10][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[10][15] [6:0] }),
     .b({ \level_2_sums[10][14] [6:0] }), .sum({ \level_3_sums[10][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[10][7] [7:0] }),
     .b({ \level_3_sums[10][6] [7:0] }), .sum({ \level_4_sums[10][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[10][3] [8:0] }),
     .b({ \level_4_sums[10][2] [8:0] }), .sum({ \level_5_sums[10][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[10][1] [9:0] }),
     .b({ \level_5_sums[10][0] [9:0] }), .sum({ \level_6_sums[10][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[65] [4:0] }), .sum({ \level_1_sums[10][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[67] [4:0] }), .sum({ \level_1_sums[10][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[10][33] [5:0] }),
     .b({ \level_1_sums[10][32] [5:0] }), .sum({ \level_2_sums[10][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[69] [4:0] }), .sum({ \level_1_sums[10][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[71] [4:0] }), .sum({ \level_1_sums[10][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[10][35] [5:0] }),
     .b({ \level_1_sums[10][34] [5:0] }), .sum({ \level_2_sums[10][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[10][17] [6:0] }),
     .b({ \level_2_sums[10][16] [6:0] }), .sum({ \level_3_sums[10][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[73] [4:0] }), .sum({ \level_1_sums[10][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[75] [4:0] }), .sum({ \level_1_sums[10][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[10][37] [5:0] }),
     .b({ \level_1_sums[10][36] [5:0] }), .sum({ \level_2_sums[10][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[77] [4:0] }), .sum({ \level_1_sums[10][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[79] [4:0] }), .sum({ \level_1_sums[10][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[10][39] [5:0] }),
     .b({ \level_1_sums[10][38] [5:0] }), .sum({ \level_2_sums[10][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[10][19] [6:0] }),
     .b({ \level_2_sums[10][18] [6:0] }), .sum({ \level_3_sums[10][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[10][9] [7:0] }),
     .b({ \level_3_sums[10][8] [7:0] }), .sum({ \level_4_sums[10][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[81] [4:0] }), .sum({ \level_1_sums[10][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[83] [4:0] }), .sum({ \level_1_sums[10][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[10][41] [5:0] }),
     .b({ \level_1_sums[10][40] [5:0] }), .sum({ \level_2_sums[10][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[85] [4:0] }), .sum({ \level_1_sums[10][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[87] [4:0] }), .sum({ \level_1_sums[10][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[10][43] [5:0] }),
     .b({ \level_1_sums[10][42] [5:0] }), .sum({ \level_2_sums[10][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[10][21] [6:0] }),
     .b({ \level_2_sums[10][20] [6:0] }), .sum({ \level_3_sums[10][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[89] [4:0] }), .sum({ \level_1_sums[10][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[91] [4:0] }), .sum({ \level_1_sums[10][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[10][45] [5:0] }),
     .b({ \level_1_sums[10][44] [5:0] }), .sum({ \level_2_sums[10][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[93] [4:0] }), .sum({ \level_1_sums[10][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[95] [4:0] }), .sum({ \level_1_sums[10][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[10][47] [5:0] }),
     .b({ \level_1_sums[10][46] [5:0] }), .sum({ \level_2_sums[10][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[10][23] [6:0] }),
     .b({ \level_2_sums[10][22] [6:0] }), .sum({ \level_3_sums[10][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[10][11] [7:0] }),
     .b({ \level_3_sums[10][10] [7:0] }), .sum({ \level_4_sums[10][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[10][5] [8:0] }),
     .b({ \level_4_sums[10][4] [8:0] }), .sum({ \level_5_sums[10][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[97] [4:0] }), .sum({ \level_1_sums[10][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[99] [4:0] }), .sum({ \level_1_sums[10][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[10][49] [5:0] }),
     .b({ \level_1_sums[10][48] [5:0] }), .sum({ \level_2_sums[10][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[101] [4:0] }), .sum({ \level_1_sums[10][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[103] [4:0] }), .sum({ \level_1_sums[10][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[10][51] [5:0] }),
     .b({ \level_1_sums[10][50] [5:0] }), .sum({ \level_2_sums[10][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[10][25] [6:0] }), .b({ \level_2_sums[10][24] [6:0] }), .sum({ \level_3_sums[10][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[105] [4:0] }), .sum({ \level_1_sums[10][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[107] [4:0] }), .sum({ \level_1_sums[10][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[10][53] [5:0] }),
     .b({ \level_1_sums[10][52] [5:0] }), .sum({ \level_2_sums[10][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[109] [4:0] }), .sum({ \level_1_sums[10][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[111] [4:0] }), .sum({ \level_1_sums[10][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[10][55] [5:0] }),
     .b({ \level_1_sums[10][54] [5:0] }), .sum({ \level_2_sums[10][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[10][27] [6:0] }), .b({ \level_2_sums[10][26] [6:0] }), .sum({ \level_3_sums[10][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[10][13] [7:0] }),
     .b({ \level_3_sums[10][12] [7:0] }), .sum({ \level_4_sums[10][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[113] [4:0] }), .sum({ \level_1_sums[10][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[115] [4:0] }), .sum({ \level_1_sums[10][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[10][57] [5:0] }),
     .b({ \level_1_sums[10][56] [5:0] }), .sum({ \level_2_sums[10][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[117] [4:0] }), .sum({ \level_1_sums[10][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[119] [4:0] }), .sum({ \level_1_sums[10][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[10][59] [5:0] }),
     .b({ \level_1_sums[10][58] [5:0] }), .sum({ \level_2_sums[10][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[10][29] [6:0] }), .b({ \level_2_sums[10][28] [6:0] }), .sum({ \level_3_sums[10][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[121] [4:0] }), .sum({ \level_1_sums[10][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[123] [4:0] }), .sum({ \level_1_sums[10][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[10][61] [5:0] }),
     .b({ \level_1_sums[10][60] [5:0] }), .sum({ \level_2_sums[10][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[125] [4:0] }), .sum({ \level_1_sums[10][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[127] [4:0] }), .sum({ \level_1_sums[10][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[10][63] [5:0] }),
     .b({ \level_1_sums[10][62] [5:0] }), .sum({ \level_2_sums[10][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[10][31] [6:0] }), .b({ \level_2_sums[10][30] [6:0] }), .sum({ \level_3_sums[10][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[10][15] [7:0] }),
     .b({ \level_3_sums[10][14] [7:0] }), .sum({ \level_4_sums[10][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[10][7] [8:0] }),
     .b({ \level_4_sums[10][6] [8:0] }), .sum({ \level_5_sums[10][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[10][3] [9:0] }),
     .b({ \level_5_sums[10][2] [9:0] }), .sum({ \level_6_sums[10][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[10][1] [9:0] }),
     .b({ \level_6_sums[10][0] [9:0] }), .sum({ \level_7_sums[10][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[129] [4:0] }), .sum({ \level_1_sums[10][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[131] [4:0] }), .sum({ \level_1_sums[10][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[10][65] [5:0] }),
     .b({ \level_1_sums[10][64] [5:0] }), .sum({ \level_2_sums[10][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[133] [4:0] }), .sum({ \level_1_sums[10][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[135] [4:0] }), .sum({ \level_1_sums[10][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[10][67] [5:0] }),
     .b({ \level_1_sums[10][66] [5:0] }), .sum({ \level_2_sums[10][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[10][33] [6:0] }), .b({ \level_2_sums[10][32] [6:0] }), .sum({ \level_3_sums[10][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[137] [4:0] }), .sum({ \level_1_sums[10][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[139] [4:0] }), .sum({ \level_1_sums[10][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[10][69] [5:0] }),
     .b({ \level_1_sums[10][68] [5:0] }), .sum({ \level_2_sums[10][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[141] [4:0] }), .sum({ \level_1_sums[10][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[143] [4:0] }), .sum({ \level_1_sums[10][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[10][71] [5:0] }),
     .b({ \level_1_sums[10][70] [5:0] }), .sum({ \level_2_sums[10][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[10][35] [6:0] }), .b({ \level_2_sums[10][34] [6:0] }), .sum({ \level_3_sums[10][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[10][17] [7:0] }),
     .b({ \level_3_sums[10][16] [7:0] }), .sum({ \level_4_sums[10][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[145] [4:0] }), .sum({ \level_1_sums[10][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[147] [4:0] }), .sum({ \level_1_sums[10][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[10][73] [5:0] }),
     .b({ \level_1_sums[10][72] [5:0] }), .sum({ \level_2_sums[10][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[149] [4:0] }), .sum({ \level_1_sums[10][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[151] [4:0] }), .sum({ \level_1_sums[10][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[10][75] [5:0] }),
     .b({ \level_1_sums[10][74] [5:0] }), .sum({ \level_2_sums[10][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[10][37] [6:0] }), .b({ \level_2_sums[10][36] [6:0] }), .sum({ \level_3_sums[10][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[153] [4:0] }), .sum({ \level_1_sums[10][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[155] [4:0] }), .sum({ \level_1_sums[10][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[10][77] [5:0] }),
     .b({ \level_1_sums[10][76] [5:0] }), .sum({ \level_2_sums[10][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[157] [4:0] }), .sum({ \level_1_sums[10][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[159] [4:0] }), .sum({ \level_1_sums[10][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[10][79] [5:0] }),
     .b({ \level_1_sums[10][78] [5:0] }), .sum({ \level_2_sums[10][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[10][39] [6:0] }), .b({ \level_2_sums[10][38] [6:0] }), .sum({ \level_3_sums[10][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[10][19] [7:0] }),
     .b({ \level_3_sums[10][18] [7:0] }), .sum({ \level_4_sums[10][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[10][9] [8:0] }),
     .b({ \level_4_sums[10][8] [8:0] }), .sum({ \level_5_sums[10][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[161] [4:0] }), .sum({ \level_1_sums[10][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[163] [4:0] }), .sum({ \level_1_sums[10][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[10][81] [5:0] }),
     .b({ \level_1_sums[10][80] [5:0] }), .sum({ \level_2_sums[10][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[165] [4:0] }), .sum({ \level_1_sums[10][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[167] [4:0] }), .sum({ \level_1_sums[10][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[10][83] [5:0] }),
     .b({ \level_1_sums[10][82] [5:0] }), .sum({ \level_2_sums[10][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[10][41] [6:0] }), .b({ \level_2_sums[10][40] [6:0] }), .sum({ \level_3_sums[10][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[169] [4:0] }), .sum({ \level_1_sums[10][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[171] [4:0] }), .sum({ \level_1_sums[10][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[10][85] [5:0] }),
     .b({ \level_1_sums[10][84] [5:0] }), .sum({ \level_2_sums[10][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[173] [4:0] }), .sum({ \level_1_sums[10][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[175] [4:0] }), .sum({ \level_1_sums[10][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[10][87] [5:0] }),
     .b({ \level_1_sums[10][86] [5:0] }), .sum({ \level_2_sums[10][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[10][43] [6:0] }), .b({ \level_2_sums[10][42] [6:0] }), .sum({ \level_3_sums[10][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[10][21] [7:0] }),
     .b({ \level_3_sums[10][20] [7:0] }), .sum({ \level_4_sums[10][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[177] [4:0] }), .sum({ \level_1_sums[10][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[179] [4:0] }), .sum({ \level_1_sums[10][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[10][89] [5:0] }),
     .b({ \level_1_sums[10][88] [5:0] }), .sum({ \level_2_sums[10][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[181] [4:0] }), .sum({ \level_1_sums[10][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[183] [4:0] }), .sum({ \level_1_sums[10][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[10][91] [5:0] }),
     .b({ \level_1_sums[10][90] [5:0] }), .sum({ \level_2_sums[10][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[10][45] [6:0] }), .b({ \level_2_sums[10][44] [6:0] }), .sum({ \level_3_sums[10][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[185] [4:0] }), .sum({ \level_1_sums[10][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[187] [4:0] }), .sum({ \level_1_sums[10][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[10][93] [5:0] }),
     .b({ \level_1_sums[10][92] [5:0] }), .sum({ \level_2_sums[10][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[189] [4:0] }), .sum({ \level_1_sums[10][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[191] [4:0] }), .sum({ \level_1_sums[10][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[10][95] [5:0] }),
     .b({ \level_1_sums[10][94] [5:0] }), .sum({ \level_2_sums[10][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[10][47] [6:0] }), .b({ \level_2_sums[10][46] [6:0] }), .sum({ \level_3_sums[10][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[10][23] [7:0] }),
     .b({ \level_3_sums[10][22] [7:0] }), .sum({ \level_4_sums[10][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[10][11] [8:0] }),
     .b({ \level_4_sums[10][10] [8:0] }), .sum({ \level_5_sums[10][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[10][5] [9:0] }),
     .b({ \level_5_sums[10][4] [9:0] }), .sum({ \level_6_sums[10][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[193] [4:0] }), .sum({ \level_1_sums[10][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[195] [4:0] }), .sum({ \level_1_sums[10][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[10][97] [5:0] }),
     .b({ \level_1_sums[10][96] [5:0] }), .sum({ \level_2_sums[10][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[197] [4:0] }), .sum({ \level_1_sums[10][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[199] [4:0] }), .sum({ \level_1_sums[10][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[10][99] [5:0] }),
     .b({ \level_1_sums[10][98] [5:0] }), .sum({ \level_2_sums[10][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[10][49] [6:0] }), .b({ \level_2_sums[10][48] [6:0] }), .sum({ \level_3_sums[10][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[201] [4:0] }), .sum({ \level_1_sums[10][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[203] [4:0] }), .sum({ \level_1_sums[10][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[10][101] [5:0] }),
     .b({ \level_1_sums[10][100] [5:0] }), .sum({ \level_2_sums[10][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[205] [4:0] }), .sum({ \level_1_sums[10][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[207] [4:0] }), .sum({ \level_1_sums[10][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[10][103] [5:0] }),
     .b({ \level_1_sums[10][102] [5:0] }), .sum({ \level_2_sums[10][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[10][51] [6:0] }), .b({ \level_2_sums[10][50] [6:0] }), .sum({ \level_3_sums[10][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[10][25] [7:0] }),
     .b({ \level_3_sums[10][24] [7:0] }), .sum({ \level_4_sums[10][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[209] [4:0] }), .sum({ \level_1_sums[10][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[211] [4:0] }), .sum({ \level_1_sums[10][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[10][105] [5:0] }),
     .b({ \level_1_sums[10][104] [5:0] }), .sum({ \level_2_sums[10][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[213] [4:0] }), .sum({ \level_1_sums[10][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[215] [4:0] }), .sum({ \level_1_sums[10][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[10][107] [5:0] }),
     .b({ \level_1_sums[10][106] [5:0] }), .sum({ \level_2_sums[10][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[10][53] [6:0] }), .b({ \level_2_sums[10][52] [6:0] }), .sum({ \level_3_sums[10][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[217] [4:0] }), .sum({ \level_1_sums[10][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[219] [4:0] }), .sum({ \level_1_sums[10][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[10][109] [5:0] }),
     .b({ \level_1_sums[10][108] [5:0] }), .sum({ \level_2_sums[10][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[221] [4:0] }), .sum({ \level_1_sums[10][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[223] [4:0] }), .sum({ \level_1_sums[10][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[10][111] [5:0] }),
     .b({ \level_1_sums[10][110] [5:0] }), .sum({ \level_2_sums[10][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[10][55] [6:0] }), .b({ \level_2_sums[10][54] [6:0] }), .sum({ \level_3_sums[10][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[10][27] [7:0] }),
     .b({ \level_3_sums[10][26] [7:0] }), .sum({ \level_4_sums[10][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[10][13] [8:0] }),
     .b({ \level_4_sums[10][12] [8:0] }), .sum({ \level_5_sums[10][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[225] [4:0] }), .sum({ \level_1_sums[10][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[227] [4:0] }), .sum({ \level_1_sums[10][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[10][113] [5:0] }),
     .b({ \level_1_sums[10][112] [5:0] }), .sum({ \level_2_sums[10][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[229] [4:0] }), .sum({ \level_1_sums[10][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[231] [4:0] }), .sum({ \level_1_sums[10][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[10][115] [5:0] }),
     .b({ \level_1_sums[10][114] [5:0] }), .sum({ \level_2_sums[10][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[10][57] [6:0] }), .b({ \level_2_sums[10][56] [6:0] }), .sum({ \level_3_sums[10][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[233] [4:0] }), .sum({ \level_1_sums[10][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[235] [4:0] }), .sum({ \level_1_sums[10][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[10][117] [5:0] }),
     .b({ \level_1_sums[10][116] [5:0] }), .sum({ \level_2_sums[10][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[237] [4:0] }), .sum({ \level_1_sums[10][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[239] [4:0] }), .sum({ \level_1_sums[10][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[10][119] [5:0] }),
     .b({ \level_1_sums[10][118] [5:0] }), .sum({ \level_2_sums[10][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[10][59] [6:0] }), .b({ \level_2_sums[10][58] [6:0] }), .sum({ \level_3_sums[10][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[10][29] [7:0] }),
     .b({ \level_3_sums[10][28] [7:0] }), .sum({ \level_4_sums[10][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[241] [4:0] }), .sum({ \level_1_sums[10][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[243] [4:0] }), .sum({ \level_1_sums[10][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[10][121] [5:0] }),
     .b({ \level_1_sums[10][120] [5:0] }), .sum({ \level_2_sums[10][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[245] [4:0] }), .sum({ \level_1_sums[10][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[247] [4:0] }), .sum({ \level_1_sums[10][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[10][123] [5:0] }),
     .b({ \level_1_sums[10][122] [5:0] }), .sum({ \level_2_sums[10][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[10][61] [6:0] }), .b({ \level_2_sums[10][60] [6:0] }), .sum({ \level_3_sums[10][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[249] [4:0] }), .sum({ \level_1_sums[10][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[251] [4:0] }), .sum({ \level_1_sums[10][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[10][125] [5:0] }),
     .b({ \level_1_sums[10][124] [5:0] }), .sum({ \level_2_sums[10][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[253] [4:0] }), .sum({ \level_1_sums[10][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[10].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[10].product_terms[255] [4:0] }), .sum({ \level_1_sums[10][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[10][127] [5:0] }),
     .b({ \level_1_sums[10][126] [5:0] }), .sum({ \level_2_sums[10][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[10][63] [6:0] }), .b({ \level_2_sums[10][62] [6:0] }), .sum({ \level_3_sums[10][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[10][31] [7:0] }),
     .b({ \level_3_sums[10][30] [7:0] }), .sum({ \level_4_sums[10][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[10][15] [8:0] }),
     .b({ \level_4_sums[10][14] [8:0] }), .sum({ \level_5_sums[10][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[10][7] [9:0] }),
     .b({ \level_5_sums[10][6] [9:0] }), .sum({ \level_6_sums[10][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[10][3] [9:0] }),
     .b({ \level_6_sums[10][2] [9:0] }), .sum({ \level_7_sums[10][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[10].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[10][0] [9:0] }),
     .b({ \level_7_sums[10][1] [9:0] }), .sum({ \level_8_sums[10] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[11].relu_inst (.in_data({ \final_sums[11] [9:0] }), .out_data({ \out_sig[11] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[1] [4:0] }), .sum({ \level_1_sums[11][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[3] [4:0] }), .sum({ \level_1_sums[11][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[11][1] [5:0] }),
     .b({ \level_1_sums[11][0] [5:0] }), .sum({ \level_2_sums[11][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[5] [4:0] }), .sum({ \level_1_sums[11][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[7] [4:0] }), .sum({ \level_1_sums[11][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[11][3] [5:0] }),
     .b({ \level_1_sums[11][2] [5:0] }), .sum({ \level_2_sums[11][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[11][1] [6:0] }),
     .b({ \level_2_sums[11][0] [6:0] }), .sum({ \level_3_sums[11][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[9] [4:0] }), .sum({ \level_1_sums[11][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[11] [4:0] }), .sum({ \level_1_sums[11][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[11][5] [5:0] }),
     .b({ \level_1_sums[11][4] [5:0] }), .sum({ \level_2_sums[11][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[13] [4:0] }), .sum({ \level_1_sums[11][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[15] [4:0] }), .sum({ \level_1_sums[11][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[11][7] [5:0] }),
     .b({ \level_1_sums[11][6] [5:0] }), .sum({ \level_2_sums[11][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[11][3] [6:0] }),
     .b({ \level_2_sums[11][2] [6:0] }), .sum({ \level_3_sums[11][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[11][1] [7:0] }),
     .b({ \level_3_sums[11][0] [7:0] }), .sum({ \level_4_sums[11][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[17] [4:0] }), .sum({ \level_1_sums[11][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[19] [4:0] }), .sum({ \level_1_sums[11][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[11][9] [5:0] }),
     .b({ \level_1_sums[11][8] [5:0] }), .sum({ \level_2_sums[11][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[21] [4:0] }), .sum({ \level_1_sums[11][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[23] [4:0] }), .sum({ \level_1_sums[11][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[11][11] [5:0] }),
     .b({ \level_1_sums[11][10] [5:0] }), .sum({ \level_2_sums[11][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[11][5] [6:0] }),
     .b({ \level_2_sums[11][4] [6:0] }), .sum({ \level_3_sums[11][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[25] [4:0] }), .sum({ \level_1_sums[11][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[27] [4:0] }), .sum({ \level_1_sums[11][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[11][13] [5:0] }),
     .b({ \level_1_sums[11][12] [5:0] }), .sum({ \level_2_sums[11][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[29] [4:0] }), .sum({ \level_1_sums[11][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[31] [4:0] }), .sum({ \level_1_sums[11][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[11][15] [5:0] }),
     .b({ \level_1_sums[11][14] [5:0] }), .sum({ \level_2_sums[11][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[11][7] [6:0] }),
     .b({ \level_2_sums[11][6] [6:0] }), .sum({ \level_3_sums[11][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[11][3] [7:0] }),
     .b({ \level_3_sums[11][2] [7:0] }), .sum({ \level_4_sums[11][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[11][1] [8:0] }),
     .b({ \level_4_sums[11][0] [8:0] }), .sum({ \level_5_sums[11][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[33] [4:0] }), .sum({ \level_1_sums[11][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[35] [4:0] }), .sum({ \level_1_sums[11][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[11][17] [5:0] }),
     .b({ \level_1_sums[11][16] [5:0] }), .sum({ \level_2_sums[11][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[37] [4:0] }), .sum({ \level_1_sums[11][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[39] [4:0] }), .sum({ \level_1_sums[11][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[11][19] [5:0] }),
     .b({ \level_1_sums[11][18] [5:0] }), .sum({ \level_2_sums[11][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[11][9] [6:0] }),
     .b({ \level_2_sums[11][8] [6:0] }), .sum({ \level_3_sums[11][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[41] [4:0] }), .sum({ \level_1_sums[11][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[43] [4:0] }), .sum({ \level_1_sums[11][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[11][21] [5:0] }),
     .b({ \level_1_sums[11][20] [5:0] }), .sum({ \level_2_sums[11][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[45] [4:0] }), .sum({ \level_1_sums[11][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[47] [4:0] }), .sum({ \level_1_sums[11][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[11][23] [5:0] }),
     .b({ \level_1_sums[11][22] [5:0] }), .sum({ \level_2_sums[11][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[11][11] [6:0] }),
     .b({ \level_2_sums[11][10] [6:0] }), .sum({ \level_3_sums[11][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[11][5] [7:0] }),
     .b({ \level_3_sums[11][4] [7:0] }), .sum({ \level_4_sums[11][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[49] [4:0] }), .sum({ \level_1_sums[11][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[51] [4:0] }), .sum({ \level_1_sums[11][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[11][25] [5:0] }),
     .b({ \level_1_sums[11][24] [5:0] }), .sum({ \level_2_sums[11][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[53] [4:0] }), .sum({ \level_1_sums[11][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[55] [4:0] }), .sum({ \level_1_sums[11][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[11][27] [5:0] }),
     .b({ \level_1_sums[11][26] [5:0] }), .sum({ \level_2_sums[11][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[11][13] [6:0] }),
     .b({ \level_2_sums[11][12] [6:0] }), .sum({ \level_3_sums[11][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[57] [4:0] }), .sum({ \level_1_sums[11][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[59] [4:0] }), .sum({ \level_1_sums[11][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[11][29] [5:0] }),
     .b({ \level_1_sums[11][28] [5:0] }), .sum({ \level_2_sums[11][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[61] [4:0] }), .sum({ \level_1_sums[11][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[63] [4:0] }), .sum({ \level_1_sums[11][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[11][31] [5:0] }),
     .b({ \level_1_sums[11][30] [5:0] }), .sum({ \level_2_sums[11][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[11][15] [6:0] }),
     .b({ \level_2_sums[11][14] [6:0] }), .sum({ \level_3_sums[11][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[11][7] [7:0] }),
     .b({ \level_3_sums[11][6] [7:0] }), .sum({ \level_4_sums[11][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[11][3] [8:0] }),
     .b({ \level_4_sums[11][2] [8:0] }), .sum({ \level_5_sums[11][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[11][1] [9:0] }),
     .b({ \level_5_sums[11][0] [9:0] }), .sum({ \level_6_sums[11][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[65] [4:0] }), .sum({ \level_1_sums[11][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[67] [4:0] }), .sum({ \level_1_sums[11][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[11][33] [5:0] }),
     .b({ \level_1_sums[11][32] [5:0] }), .sum({ \level_2_sums[11][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[69] [4:0] }), .sum({ \level_1_sums[11][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[71] [4:0] }), .sum({ \level_1_sums[11][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[11][35] [5:0] }),
     .b({ \level_1_sums[11][34] [5:0] }), .sum({ \level_2_sums[11][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[11][17] [6:0] }),
     .b({ \level_2_sums[11][16] [6:0] }), .sum({ \level_3_sums[11][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[73] [4:0] }), .sum({ \level_1_sums[11][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[75] [4:0] }), .sum({ \level_1_sums[11][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[11][37] [5:0] }),
     .b({ \level_1_sums[11][36] [5:0] }), .sum({ \level_2_sums[11][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[77] [4:0] }), .sum({ \level_1_sums[11][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[79] [4:0] }), .sum({ \level_1_sums[11][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[11][39] [5:0] }),
     .b({ \level_1_sums[11][38] [5:0] }), .sum({ \level_2_sums[11][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[11][19] [6:0] }),
     .b({ \level_2_sums[11][18] [6:0] }), .sum({ \level_3_sums[11][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[11][9] [7:0] }),
     .b({ \level_3_sums[11][8] [7:0] }), .sum({ \level_4_sums[11][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[81] [4:0] }), .sum({ \level_1_sums[11][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[83] [4:0] }), .sum({ \level_1_sums[11][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[11][41] [5:0] }),
     .b({ \level_1_sums[11][40] [5:0] }), .sum({ \level_2_sums[11][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[85] [4:0] }), .sum({ \level_1_sums[11][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[87] [4:0] }), .sum({ \level_1_sums[11][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[11][43] [5:0] }),
     .b({ \level_1_sums[11][42] [5:0] }), .sum({ \level_2_sums[11][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[11][21] [6:0] }),
     .b({ \level_2_sums[11][20] [6:0] }), .sum({ \level_3_sums[11][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[89] [4:0] }), .sum({ \level_1_sums[11][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[91] [4:0] }), .sum({ \level_1_sums[11][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[11][45] [5:0] }),
     .b({ \level_1_sums[11][44] [5:0] }), .sum({ \level_2_sums[11][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[93] [4:0] }), .sum({ \level_1_sums[11][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[95] [4:0] }), .sum({ \level_1_sums[11][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[11][47] [5:0] }),
     .b({ \level_1_sums[11][46] [5:0] }), .sum({ \level_2_sums[11][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[11][23] [6:0] }),
     .b({ \level_2_sums[11][22] [6:0] }), .sum({ \level_3_sums[11][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[11][11] [7:0] }),
     .b({ \level_3_sums[11][10] [7:0] }), .sum({ \level_4_sums[11][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[11][5] [8:0] }),
     .b({ \level_4_sums[11][4] [8:0] }), .sum({ \level_5_sums[11][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[97] [4:0] }), .sum({ \level_1_sums[11][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[99] [4:0] }), .sum({ \level_1_sums[11][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[11][49] [5:0] }),
     .b({ \level_1_sums[11][48] [5:0] }), .sum({ \level_2_sums[11][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[101] [4:0] }), .sum({ \level_1_sums[11][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[103] [4:0] }), .sum({ \level_1_sums[11][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[11][51] [5:0] }),
     .b({ \level_1_sums[11][50] [5:0] }), .sum({ \level_2_sums[11][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[11][25] [6:0] }), .b({ \level_2_sums[11][24] [6:0] }), .sum({ \level_3_sums[11][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[105] [4:0] }), .sum({ \level_1_sums[11][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[107] [4:0] }), .sum({ \level_1_sums[11][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[11][53] [5:0] }),
     .b({ \level_1_sums[11][52] [5:0] }), .sum({ \level_2_sums[11][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[109] [4:0] }), .sum({ \level_1_sums[11][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[111] [4:0] }), .sum({ \level_1_sums[11][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[11][55] [5:0] }),
     .b({ \level_1_sums[11][54] [5:0] }), .sum({ \level_2_sums[11][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[11][27] [6:0] }), .b({ \level_2_sums[11][26] [6:0] }), .sum({ \level_3_sums[11][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[11][13] [7:0] }),
     .b({ \level_3_sums[11][12] [7:0] }), .sum({ \level_4_sums[11][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[113] [4:0] }), .sum({ \level_1_sums[11][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[115] [4:0] }), .sum({ \level_1_sums[11][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[11][57] [5:0] }),
     .b({ \level_1_sums[11][56] [5:0] }), .sum({ \level_2_sums[11][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[117] [4:0] }), .sum({ \level_1_sums[11][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[119] [4:0] }), .sum({ \level_1_sums[11][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[11][59] [5:0] }),
     .b({ \level_1_sums[11][58] [5:0] }), .sum({ \level_2_sums[11][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[11][29] [6:0] }), .b({ \level_2_sums[11][28] [6:0] }), .sum({ \level_3_sums[11][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[121] [4:0] }), .sum({ \level_1_sums[11][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[123] [4:0] }), .sum({ \level_1_sums[11][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[11][61] [5:0] }),
     .b({ \level_1_sums[11][60] [5:0] }), .sum({ \level_2_sums[11][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[125] [4:0] }), .sum({ \level_1_sums[11][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[127] [4:0] }), .sum({ \level_1_sums[11][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[11][63] [5:0] }),
     .b({ \level_1_sums[11][62] [5:0] }), .sum({ \level_2_sums[11][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[11][31] [6:0] }), .b({ \level_2_sums[11][30] [6:0] }), .sum({ \level_3_sums[11][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[11][15] [7:0] }),
     .b({ \level_3_sums[11][14] [7:0] }), .sum({ \level_4_sums[11][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[11][7] [8:0] }),
     .b({ \level_4_sums[11][6] [8:0] }), .sum({ \level_5_sums[11][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[11][3] [9:0] }),
     .b({ \level_5_sums[11][2] [9:0] }), .sum({ \level_6_sums[11][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[11][1] [9:0] }),
     .b({ \level_6_sums[11][0] [9:0] }), .sum({ \level_7_sums[11][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[129] [4:0] }), .sum({ \level_1_sums[11][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[131] [4:0] }), .sum({ \level_1_sums[11][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[11][65] [5:0] }),
     .b({ \level_1_sums[11][64] [5:0] }), .sum({ \level_2_sums[11][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[133] [4:0] }), .sum({ \level_1_sums[11][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[135] [4:0] }), .sum({ \level_1_sums[11][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[11][67] [5:0] }),
     .b({ \level_1_sums[11][66] [5:0] }), .sum({ \level_2_sums[11][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[11][33] [6:0] }), .b({ \level_2_sums[11][32] [6:0] }), .sum({ \level_3_sums[11][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[137] [4:0] }), .sum({ \level_1_sums[11][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[139] [4:0] }), .sum({ \level_1_sums[11][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[11][69] [5:0] }),
     .b({ \level_1_sums[11][68] [5:0] }), .sum({ \level_2_sums[11][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[141] [4:0] }), .sum({ \level_1_sums[11][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[143] [4:0] }), .sum({ \level_1_sums[11][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[11][71] [5:0] }),
     .b({ \level_1_sums[11][70] [5:0] }), .sum({ \level_2_sums[11][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[11][35] [6:0] }), .b({ \level_2_sums[11][34] [6:0] }), .sum({ \level_3_sums[11][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[11][17] [7:0] }),
     .b({ \level_3_sums[11][16] [7:0] }), .sum({ \level_4_sums[11][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[145] [4:0] }), .sum({ \level_1_sums[11][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[147] [4:0] }), .sum({ \level_1_sums[11][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[11][73] [5:0] }),
     .b({ \level_1_sums[11][72] [5:0] }), .sum({ \level_2_sums[11][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[149] [4:0] }), .sum({ \level_1_sums[11][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[151] [4:0] }), .sum({ \level_1_sums[11][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[11][75] [5:0] }),
     .b({ \level_1_sums[11][74] [5:0] }), .sum({ \level_2_sums[11][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[11][37] [6:0] }), .b({ \level_2_sums[11][36] [6:0] }), .sum({ \level_3_sums[11][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[153] [4:0] }), .sum({ \level_1_sums[11][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[155] [4:0] }), .sum({ \level_1_sums[11][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[11][77] [5:0] }),
     .b({ \level_1_sums[11][76] [5:0] }), .sum({ \level_2_sums[11][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[157] [4:0] }), .sum({ \level_1_sums[11][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[159] [4:0] }), .sum({ \level_1_sums[11][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[11][79] [5:0] }),
     .b({ \level_1_sums[11][78] [5:0] }), .sum({ \level_2_sums[11][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[11][39] [6:0] }), .b({ \level_2_sums[11][38] [6:0] }), .sum({ \level_3_sums[11][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[11][19] [7:0] }),
     .b({ \level_3_sums[11][18] [7:0] }), .sum({ \level_4_sums[11][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[11][9] [8:0] }),
     .b({ \level_4_sums[11][8] [8:0] }), .sum({ \level_5_sums[11][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[161] [4:0] }), .sum({ \level_1_sums[11][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[163] [4:0] }), .sum({ \level_1_sums[11][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[11][81] [5:0] }),
     .b({ \level_1_sums[11][80] [5:0] }), .sum({ \level_2_sums[11][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[165] [4:0] }), .sum({ \level_1_sums[11][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[167] [4:0] }), .sum({ \level_1_sums[11][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[11][83] [5:0] }),
     .b({ \level_1_sums[11][82] [5:0] }), .sum({ \level_2_sums[11][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[11][41] [6:0] }), .b({ \level_2_sums[11][40] [6:0] }), .sum({ \level_3_sums[11][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[169] [4:0] }), .sum({ \level_1_sums[11][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[171] [4:0] }), .sum({ \level_1_sums[11][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[11][85] [5:0] }),
     .b({ \level_1_sums[11][84] [5:0] }), .sum({ \level_2_sums[11][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[173] [4:0] }), .sum({ \level_1_sums[11][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[175] [4:0] }), .sum({ \level_1_sums[11][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[11][87] [5:0] }),
     .b({ \level_1_sums[11][86] [5:0] }), .sum({ \level_2_sums[11][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[11][43] [6:0] }), .b({ \level_2_sums[11][42] [6:0] }), .sum({ \level_3_sums[11][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[11][21] [7:0] }),
     .b({ \level_3_sums[11][20] [7:0] }), .sum({ \level_4_sums[11][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[177] [4:0] }), .sum({ \level_1_sums[11][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[179] [4:0] }), .sum({ \level_1_sums[11][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[11][89] [5:0] }),
     .b({ \level_1_sums[11][88] [5:0] }), .sum({ \level_2_sums[11][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[181] [4:0] }), .sum({ \level_1_sums[11][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[183] [4:0] }), .sum({ \level_1_sums[11][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[11][91] [5:0] }),
     .b({ \level_1_sums[11][90] [5:0] }), .sum({ \level_2_sums[11][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[11][45] [6:0] }), .b({ \level_2_sums[11][44] [6:0] }), .sum({ \level_3_sums[11][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[185] [4:0] }), .sum({ \level_1_sums[11][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[187] [4:0] }), .sum({ \level_1_sums[11][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[11][93] [5:0] }),
     .b({ \level_1_sums[11][92] [5:0] }), .sum({ \level_2_sums[11][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[189] [4:0] }), .sum({ \level_1_sums[11][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[191] [4:0] }), .sum({ \level_1_sums[11][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[11][95] [5:0] }),
     .b({ \level_1_sums[11][94] [5:0] }), .sum({ \level_2_sums[11][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[11][47] [6:0] }), .b({ \level_2_sums[11][46] [6:0] }), .sum({ \level_3_sums[11][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[11][23] [7:0] }),
     .b({ \level_3_sums[11][22] [7:0] }), .sum({ \level_4_sums[11][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[11][11] [8:0] }),
     .b({ \level_4_sums[11][10] [8:0] }), .sum({ \level_5_sums[11][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[11][5] [9:0] }),
     .b({ \level_5_sums[11][4] [9:0] }), .sum({ \level_6_sums[11][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[193] [4:0] }), .sum({ \level_1_sums[11][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[195] [4:0] }), .sum({ \level_1_sums[11][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[11][97] [5:0] }),
     .b({ \level_1_sums[11][96] [5:0] }), .sum({ \level_2_sums[11][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[197] [4:0] }), .sum({ \level_1_sums[11][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[199] [4:0] }), .sum({ \level_1_sums[11][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[11][99] [5:0] }),
     .b({ \level_1_sums[11][98] [5:0] }), .sum({ \level_2_sums[11][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[11][49] [6:0] }), .b({ \level_2_sums[11][48] [6:0] }), .sum({ \level_3_sums[11][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[201] [4:0] }), .sum({ \level_1_sums[11][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[203] [4:0] }), .sum({ \level_1_sums[11][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[11][101] [5:0] }),
     .b({ \level_1_sums[11][100] [5:0] }), .sum({ \level_2_sums[11][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[205] [4:0] }), .sum({ \level_1_sums[11][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[207] [4:0] }), .sum({ \level_1_sums[11][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[11][103] [5:0] }),
     .b({ \level_1_sums[11][102] [5:0] }), .sum({ \level_2_sums[11][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[11][51] [6:0] }), .b({ \level_2_sums[11][50] [6:0] }), .sum({ \level_3_sums[11][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[11][25] [7:0] }),
     .b({ \level_3_sums[11][24] [7:0] }), .sum({ \level_4_sums[11][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[209] [4:0] }), .sum({ \level_1_sums[11][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[211] [4:0] }), .sum({ \level_1_sums[11][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[11][105] [5:0] }),
     .b({ \level_1_sums[11][104] [5:0] }), .sum({ \level_2_sums[11][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[213] [4:0] }), .sum({ \level_1_sums[11][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[215] [4:0] }), .sum({ \level_1_sums[11][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[11][107] [5:0] }),
     .b({ \level_1_sums[11][106] [5:0] }), .sum({ \level_2_sums[11][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[11][53] [6:0] }), .b({ \level_2_sums[11][52] [6:0] }), .sum({ \level_3_sums[11][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[217] [4:0] }), .sum({ \level_1_sums[11][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[219] [4:0] }), .sum({ \level_1_sums[11][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[11][109] [5:0] }),
     .b({ \level_1_sums[11][108] [5:0] }), .sum({ \level_2_sums[11][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[221] [4:0] }), .sum({ \level_1_sums[11][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[223] [4:0] }), .sum({ \level_1_sums[11][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[11][111] [5:0] }),
     .b({ \level_1_sums[11][110] [5:0] }), .sum({ \level_2_sums[11][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[11][55] [6:0] }), .b({ \level_2_sums[11][54] [6:0] }), .sum({ \level_3_sums[11][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[11][27] [7:0] }),
     .b({ \level_3_sums[11][26] [7:0] }), .sum({ \level_4_sums[11][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[11][13] [8:0] }),
     .b({ \level_4_sums[11][12] [8:0] }), .sum({ \level_5_sums[11][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[225] [4:0] }), .sum({ \level_1_sums[11][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[227] [4:0] }), .sum({ \level_1_sums[11][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[11][113] [5:0] }),
     .b({ \level_1_sums[11][112] [5:0] }), .sum({ \level_2_sums[11][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[229] [4:0] }), .sum({ \level_1_sums[11][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[231] [4:0] }), .sum({ \level_1_sums[11][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[11][115] [5:0] }),
     .b({ \level_1_sums[11][114] [5:0] }), .sum({ \level_2_sums[11][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[11][57] [6:0] }), .b({ \level_2_sums[11][56] [6:0] }), .sum({ \level_3_sums[11][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[233] [4:0] }), .sum({ \level_1_sums[11][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[235] [4:0] }), .sum({ \level_1_sums[11][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[11][117] [5:0] }),
     .b({ \level_1_sums[11][116] [5:0] }), .sum({ \level_2_sums[11][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[237] [4:0] }), .sum({ \level_1_sums[11][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[239] [4:0] }), .sum({ \level_1_sums[11][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[11][119] [5:0] }),
     .b({ \level_1_sums[11][118] [5:0] }), .sum({ \level_2_sums[11][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[11][59] [6:0] }), .b({ \level_2_sums[11][58] [6:0] }), .sum({ \level_3_sums[11][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[11][29] [7:0] }),
     .b({ \level_3_sums[11][28] [7:0] }), .sum({ \level_4_sums[11][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[241] [4:0] }), .sum({ \level_1_sums[11][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[243] [4:0] }), .sum({ \level_1_sums[11][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[11][121] [5:0] }),
     .b({ \level_1_sums[11][120] [5:0] }), .sum({ \level_2_sums[11][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[245] [4:0] }), .sum({ \level_1_sums[11][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[247] [4:0] }), .sum({ \level_1_sums[11][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[11][123] [5:0] }),
     .b({ \level_1_sums[11][122] [5:0] }), .sum({ \level_2_sums[11][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[11][61] [6:0] }), .b({ \level_2_sums[11][60] [6:0] }), .sum({ \level_3_sums[11][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[249] [4:0] }), .sum({ \level_1_sums[11][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[251] [4:0] }), .sum({ \level_1_sums[11][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[11][125] [5:0] }),
     .b({ \level_1_sums[11][124] [5:0] }), .sum({ \level_2_sums[11][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[253] [4:0] }), .sum({ \level_1_sums[11][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[11].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[11].product_terms[255] [4:0] }), .sum({ \level_1_sums[11][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[11][127] [5:0] }),
     .b({ \level_1_sums[11][126] [5:0] }), .sum({ \level_2_sums[11][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[11][63] [6:0] }), .b({ \level_2_sums[11][62] [6:0] }), .sum({ \level_3_sums[11][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[11][31] [7:0] }),
     .b({ \level_3_sums[11][30] [7:0] }), .sum({ \level_4_sums[11][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[11][15] [8:0] }),
     .b({ \level_4_sums[11][14] [8:0] }), .sum({ \level_5_sums[11][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[11][7] [9:0] }),
     .b({ \level_5_sums[11][6] [9:0] }), .sum({ \level_6_sums[11][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[11][3] [9:0] }),
     .b({ \level_6_sums[11][2] [9:0] }), .sum({ \level_7_sums[11][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[11].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[11][0] [9:0] }),
     .b({ \level_7_sums[11][1] [9:0] }), .sum({ \level_8_sums[11] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[12].relu_inst (.in_data({ \final_sums[12] [9:0] }), .out_data({ \out_sig[12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[1] [4:0] }), .sum({ \level_1_sums[12][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[3] [4:0] }), .sum({ \level_1_sums[12][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[12][1] [5:0] }),
     .b({ \level_1_sums[12][0] [5:0] }), .sum({ \level_2_sums[12][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[5] [4:0] }), .sum({ \level_1_sums[12][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[7] [4:0] }), .sum({ \level_1_sums[12][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[12][3] [5:0] }),
     .b({ \level_1_sums[12][2] [5:0] }), .sum({ \level_2_sums[12][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[12][1] [6:0] }),
     .b({ \level_2_sums[12][0] [6:0] }), .sum({ \level_3_sums[12][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[9] [4:0] }), .sum({ \level_1_sums[12][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[11] [4:0] }), .sum({ \level_1_sums[12][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[12][5] [5:0] }),
     .b({ \level_1_sums[12][4] [5:0] }), .sum({ \level_2_sums[12][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[13] [4:0] }), .sum({ \level_1_sums[12][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[15] [4:0] }), .sum({ \level_1_sums[12][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[12][7] [5:0] }),
     .b({ \level_1_sums[12][6] [5:0] }), .sum({ \level_2_sums[12][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[12][3] [6:0] }),
     .b({ \level_2_sums[12][2] [6:0] }), .sum({ \level_3_sums[12][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[12][1] [7:0] }),
     .b({ \level_3_sums[12][0] [7:0] }), .sum({ \level_4_sums[12][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[17] [4:0] }), .sum({ \level_1_sums[12][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[19] [4:0] }), .sum({ \level_1_sums[12][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[12][9] [5:0] }),
     .b({ \level_1_sums[12][8] [5:0] }), .sum({ \level_2_sums[12][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[21] [4:0] }), .sum({ \level_1_sums[12][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[23] [4:0] }), .sum({ \level_1_sums[12][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[12][11] [5:0] }),
     .b({ \level_1_sums[12][10] [5:0] }), .sum({ \level_2_sums[12][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[12][5] [6:0] }),
     .b({ \level_2_sums[12][4] [6:0] }), .sum({ \level_3_sums[12][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[25] [4:0] }), .sum({ \level_1_sums[12][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[27] [4:0] }), .sum({ \level_1_sums[12][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[12][13] [5:0] }),
     .b({ \level_1_sums[12][12] [5:0] }), .sum({ \level_2_sums[12][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[29] [4:0] }), .sum({ \level_1_sums[12][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[31] [4:0] }), .sum({ \level_1_sums[12][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[12][15] [5:0] }),
     .b({ \level_1_sums[12][14] [5:0] }), .sum({ \level_2_sums[12][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[12][7] [6:0] }),
     .b({ \level_2_sums[12][6] [6:0] }), .sum({ \level_3_sums[12][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[12][3] [7:0] }),
     .b({ \level_3_sums[12][2] [7:0] }), .sum({ \level_4_sums[12][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[12][1] [8:0] }),
     .b({ \level_4_sums[12][0] [8:0] }), .sum({ \level_5_sums[12][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[33] [4:0] }), .sum({ \level_1_sums[12][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[35] [4:0] }), .sum({ \level_1_sums[12][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[12][17] [5:0] }),
     .b({ \level_1_sums[12][16] [5:0] }), .sum({ \level_2_sums[12][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[37] [4:0] }), .sum({ \level_1_sums[12][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[39] [4:0] }), .sum({ \level_1_sums[12][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[12][19] [5:0] }),
     .b({ \level_1_sums[12][18] [5:0] }), .sum({ \level_2_sums[12][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[12][9] [6:0] }),
     .b({ \level_2_sums[12][8] [6:0] }), .sum({ \level_3_sums[12][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[41] [4:0] }), .sum({ \level_1_sums[12][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[43] [4:0] }), .sum({ \level_1_sums[12][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[12][21] [5:0] }),
     .b({ \level_1_sums[12][20] [5:0] }), .sum({ \level_2_sums[12][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[45] [4:0] }), .sum({ \level_1_sums[12][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[47] [4:0] }), .sum({ \level_1_sums[12][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[12][23] [5:0] }),
     .b({ \level_1_sums[12][22] [5:0] }), .sum({ \level_2_sums[12][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[12][11] [6:0] }),
     .b({ \level_2_sums[12][10] [6:0] }), .sum({ \level_3_sums[12][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[12][5] [7:0] }),
     .b({ \level_3_sums[12][4] [7:0] }), .sum({ \level_4_sums[12][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[49] [4:0] }), .sum({ \level_1_sums[12][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[51] [4:0] }), .sum({ \level_1_sums[12][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[12][25] [5:0] }),
     .b({ \level_1_sums[12][24] [5:0] }), .sum({ \level_2_sums[12][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[53] [4:0] }), .sum({ \level_1_sums[12][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[55] [4:0] }), .sum({ \level_1_sums[12][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[12][27] [5:0] }),
     .b({ \level_1_sums[12][26] [5:0] }), .sum({ \level_2_sums[12][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[12][13] [6:0] }),
     .b({ \level_2_sums[12][12] [6:0] }), .sum({ \level_3_sums[12][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[57] [4:0] }), .sum({ \level_1_sums[12][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[59] [4:0] }), .sum({ \level_1_sums[12][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[12][29] [5:0] }),
     .b({ \level_1_sums[12][28] [5:0] }), .sum({ \level_2_sums[12][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[61] [4:0] }), .sum({ \level_1_sums[12][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[63] [4:0] }), .sum({ \level_1_sums[12][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[12][31] [5:0] }),
     .b({ \level_1_sums[12][30] [5:0] }), .sum({ \level_2_sums[12][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[12][15] [6:0] }),
     .b({ \level_2_sums[12][14] [6:0] }), .sum({ \level_3_sums[12][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[12][7] [7:0] }),
     .b({ \level_3_sums[12][6] [7:0] }), .sum({ \level_4_sums[12][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[12][3] [8:0] }),
     .b({ \level_4_sums[12][2] [8:0] }), .sum({ \level_5_sums[12][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[12][1] [9:0] }),
     .b({ \level_5_sums[12][0] [9:0] }), .sum({ \level_6_sums[12][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[65] [4:0] }), .sum({ \level_1_sums[12][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[67] [4:0] }), .sum({ \level_1_sums[12][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[12][33] [5:0] }),
     .b({ \level_1_sums[12][32] [5:0] }), .sum({ \level_2_sums[12][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[69] [4:0] }), .sum({ \level_1_sums[12][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[71] [4:0] }), .sum({ \level_1_sums[12][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[12][35] [5:0] }),
     .b({ \level_1_sums[12][34] [5:0] }), .sum({ \level_2_sums[12][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[12][17] [6:0] }),
     .b({ \level_2_sums[12][16] [6:0] }), .sum({ \level_3_sums[12][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[73] [4:0] }), .sum({ \level_1_sums[12][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[75] [4:0] }), .sum({ \level_1_sums[12][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[12][37] [5:0] }),
     .b({ \level_1_sums[12][36] [5:0] }), .sum({ \level_2_sums[12][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[77] [4:0] }), .sum({ \level_1_sums[12][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[79] [4:0] }), .sum({ \level_1_sums[12][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[12][39] [5:0] }),
     .b({ \level_1_sums[12][38] [5:0] }), .sum({ \level_2_sums[12][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[12][19] [6:0] }),
     .b({ \level_2_sums[12][18] [6:0] }), .sum({ \level_3_sums[12][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[12][9] [7:0] }),
     .b({ \level_3_sums[12][8] [7:0] }), .sum({ \level_4_sums[12][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[81] [4:0] }), .sum({ \level_1_sums[12][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[83] [4:0] }), .sum({ \level_1_sums[12][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[12][41] [5:0] }),
     .b({ \level_1_sums[12][40] [5:0] }), .sum({ \level_2_sums[12][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[85] [4:0] }), .sum({ \level_1_sums[12][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[87] [4:0] }), .sum({ \level_1_sums[12][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[12][43] [5:0] }),
     .b({ \level_1_sums[12][42] [5:0] }), .sum({ \level_2_sums[12][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[12][21] [6:0] }),
     .b({ \level_2_sums[12][20] [6:0] }), .sum({ \level_3_sums[12][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[89] [4:0] }), .sum({ \level_1_sums[12][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[91] [4:0] }), .sum({ \level_1_sums[12][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[12][45] [5:0] }),
     .b({ \level_1_sums[12][44] [5:0] }), .sum({ \level_2_sums[12][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[93] [4:0] }), .sum({ \level_1_sums[12][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[95] [4:0] }), .sum({ \level_1_sums[12][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[12][47] [5:0] }),
     .b({ \level_1_sums[12][46] [5:0] }), .sum({ \level_2_sums[12][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[12][23] [6:0] }),
     .b({ \level_2_sums[12][22] [6:0] }), .sum({ \level_3_sums[12][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[12][11] [7:0] }),
     .b({ \level_3_sums[12][10] [7:0] }), .sum({ \level_4_sums[12][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[12][5] [8:0] }),
     .b({ \level_4_sums[12][4] [8:0] }), .sum({ \level_5_sums[12][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[97] [4:0] }), .sum({ \level_1_sums[12][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[99] [4:0] }), .sum({ \level_1_sums[12][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[12][49] [5:0] }),
     .b({ \level_1_sums[12][48] [5:0] }), .sum({ \level_2_sums[12][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[101] [4:0] }), .sum({ \level_1_sums[12][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[103] [4:0] }), .sum({ \level_1_sums[12][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[12][51] [5:0] }),
     .b({ \level_1_sums[12][50] [5:0] }), .sum({ \level_2_sums[12][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[12][25] [6:0] }), .b({ \level_2_sums[12][24] [6:0] }), .sum({ \level_3_sums[12][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[105] [4:0] }), .sum({ \level_1_sums[12][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[107] [4:0] }), .sum({ \level_1_sums[12][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[12][53] [5:0] }),
     .b({ \level_1_sums[12][52] [5:0] }), .sum({ \level_2_sums[12][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[109] [4:0] }), .sum({ \level_1_sums[12][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[111] [4:0] }), .sum({ \level_1_sums[12][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[12][55] [5:0] }),
     .b({ \level_1_sums[12][54] [5:0] }), .sum({ \level_2_sums[12][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[12][27] [6:0] }), .b({ \level_2_sums[12][26] [6:0] }), .sum({ \level_3_sums[12][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[12][13] [7:0] }),
     .b({ \level_3_sums[12][12] [7:0] }), .sum({ \level_4_sums[12][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[113] [4:0] }), .sum({ \level_1_sums[12][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[115] [4:0] }), .sum({ \level_1_sums[12][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[12][57] [5:0] }),
     .b({ \level_1_sums[12][56] [5:0] }), .sum({ \level_2_sums[12][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[117] [4:0] }), .sum({ \level_1_sums[12][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[119] [4:0] }), .sum({ \level_1_sums[12][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[12][59] [5:0] }),
     .b({ \level_1_sums[12][58] [5:0] }), .sum({ \level_2_sums[12][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[12][29] [6:0] }), .b({ \level_2_sums[12][28] [6:0] }), .sum({ \level_3_sums[12][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[121] [4:0] }), .sum({ \level_1_sums[12][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[123] [4:0] }), .sum({ \level_1_sums[12][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[12][61] [5:0] }),
     .b({ \level_1_sums[12][60] [5:0] }), .sum({ \level_2_sums[12][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[125] [4:0] }), .sum({ \level_1_sums[12][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[127] [4:0] }), .sum({ \level_1_sums[12][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[12][63] [5:0] }),
     .b({ \level_1_sums[12][62] [5:0] }), .sum({ \level_2_sums[12][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[12][31] [6:0] }), .b({ \level_2_sums[12][30] [6:0] }), .sum({ \level_3_sums[12][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[12][15] [7:0] }),
     .b({ \level_3_sums[12][14] [7:0] }), .sum({ \level_4_sums[12][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[12][7] [8:0] }),
     .b({ \level_4_sums[12][6] [8:0] }), .sum({ \level_5_sums[12][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[12][3] [9:0] }),
     .b({ \level_5_sums[12][2] [9:0] }), .sum({ \level_6_sums[12][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[12][1] [9:0] }),
     .b({ \level_6_sums[12][0] [9:0] }), .sum({ \level_7_sums[12][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[129] [4:0] }), .sum({ \level_1_sums[12][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[131] [4:0] }), .sum({ \level_1_sums[12][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[12][65] [5:0] }),
     .b({ \level_1_sums[12][64] [5:0] }), .sum({ \level_2_sums[12][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[133] [4:0] }), .sum({ \level_1_sums[12][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[135] [4:0] }), .sum({ \level_1_sums[12][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[12][67] [5:0] }),
     .b({ \level_1_sums[12][66] [5:0] }), .sum({ \level_2_sums[12][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[12][33] [6:0] }), .b({ \level_2_sums[12][32] [6:0] }), .sum({ \level_3_sums[12][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[137] [4:0] }), .sum({ \level_1_sums[12][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[139] [4:0] }), .sum({ \level_1_sums[12][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[12][69] [5:0] }),
     .b({ \level_1_sums[12][68] [5:0] }), .sum({ \level_2_sums[12][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[141] [4:0] }), .sum({ \level_1_sums[12][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[143] [4:0] }), .sum({ \level_1_sums[12][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[12][71] [5:0] }),
     .b({ \level_1_sums[12][70] [5:0] }), .sum({ \level_2_sums[12][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[12][35] [6:0] }), .b({ \level_2_sums[12][34] [6:0] }), .sum({ \level_3_sums[12][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[12][17] [7:0] }),
     .b({ \level_3_sums[12][16] [7:0] }), .sum({ \level_4_sums[12][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[145] [4:0] }), .sum({ \level_1_sums[12][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[147] [4:0] }), .sum({ \level_1_sums[12][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[12][73] [5:0] }),
     .b({ \level_1_sums[12][72] [5:0] }), .sum({ \level_2_sums[12][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[149] [4:0] }), .sum({ \level_1_sums[12][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[151] [4:0] }), .sum({ \level_1_sums[12][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[12][75] [5:0] }),
     .b({ \level_1_sums[12][74] [5:0] }), .sum({ \level_2_sums[12][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[12][37] [6:0] }), .b({ \level_2_sums[12][36] [6:0] }), .sum({ \level_3_sums[12][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[153] [4:0] }), .sum({ \level_1_sums[12][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[155] [4:0] }), .sum({ \level_1_sums[12][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[12][77] [5:0] }),
     .b({ \level_1_sums[12][76] [5:0] }), .sum({ \level_2_sums[12][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[157] [4:0] }), .sum({ \level_1_sums[12][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[159] [4:0] }), .sum({ \level_1_sums[12][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[12][79] [5:0] }),
     .b({ \level_1_sums[12][78] [5:0] }), .sum({ \level_2_sums[12][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[12][39] [6:0] }), .b({ \level_2_sums[12][38] [6:0] }), .sum({ \level_3_sums[12][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[12][19] [7:0] }),
     .b({ \level_3_sums[12][18] [7:0] }), .sum({ \level_4_sums[12][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[12][9] [8:0] }),
     .b({ \level_4_sums[12][8] [8:0] }), .sum({ \level_5_sums[12][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[161] [4:0] }), .sum({ \level_1_sums[12][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[163] [4:0] }), .sum({ \level_1_sums[12][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[12][81] [5:0] }),
     .b({ \level_1_sums[12][80] [5:0] }), .sum({ \level_2_sums[12][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[165] [4:0] }), .sum({ \level_1_sums[12][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[167] [4:0] }), .sum({ \level_1_sums[12][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[12][83] [5:0] }),
     .b({ \level_1_sums[12][82] [5:0] }), .sum({ \level_2_sums[12][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[12][41] [6:0] }), .b({ \level_2_sums[12][40] [6:0] }), .sum({ \level_3_sums[12][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[169] [4:0] }), .sum({ \level_1_sums[12][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[171] [4:0] }), .sum({ \level_1_sums[12][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[12][85] [5:0] }),
     .b({ \level_1_sums[12][84] [5:0] }), .sum({ \level_2_sums[12][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[173] [4:0] }), .sum({ \level_1_sums[12][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[175] [4:0] }), .sum({ \level_1_sums[12][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[12][87] [5:0] }),
     .b({ \level_1_sums[12][86] [5:0] }), .sum({ \level_2_sums[12][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[12][43] [6:0] }), .b({ \level_2_sums[12][42] [6:0] }), .sum({ \level_3_sums[12][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[12][21] [7:0] }),
     .b({ \level_3_sums[12][20] [7:0] }), .sum({ \level_4_sums[12][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[177] [4:0] }), .sum({ \level_1_sums[12][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[179] [4:0] }), .sum({ \level_1_sums[12][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[12][89] [5:0] }),
     .b({ \level_1_sums[12][88] [5:0] }), .sum({ \level_2_sums[12][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[181] [4:0] }), .sum({ \level_1_sums[12][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[183] [4:0] }), .sum({ \level_1_sums[12][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[12][91] [5:0] }),
     .b({ \level_1_sums[12][90] [5:0] }), .sum({ \level_2_sums[12][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[12][45] [6:0] }), .b({ \level_2_sums[12][44] [6:0] }), .sum({ \level_3_sums[12][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[185] [4:0] }), .sum({ \level_1_sums[12][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[187] [4:0] }), .sum({ \level_1_sums[12][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[12][93] [5:0] }),
     .b({ \level_1_sums[12][92] [5:0] }), .sum({ \level_2_sums[12][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[189] [4:0] }), .sum({ \level_1_sums[12][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[191] [4:0] }), .sum({ \level_1_sums[12][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[12][95] [5:0] }),
     .b({ \level_1_sums[12][94] [5:0] }), .sum({ \level_2_sums[12][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[12][47] [6:0] }), .b({ \level_2_sums[12][46] [6:0] }), .sum({ \level_3_sums[12][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[12][23] [7:0] }),
     .b({ \level_3_sums[12][22] [7:0] }), .sum({ \level_4_sums[12][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[12][11] [8:0] }),
     .b({ \level_4_sums[12][10] [8:0] }), .sum({ \level_5_sums[12][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[12][5] [9:0] }),
     .b({ \level_5_sums[12][4] [9:0] }), .sum({ \level_6_sums[12][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[193] [4:0] }), .sum({ \level_1_sums[12][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[195] [4:0] }), .sum({ \level_1_sums[12][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[12][97] [5:0] }),
     .b({ \level_1_sums[12][96] [5:0] }), .sum({ \level_2_sums[12][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[197] [4:0] }), .sum({ \level_1_sums[12][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[199] [4:0] }), .sum({ \level_1_sums[12][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[12][99] [5:0] }),
     .b({ \level_1_sums[12][98] [5:0] }), .sum({ \level_2_sums[12][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[12][49] [6:0] }), .b({ \level_2_sums[12][48] [6:0] }), .sum({ \level_3_sums[12][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[201] [4:0] }), .sum({ \level_1_sums[12][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[203] [4:0] }), .sum({ \level_1_sums[12][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[12][101] [5:0] }),
     .b({ \level_1_sums[12][100] [5:0] }), .sum({ \level_2_sums[12][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[205] [4:0] }), .sum({ \level_1_sums[12][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[207] [4:0] }), .sum({ \level_1_sums[12][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[12][103] [5:0] }),
     .b({ \level_1_sums[12][102] [5:0] }), .sum({ \level_2_sums[12][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[12][51] [6:0] }), .b({ \level_2_sums[12][50] [6:0] }), .sum({ \level_3_sums[12][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[12][25] [7:0] }),
     .b({ \level_3_sums[12][24] [7:0] }), .sum({ \level_4_sums[12][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[209] [4:0] }), .sum({ \level_1_sums[12][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[211] [4:0] }), .sum({ \level_1_sums[12][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[12][105] [5:0] }),
     .b({ \level_1_sums[12][104] [5:0] }), .sum({ \level_2_sums[12][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[213] [4:0] }), .sum({ \level_1_sums[12][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[215] [4:0] }), .sum({ \level_1_sums[12][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[12][107] [5:0] }),
     .b({ \level_1_sums[12][106] [5:0] }), .sum({ \level_2_sums[12][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[12][53] [6:0] }), .b({ \level_2_sums[12][52] [6:0] }), .sum({ \level_3_sums[12][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[217] [4:0] }), .sum({ \level_1_sums[12][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[219] [4:0] }), .sum({ \level_1_sums[12][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[12][109] [5:0] }),
     .b({ \level_1_sums[12][108] [5:0] }), .sum({ \level_2_sums[12][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[221] [4:0] }), .sum({ \level_1_sums[12][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[223] [4:0] }), .sum({ \level_1_sums[12][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[12][111] [5:0] }),
     .b({ \level_1_sums[12][110] [5:0] }), .sum({ \level_2_sums[12][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[12][55] [6:0] }), .b({ \level_2_sums[12][54] [6:0] }), .sum({ \level_3_sums[12][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[12][27] [7:0] }),
     .b({ \level_3_sums[12][26] [7:0] }), .sum({ \level_4_sums[12][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[12][13] [8:0] }),
     .b({ \level_4_sums[12][12] [8:0] }), .sum({ \level_5_sums[12][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[225] [4:0] }), .sum({ \level_1_sums[12][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[227] [4:0] }), .sum({ \level_1_sums[12][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[12][113] [5:0] }),
     .b({ \level_1_sums[12][112] [5:0] }), .sum({ \level_2_sums[12][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[229] [4:0] }), .sum({ \level_1_sums[12][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[231] [4:0] }), .sum({ \level_1_sums[12][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[12][115] [5:0] }),
     .b({ \level_1_sums[12][114] [5:0] }), .sum({ \level_2_sums[12][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[12][57] [6:0] }), .b({ \level_2_sums[12][56] [6:0] }), .sum({ \level_3_sums[12][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[233] [4:0] }), .sum({ \level_1_sums[12][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[235] [4:0] }), .sum({ \level_1_sums[12][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[12][117] [5:0] }),
     .b({ \level_1_sums[12][116] [5:0] }), .sum({ \level_2_sums[12][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[237] [4:0] }), .sum({ \level_1_sums[12][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[239] [4:0] }), .sum({ \level_1_sums[12][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[12][119] [5:0] }),
     .b({ \level_1_sums[12][118] [5:0] }), .sum({ \level_2_sums[12][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[12][59] [6:0] }), .b({ \level_2_sums[12][58] [6:0] }), .sum({ \level_3_sums[12][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[12][29] [7:0] }),
     .b({ \level_3_sums[12][28] [7:0] }), .sum({ \level_4_sums[12][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[241] [4:0] }), .sum({ \level_1_sums[12][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[243] [4:0] }), .sum({ \level_1_sums[12][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[12][121] [5:0] }),
     .b({ \level_1_sums[12][120] [5:0] }), .sum({ \level_2_sums[12][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[245] [4:0] }), .sum({ \level_1_sums[12][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[247] [4:0] }), .sum({ \level_1_sums[12][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[12][123] [5:0] }),
     .b({ \level_1_sums[12][122] [5:0] }), .sum({ \level_2_sums[12][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[12][61] [6:0] }), .b({ \level_2_sums[12][60] [6:0] }), .sum({ \level_3_sums[12][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[249] [4:0] }), .sum({ \level_1_sums[12][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[251] [4:0] }), .sum({ \level_1_sums[12][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[12][125] [5:0] }),
     .b({ \level_1_sums[12][124] [5:0] }), .sum({ \level_2_sums[12][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[253] [4:0] }), .sum({ \level_1_sums[12][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[12].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[12].product_terms[255] [4:0] }), .sum({ \level_1_sums[12][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[12][127] [5:0] }),
     .b({ \level_1_sums[12][126] [5:0] }), .sum({ \level_2_sums[12][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[12][63] [6:0] }), .b({ \level_2_sums[12][62] [6:0] }), .sum({ \level_3_sums[12][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[12][31] [7:0] }),
     .b({ \level_3_sums[12][30] [7:0] }), .sum({ \level_4_sums[12][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[12][15] [8:0] }),
     .b({ \level_4_sums[12][14] [8:0] }), .sum({ \level_5_sums[12][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[12][7] [9:0] }),
     .b({ \level_5_sums[12][6] [9:0] }), .sum({ \level_6_sums[12][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[12][3] [9:0] }),
     .b({ \level_6_sums[12][2] [9:0] }), .sum({ \level_7_sums[12][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[12].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[12][0] [9:0] }),
     .b({ \level_7_sums[12][1] [9:0] }), .sum({ \level_8_sums[12] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[13].relu_inst (.in_data({ \final_sums[13] [9:0] }), .out_data({ \out_sig[13] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[1] [4:0] }), .sum({ \level_1_sums[13][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[3] [4:0] }), .sum({ \level_1_sums[13][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[13][1] [5:0] }),
     .b({ \level_1_sums[13][0] [5:0] }), .sum({ \level_2_sums[13][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[5] [4:0] }), .sum({ \level_1_sums[13][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[7] [4:0] }), .sum({ \level_1_sums[13][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[13][3] [5:0] }),
     .b({ \level_1_sums[13][2] [5:0] }), .sum({ \level_2_sums[13][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[13][1] [6:0] }),
     .b({ \level_2_sums[13][0] [6:0] }), .sum({ \level_3_sums[13][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[9] [4:0] }), .sum({ \level_1_sums[13][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[11] [4:0] }), .sum({ \level_1_sums[13][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[13][5] [5:0] }),
     .b({ \level_1_sums[13][4] [5:0] }), .sum({ \level_2_sums[13][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[13] [4:0] }), .sum({ \level_1_sums[13][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[15] [4:0] }), .sum({ \level_1_sums[13][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[13][7] [5:0] }),
     .b({ \level_1_sums[13][6] [5:0] }), .sum({ \level_2_sums[13][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[13][3] [6:0] }),
     .b({ \level_2_sums[13][2] [6:0] }), .sum({ \level_3_sums[13][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[13][1] [7:0] }),
     .b({ \level_3_sums[13][0] [7:0] }), .sum({ \level_4_sums[13][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[17] [4:0] }), .sum({ \level_1_sums[13][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[19] [4:0] }), .sum({ \level_1_sums[13][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[13][9] [5:0] }),
     .b({ \level_1_sums[13][8] [5:0] }), .sum({ \level_2_sums[13][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[21] [4:0] }), .sum({ \level_1_sums[13][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[23] [4:0] }), .sum({ \level_1_sums[13][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[13][11] [5:0] }),
     .b({ \level_1_sums[13][10] [5:0] }), .sum({ \level_2_sums[13][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[13][5] [6:0] }),
     .b({ \level_2_sums[13][4] [6:0] }), .sum({ \level_3_sums[13][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[25] [4:0] }), .sum({ \level_1_sums[13][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[27] [4:0] }), .sum({ \level_1_sums[13][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[13][13] [5:0] }),
     .b({ \level_1_sums[13][12] [5:0] }), .sum({ \level_2_sums[13][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[29] [4:0] }), .sum({ \level_1_sums[13][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[31] [4:0] }), .sum({ \level_1_sums[13][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[13][15] [5:0] }),
     .b({ \level_1_sums[13][14] [5:0] }), .sum({ \level_2_sums[13][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[13][7] [6:0] }),
     .b({ \level_2_sums[13][6] [6:0] }), .sum({ \level_3_sums[13][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[13][3] [7:0] }),
     .b({ \level_3_sums[13][2] [7:0] }), .sum({ \level_4_sums[13][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[13][1] [8:0] }),
     .b({ \level_4_sums[13][0] [8:0] }), .sum({ \level_5_sums[13][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[33] [4:0] }), .sum({ \level_1_sums[13][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[35] [4:0] }), .sum({ \level_1_sums[13][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[13][17] [5:0] }),
     .b({ \level_1_sums[13][16] [5:0] }), .sum({ \level_2_sums[13][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[37] [4:0] }), .sum({ \level_1_sums[13][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[39] [4:0] }), .sum({ \level_1_sums[13][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[13][19] [5:0] }),
     .b({ \level_1_sums[13][18] [5:0] }), .sum({ \level_2_sums[13][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[13][9] [6:0] }),
     .b({ \level_2_sums[13][8] [6:0] }), .sum({ \level_3_sums[13][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[41] [4:0] }), .sum({ \level_1_sums[13][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[43] [4:0] }), .sum({ \level_1_sums[13][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[13][21] [5:0] }),
     .b({ \level_1_sums[13][20] [5:0] }), .sum({ \level_2_sums[13][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[45] [4:0] }), .sum({ \level_1_sums[13][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[47] [4:0] }), .sum({ \level_1_sums[13][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[13][23] [5:0] }),
     .b({ \level_1_sums[13][22] [5:0] }), .sum({ \level_2_sums[13][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[13][11] [6:0] }),
     .b({ \level_2_sums[13][10] [6:0] }), .sum({ \level_3_sums[13][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[13][5] [7:0] }),
     .b({ \level_3_sums[13][4] [7:0] }), .sum({ \level_4_sums[13][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[49] [4:0] }), .sum({ \level_1_sums[13][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[51] [4:0] }), .sum({ \level_1_sums[13][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[13][25] [5:0] }),
     .b({ \level_1_sums[13][24] [5:0] }), .sum({ \level_2_sums[13][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[53] [4:0] }), .sum({ \level_1_sums[13][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[55] [4:0] }), .sum({ \level_1_sums[13][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[13][27] [5:0] }),
     .b({ \level_1_sums[13][26] [5:0] }), .sum({ \level_2_sums[13][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[13][13] [6:0] }),
     .b({ \level_2_sums[13][12] [6:0] }), .sum({ \level_3_sums[13][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[57] [4:0] }), .sum({ \level_1_sums[13][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[59] [4:0] }), .sum({ \level_1_sums[13][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[13][29] [5:0] }),
     .b({ \level_1_sums[13][28] [5:0] }), .sum({ \level_2_sums[13][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[61] [4:0] }), .sum({ \level_1_sums[13][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[63] [4:0] }), .sum({ \level_1_sums[13][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[13][31] [5:0] }),
     .b({ \level_1_sums[13][30] [5:0] }), .sum({ \level_2_sums[13][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[13][15] [6:0] }),
     .b({ \level_2_sums[13][14] [6:0] }), .sum({ \level_3_sums[13][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[13][7] [7:0] }),
     .b({ \level_3_sums[13][6] [7:0] }), .sum({ \level_4_sums[13][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[13][3] [8:0] }),
     .b({ \level_4_sums[13][2] [8:0] }), .sum({ \level_5_sums[13][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[13][1] [9:0] }),
     .b({ \level_5_sums[13][0] [9:0] }), .sum({ \level_6_sums[13][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[65] [4:0] }), .sum({ \level_1_sums[13][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[67] [4:0] }), .sum({ \level_1_sums[13][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[13][33] [5:0] }),
     .b({ \level_1_sums[13][32] [5:0] }), .sum({ \level_2_sums[13][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[69] [4:0] }), .sum({ \level_1_sums[13][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[71] [4:0] }), .sum({ \level_1_sums[13][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[13][35] [5:0] }),
     .b({ \level_1_sums[13][34] [5:0] }), .sum({ \level_2_sums[13][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[13][17] [6:0] }),
     .b({ \level_2_sums[13][16] [6:0] }), .sum({ \level_3_sums[13][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[73] [4:0] }), .sum({ \level_1_sums[13][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[75] [4:0] }), .sum({ \level_1_sums[13][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[13][37] [5:0] }),
     .b({ \level_1_sums[13][36] [5:0] }), .sum({ \level_2_sums[13][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[77] [4:0] }), .sum({ \level_1_sums[13][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[79] [4:0] }), .sum({ \level_1_sums[13][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[13][39] [5:0] }),
     .b({ \level_1_sums[13][38] [5:0] }), .sum({ \level_2_sums[13][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[13][19] [6:0] }),
     .b({ \level_2_sums[13][18] [6:0] }), .sum({ \level_3_sums[13][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[13][9] [7:0] }),
     .b({ \level_3_sums[13][8] [7:0] }), .sum({ \level_4_sums[13][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[81] [4:0] }), .sum({ \level_1_sums[13][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[83] [4:0] }), .sum({ \level_1_sums[13][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[13][41] [5:0] }),
     .b({ \level_1_sums[13][40] [5:0] }), .sum({ \level_2_sums[13][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[85] [4:0] }), .sum({ \level_1_sums[13][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[87] [4:0] }), .sum({ \level_1_sums[13][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[13][43] [5:0] }),
     .b({ \level_1_sums[13][42] [5:0] }), .sum({ \level_2_sums[13][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[13][21] [6:0] }),
     .b({ \level_2_sums[13][20] [6:0] }), .sum({ \level_3_sums[13][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[89] [4:0] }), .sum({ \level_1_sums[13][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[91] [4:0] }), .sum({ \level_1_sums[13][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[13][45] [5:0] }),
     .b({ \level_1_sums[13][44] [5:0] }), .sum({ \level_2_sums[13][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[93] [4:0] }), .sum({ \level_1_sums[13][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[95] [4:0] }), .sum({ \level_1_sums[13][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[13][47] [5:0] }),
     .b({ \level_1_sums[13][46] [5:0] }), .sum({ \level_2_sums[13][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[13][23] [6:0] }),
     .b({ \level_2_sums[13][22] [6:0] }), .sum({ \level_3_sums[13][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[13][11] [7:0] }),
     .b({ \level_3_sums[13][10] [7:0] }), .sum({ \level_4_sums[13][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[13][5] [8:0] }),
     .b({ \level_4_sums[13][4] [8:0] }), .sum({ \level_5_sums[13][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[97] [4:0] }), .sum({ \level_1_sums[13][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[99] [4:0] }), .sum({ \level_1_sums[13][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[13][49] [5:0] }),
     .b({ \level_1_sums[13][48] [5:0] }), .sum({ \level_2_sums[13][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[101] [4:0] }), .sum({ \level_1_sums[13][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[103] [4:0] }), .sum({ \level_1_sums[13][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[13][51] [5:0] }),
     .b({ \level_1_sums[13][50] [5:0] }), .sum({ \level_2_sums[13][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[13][25] [6:0] }), .b({ \level_2_sums[13][24] [6:0] }), .sum({ \level_3_sums[13][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[105] [4:0] }), .sum({ \level_1_sums[13][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[107] [4:0] }), .sum({ \level_1_sums[13][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[13][53] [5:0] }),
     .b({ \level_1_sums[13][52] [5:0] }), .sum({ \level_2_sums[13][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[109] [4:0] }), .sum({ \level_1_sums[13][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[111] [4:0] }), .sum({ \level_1_sums[13][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[13][55] [5:0] }),
     .b({ \level_1_sums[13][54] [5:0] }), .sum({ \level_2_sums[13][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[13][27] [6:0] }), .b({ \level_2_sums[13][26] [6:0] }), .sum({ \level_3_sums[13][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[13][13] [7:0] }),
     .b({ \level_3_sums[13][12] [7:0] }), .sum({ \level_4_sums[13][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[113] [4:0] }), .sum({ \level_1_sums[13][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[115] [4:0] }), .sum({ \level_1_sums[13][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[13][57] [5:0] }),
     .b({ \level_1_sums[13][56] [5:0] }), .sum({ \level_2_sums[13][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[117] [4:0] }), .sum({ \level_1_sums[13][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[119] [4:0] }), .sum({ \level_1_sums[13][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[13][59] [5:0] }),
     .b({ \level_1_sums[13][58] [5:0] }), .sum({ \level_2_sums[13][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[13][29] [6:0] }), .b({ \level_2_sums[13][28] [6:0] }), .sum({ \level_3_sums[13][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[121] [4:0] }), .sum({ \level_1_sums[13][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[123] [4:0] }), .sum({ \level_1_sums[13][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[13][61] [5:0] }),
     .b({ \level_1_sums[13][60] [5:0] }), .sum({ \level_2_sums[13][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[125] [4:0] }), .sum({ \level_1_sums[13][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[127] [4:0] }), .sum({ \level_1_sums[13][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[13][63] [5:0] }),
     .b({ \level_1_sums[13][62] [5:0] }), .sum({ \level_2_sums[13][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[13][31] [6:0] }), .b({ \level_2_sums[13][30] [6:0] }), .sum({ \level_3_sums[13][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[13][15] [7:0] }),
     .b({ \level_3_sums[13][14] [7:0] }), .sum({ \level_4_sums[13][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[13][7] [8:0] }),
     .b({ \level_4_sums[13][6] [8:0] }), .sum({ \level_5_sums[13][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[13][3] [9:0] }),
     .b({ \level_5_sums[13][2] [9:0] }), .sum({ \level_6_sums[13][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[13][1] [9:0] }),
     .b({ \level_6_sums[13][0] [9:0] }), .sum({ \level_7_sums[13][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[129] [4:0] }), .sum({ \level_1_sums[13][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[131] [4:0] }), .sum({ \level_1_sums[13][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[13][65] [5:0] }),
     .b({ \level_1_sums[13][64] [5:0] }), .sum({ \level_2_sums[13][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[133] [4:0] }), .sum({ \level_1_sums[13][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[135] [4:0] }), .sum({ \level_1_sums[13][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[13][67] [5:0] }),
     .b({ \level_1_sums[13][66] [5:0] }), .sum({ \level_2_sums[13][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[13][33] [6:0] }), .b({ \level_2_sums[13][32] [6:0] }), .sum({ \level_3_sums[13][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[137] [4:0] }), .sum({ \level_1_sums[13][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[139] [4:0] }), .sum({ \level_1_sums[13][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[13][69] [5:0] }),
     .b({ \level_1_sums[13][68] [5:0] }), .sum({ \level_2_sums[13][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[141] [4:0] }), .sum({ \level_1_sums[13][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[143] [4:0] }), .sum({ \level_1_sums[13][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[13][71] [5:0] }),
     .b({ \level_1_sums[13][70] [5:0] }), .sum({ \level_2_sums[13][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[13][35] [6:0] }), .b({ \level_2_sums[13][34] [6:0] }), .sum({ \level_3_sums[13][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[13][17] [7:0] }),
     .b({ \level_3_sums[13][16] [7:0] }), .sum({ \level_4_sums[13][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[145] [4:0] }), .sum({ \level_1_sums[13][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[147] [4:0] }), .sum({ \level_1_sums[13][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[13][73] [5:0] }),
     .b({ \level_1_sums[13][72] [5:0] }), .sum({ \level_2_sums[13][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[149] [4:0] }), .sum({ \level_1_sums[13][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[151] [4:0] }), .sum({ \level_1_sums[13][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[13][75] [5:0] }),
     .b({ \level_1_sums[13][74] [5:0] }), .sum({ \level_2_sums[13][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[13][37] [6:0] }), .b({ \level_2_sums[13][36] [6:0] }), .sum({ \level_3_sums[13][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[153] [4:0] }), .sum({ \level_1_sums[13][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[155] [4:0] }), .sum({ \level_1_sums[13][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[13][77] [5:0] }),
     .b({ \level_1_sums[13][76] [5:0] }), .sum({ \level_2_sums[13][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[157] [4:0] }), .sum({ \level_1_sums[13][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[159] [4:0] }), .sum({ \level_1_sums[13][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[13][79] [5:0] }),
     .b({ \level_1_sums[13][78] [5:0] }), .sum({ \level_2_sums[13][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[13][39] [6:0] }), .b({ \level_2_sums[13][38] [6:0] }), .sum({ \level_3_sums[13][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[13][19] [7:0] }),
     .b({ \level_3_sums[13][18] [7:0] }), .sum({ \level_4_sums[13][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[13][9] [8:0] }),
     .b({ \level_4_sums[13][8] [8:0] }), .sum({ \level_5_sums[13][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[161] [4:0] }), .sum({ \level_1_sums[13][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[163] [4:0] }), .sum({ \level_1_sums[13][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[13][81] [5:0] }),
     .b({ \level_1_sums[13][80] [5:0] }), .sum({ \level_2_sums[13][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[165] [4:0] }), .sum({ \level_1_sums[13][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[167] [4:0] }), .sum({ \level_1_sums[13][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[13][83] [5:0] }),
     .b({ \level_1_sums[13][82] [5:0] }), .sum({ \level_2_sums[13][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[13][41] [6:0] }), .b({ \level_2_sums[13][40] [6:0] }), .sum({ \level_3_sums[13][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[169] [4:0] }), .sum({ \level_1_sums[13][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[171] [4:0] }), .sum({ \level_1_sums[13][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[13][85] [5:0] }),
     .b({ \level_1_sums[13][84] [5:0] }), .sum({ \level_2_sums[13][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[173] [4:0] }), .sum({ \level_1_sums[13][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[175] [4:0] }), .sum({ \level_1_sums[13][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[13][87] [5:0] }),
     .b({ \level_1_sums[13][86] [5:0] }), .sum({ \level_2_sums[13][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[13][43] [6:0] }), .b({ \level_2_sums[13][42] [6:0] }), .sum({ \level_3_sums[13][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[13][21] [7:0] }),
     .b({ \level_3_sums[13][20] [7:0] }), .sum({ \level_4_sums[13][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[177] [4:0] }), .sum({ \level_1_sums[13][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[179] [4:0] }), .sum({ \level_1_sums[13][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[13][89] [5:0] }),
     .b({ \level_1_sums[13][88] [5:0] }), .sum({ \level_2_sums[13][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[181] [4:0] }), .sum({ \level_1_sums[13][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[183] [4:0] }), .sum({ \level_1_sums[13][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[13][91] [5:0] }),
     .b({ \level_1_sums[13][90] [5:0] }), .sum({ \level_2_sums[13][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[13][45] [6:0] }), .b({ \level_2_sums[13][44] [6:0] }), .sum({ \level_3_sums[13][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[185] [4:0] }), .sum({ \level_1_sums[13][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[187] [4:0] }), .sum({ \level_1_sums[13][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[13][93] [5:0] }),
     .b({ \level_1_sums[13][92] [5:0] }), .sum({ \level_2_sums[13][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[189] [4:0] }), .sum({ \level_1_sums[13][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[191] [4:0] }), .sum({ \level_1_sums[13][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[13][95] [5:0] }),
     .b({ \level_1_sums[13][94] [5:0] }), .sum({ \level_2_sums[13][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[13][47] [6:0] }), .b({ \level_2_sums[13][46] [6:0] }), .sum({ \level_3_sums[13][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[13][23] [7:0] }),
     .b({ \level_3_sums[13][22] [7:0] }), .sum({ \level_4_sums[13][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[13][11] [8:0] }),
     .b({ \level_4_sums[13][10] [8:0] }), .sum({ \level_5_sums[13][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[13][5] [9:0] }),
     .b({ \level_5_sums[13][4] [9:0] }), .sum({ \level_6_sums[13][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[193] [4:0] }), .sum({ \level_1_sums[13][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[195] [4:0] }), .sum({ \level_1_sums[13][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[13][97] [5:0] }),
     .b({ \level_1_sums[13][96] [5:0] }), .sum({ \level_2_sums[13][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[197] [4:0] }), .sum({ \level_1_sums[13][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[199] [4:0] }), .sum({ \level_1_sums[13][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[13][99] [5:0] }),
     .b({ \level_1_sums[13][98] [5:0] }), .sum({ \level_2_sums[13][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[13][49] [6:0] }), .b({ \level_2_sums[13][48] [6:0] }), .sum({ \level_3_sums[13][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[201] [4:0] }), .sum({ \level_1_sums[13][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[203] [4:0] }), .sum({ \level_1_sums[13][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[13][101] [5:0] }),
     .b({ \level_1_sums[13][100] [5:0] }), .sum({ \level_2_sums[13][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[205] [4:0] }), .sum({ \level_1_sums[13][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[207] [4:0] }), .sum({ \level_1_sums[13][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[13][103] [5:0] }),
     .b({ \level_1_sums[13][102] [5:0] }), .sum({ \level_2_sums[13][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[13][51] [6:0] }), .b({ \level_2_sums[13][50] [6:0] }), .sum({ \level_3_sums[13][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[13][25] [7:0] }),
     .b({ \level_3_sums[13][24] [7:0] }), .sum({ \level_4_sums[13][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[209] [4:0] }), .sum({ \level_1_sums[13][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[211] [4:0] }), .sum({ \level_1_sums[13][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[13][105] [5:0] }),
     .b({ \level_1_sums[13][104] [5:0] }), .sum({ \level_2_sums[13][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[213] [4:0] }), .sum({ \level_1_sums[13][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[215] [4:0] }), .sum({ \level_1_sums[13][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[13][107] [5:0] }),
     .b({ \level_1_sums[13][106] [5:0] }), .sum({ \level_2_sums[13][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[13][53] [6:0] }), .b({ \level_2_sums[13][52] [6:0] }), .sum({ \level_3_sums[13][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[217] [4:0] }), .sum({ \level_1_sums[13][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[219] [4:0] }), .sum({ \level_1_sums[13][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[13][109] [5:0] }),
     .b({ \level_1_sums[13][108] [5:0] }), .sum({ \level_2_sums[13][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[221] [4:0] }), .sum({ \level_1_sums[13][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[223] [4:0] }), .sum({ \level_1_sums[13][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[13][111] [5:0] }),
     .b({ \level_1_sums[13][110] [5:0] }), .sum({ \level_2_sums[13][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[13][55] [6:0] }), .b({ \level_2_sums[13][54] [6:0] }), .sum({ \level_3_sums[13][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[13][27] [7:0] }),
     .b({ \level_3_sums[13][26] [7:0] }), .sum({ \level_4_sums[13][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[13][13] [8:0] }),
     .b({ \level_4_sums[13][12] [8:0] }), .sum({ \level_5_sums[13][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[225] [4:0] }), .sum({ \level_1_sums[13][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[227] [4:0] }), .sum({ \level_1_sums[13][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[13][113] [5:0] }),
     .b({ \level_1_sums[13][112] [5:0] }), .sum({ \level_2_sums[13][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[229] [4:0] }), .sum({ \level_1_sums[13][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[231] [4:0] }), .sum({ \level_1_sums[13][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[13][115] [5:0] }),
     .b({ \level_1_sums[13][114] [5:0] }), .sum({ \level_2_sums[13][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[13][57] [6:0] }), .b({ \level_2_sums[13][56] [6:0] }), .sum({ \level_3_sums[13][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[233] [4:0] }), .sum({ \level_1_sums[13][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[235] [4:0] }), .sum({ \level_1_sums[13][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[13][117] [5:0] }),
     .b({ \level_1_sums[13][116] [5:0] }), .sum({ \level_2_sums[13][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[237] [4:0] }), .sum({ \level_1_sums[13][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[239] [4:0] }), .sum({ \level_1_sums[13][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[13][119] [5:0] }),
     .b({ \level_1_sums[13][118] [5:0] }), .sum({ \level_2_sums[13][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[13][59] [6:0] }), .b({ \level_2_sums[13][58] [6:0] }), .sum({ \level_3_sums[13][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[13][29] [7:0] }),
     .b({ \level_3_sums[13][28] [7:0] }), .sum({ \level_4_sums[13][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[241] [4:0] }), .sum({ \level_1_sums[13][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[243] [4:0] }), .sum({ \level_1_sums[13][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[13][121] [5:0] }),
     .b({ \level_1_sums[13][120] [5:0] }), .sum({ \level_2_sums[13][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[245] [4:0] }), .sum({ \level_1_sums[13][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[247] [4:0] }), .sum({ \level_1_sums[13][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[13][123] [5:0] }),
     .b({ \level_1_sums[13][122] [5:0] }), .sum({ \level_2_sums[13][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[13][61] [6:0] }), .b({ \level_2_sums[13][60] [6:0] }), .sum({ \level_3_sums[13][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[249] [4:0] }), .sum({ \level_1_sums[13][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[251] [4:0] }), .sum({ \level_1_sums[13][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[13][125] [5:0] }),
     .b({ \level_1_sums[13][124] [5:0] }), .sum({ \level_2_sums[13][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[253] [4:0] }), .sum({ \level_1_sums[13][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[13].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[13].product_terms[255] [4:0] }), .sum({ \level_1_sums[13][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[13][127] [5:0] }),
     .b({ \level_1_sums[13][126] [5:0] }), .sum({ \level_2_sums[13][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[13][63] [6:0] }), .b({ \level_2_sums[13][62] [6:0] }), .sum({ \level_3_sums[13][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[13][31] [7:0] }),
     .b({ \level_3_sums[13][30] [7:0] }), .sum({ \level_4_sums[13][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[13][15] [8:0] }),
     .b({ \level_4_sums[13][14] [8:0] }), .sum({ \level_5_sums[13][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[13][7] [9:0] }),
     .b({ \level_5_sums[13][6] [9:0] }), .sum({ \level_6_sums[13][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[13][3] [9:0] }),
     .b({ \level_6_sums[13][2] [9:0] }), .sum({ \level_7_sums[13][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[13].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[13][0] [9:0] }),
     .b({ \level_7_sums[13][1] [9:0] }), .sum({ \level_8_sums[13] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[14].relu_inst (.in_data({ \final_sums[14] [9:0] }), .out_data({ \out_sig[14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[1] [4:0] }), .sum({ \level_1_sums[14][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[3] [4:0] }), .sum({ \level_1_sums[14][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[14][1] [5:0] }),
     .b({ \level_1_sums[14][0] [5:0] }), .sum({ \level_2_sums[14][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[5] [4:0] }), .sum({ \level_1_sums[14][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[7] [4:0] }), .sum({ \level_1_sums[14][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[14][3] [5:0] }),
     .b({ \level_1_sums[14][2] [5:0] }), .sum({ \level_2_sums[14][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[14][1] [6:0] }),
     .b({ \level_2_sums[14][0] [6:0] }), .sum({ \level_3_sums[14][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[9] [4:0] }), .sum({ \level_1_sums[14][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[11] [4:0] }), .sum({ \level_1_sums[14][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[14][5] [5:0] }),
     .b({ \level_1_sums[14][4] [5:0] }), .sum({ \level_2_sums[14][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[13] [4:0] }), .sum({ \level_1_sums[14][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[15] [4:0] }), .sum({ \level_1_sums[14][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[14][7] [5:0] }),
     .b({ \level_1_sums[14][6] [5:0] }), .sum({ \level_2_sums[14][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[14][3] [6:0] }),
     .b({ \level_2_sums[14][2] [6:0] }), .sum({ \level_3_sums[14][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[14][1] [7:0] }),
     .b({ \level_3_sums[14][0] [7:0] }), .sum({ \level_4_sums[14][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[17] [4:0] }), .sum({ \level_1_sums[14][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[19] [4:0] }), .sum({ \level_1_sums[14][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[14][9] [5:0] }),
     .b({ \level_1_sums[14][8] [5:0] }), .sum({ \level_2_sums[14][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[21] [4:0] }), .sum({ \level_1_sums[14][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[23] [4:0] }), .sum({ \level_1_sums[14][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[14][11] [5:0] }),
     .b({ \level_1_sums[14][10] [5:0] }), .sum({ \level_2_sums[14][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[14][5] [6:0] }),
     .b({ \level_2_sums[14][4] [6:0] }), .sum({ \level_3_sums[14][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[25] [4:0] }), .sum({ \level_1_sums[14][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[27] [4:0] }), .sum({ \level_1_sums[14][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[14][13] [5:0] }),
     .b({ \level_1_sums[14][12] [5:0] }), .sum({ \level_2_sums[14][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[29] [4:0] }), .sum({ \level_1_sums[14][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[31] [4:0] }), .sum({ \level_1_sums[14][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[14][15] [5:0] }),
     .b({ \level_1_sums[14][14] [5:0] }), .sum({ \level_2_sums[14][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[14][7] [6:0] }),
     .b({ \level_2_sums[14][6] [6:0] }), .sum({ \level_3_sums[14][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[14][3] [7:0] }),
     .b({ \level_3_sums[14][2] [7:0] }), .sum({ \level_4_sums[14][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[14][1] [8:0] }),
     .b({ \level_4_sums[14][0] [8:0] }), .sum({ \level_5_sums[14][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[33] [4:0] }), .sum({ \level_1_sums[14][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[35] [4:0] }), .sum({ \level_1_sums[14][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[14][17] [5:0] }),
     .b({ \level_1_sums[14][16] [5:0] }), .sum({ \level_2_sums[14][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[37] [4:0] }), .sum({ \level_1_sums[14][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[39] [4:0] }), .sum({ \level_1_sums[14][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[14][19] [5:0] }),
     .b({ \level_1_sums[14][18] [5:0] }), .sum({ \level_2_sums[14][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[14][9] [6:0] }),
     .b({ \level_2_sums[14][8] [6:0] }), .sum({ \level_3_sums[14][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[41] [4:0] }), .sum({ \level_1_sums[14][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[43] [4:0] }), .sum({ \level_1_sums[14][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[14][21] [5:0] }),
     .b({ \level_1_sums[14][20] [5:0] }), .sum({ \level_2_sums[14][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[45] [4:0] }), .sum({ \level_1_sums[14][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[47] [4:0] }), .sum({ \level_1_sums[14][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[14][23] [5:0] }),
     .b({ \level_1_sums[14][22] [5:0] }), .sum({ \level_2_sums[14][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[14][11] [6:0] }),
     .b({ \level_2_sums[14][10] [6:0] }), .sum({ \level_3_sums[14][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[14][5] [7:0] }),
     .b({ \level_3_sums[14][4] [7:0] }), .sum({ \level_4_sums[14][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[49] [4:0] }), .sum({ \level_1_sums[14][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[51] [4:0] }), .sum({ \level_1_sums[14][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[14][25] [5:0] }),
     .b({ \level_1_sums[14][24] [5:0] }), .sum({ \level_2_sums[14][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[53] [4:0] }), .sum({ \level_1_sums[14][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[55] [4:0] }), .sum({ \level_1_sums[14][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[14][27] [5:0] }),
     .b({ \level_1_sums[14][26] [5:0] }), .sum({ \level_2_sums[14][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[14][13] [6:0] }),
     .b({ \level_2_sums[14][12] [6:0] }), .sum({ \level_3_sums[14][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[57] [4:0] }), .sum({ \level_1_sums[14][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[59] [4:0] }), .sum({ \level_1_sums[14][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[14][29] [5:0] }),
     .b({ \level_1_sums[14][28] [5:0] }), .sum({ \level_2_sums[14][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[61] [4:0] }), .sum({ \level_1_sums[14][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[63] [4:0] }), .sum({ \level_1_sums[14][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[14][31] [5:0] }),
     .b({ \level_1_sums[14][30] [5:0] }), .sum({ \level_2_sums[14][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[14][15] [6:0] }),
     .b({ \level_2_sums[14][14] [6:0] }), .sum({ \level_3_sums[14][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[14][7] [7:0] }),
     .b({ \level_3_sums[14][6] [7:0] }), .sum({ \level_4_sums[14][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[14][3] [8:0] }),
     .b({ \level_4_sums[14][2] [8:0] }), .sum({ \level_5_sums[14][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[14][1] [9:0] }),
     .b({ \level_5_sums[14][0] [9:0] }), .sum({ \level_6_sums[14][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[65] [4:0] }), .sum({ \level_1_sums[14][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[67] [4:0] }), .sum({ \level_1_sums[14][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[14][33] [5:0] }),
     .b({ \level_1_sums[14][32] [5:0] }), .sum({ \level_2_sums[14][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[69] [4:0] }), .sum({ \level_1_sums[14][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[71] [4:0] }), .sum({ \level_1_sums[14][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[14][35] [5:0] }),
     .b({ \level_1_sums[14][34] [5:0] }), .sum({ \level_2_sums[14][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[14][17] [6:0] }),
     .b({ \level_2_sums[14][16] [6:0] }), .sum({ \level_3_sums[14][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[73] [4:0] }), .sum({ \level_1_sums[14][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[75] [4:0] }), .sum({ \level_1_sums[14][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[14][37] [5:0] }),
     .b({ \level_1_sums[14][36] [5:0] }), .sum({ \level_2_sums[14][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[77] [4:0] }), .sum({ \level_1_sums[14][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[79] [4:0] }), .sum({ \level_1_sums[14][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[14][39] [5:0] }),
     .b({ \level_1_sums[14][38] [5:0] }), .sum({ \level_2_sums[14][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[14][19] [6:0] }),
     .b({ \level_2_sums[14][18] [6:0] }), .sum({ \level_3_sums[14][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[14][9] [7:0] }),
     .b({ \level_3_sums[14][8] [7:0] }), .sum({ \level_4_sums[14][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[81] [4:0] }), .sum({ \level_1_sums[14][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[83] [4:0] }), .sum({ \level_1_sums[14][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[14][41] [5:0] }),
     .b({ \level_1_sums[14][40] [5:0] }), .sum({ \level_2_sums[14][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[85] [4:0] }), .sum({ \level_1_sums[14][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[87] [4:0] }), .sum({ \level_1_sums[14][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[14][43] [5:0] }),
     .b({ \level_1_sums[14][42] [5:0] }), .sum({ \level_2_sums[14][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[14][21] [6:0] }),
     .b({ \level_2_sums[14][20] [6:0] }), .sum({ \level_3_sums[14][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[89] [4:0] }), .sum({ \level_1_sums[14][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[91] [4:0] }), .sum({ \level_1_sums[14][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[14][45] [5:0] }),
     .b({ \level_1_sums[14][44] [5:0] }), .sum({ \level_2_sums[14][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[93] [4:0] }), .sum({ \level_1_sums[14][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[95] [4:0] }), .sum({ \level_1_sums[14][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[14][47] [5:0] }),
     .b({ \level_1_sums[14][46] [5:0] }), .sum({ \level_2_sums[14][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[14][23] [6:0] }),
     .b({ \level_2_sums[14][22] [6:0] }), .sum({ \level_3_sums[14][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[14][11] [7:0] }),
     .b({ \level_3_sums[14][10] [7:0] }), .sum({ \level_4_sums[14][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[14][5] [8:0] }),
     .b({ \level_4_sums[14][4] [8:0] }), .sum({ \level_5_sums[14][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[97] [4:0] }), .sum({ \level_1_sums[14][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[99] [4:0] }), .sum({ \level_1_sums[14][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[14][49] [5:0] }),
     .b({ \level_1_sums[14][48] [5:0] }), .sum({ \level_2_sums[14][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[101] [4:0] }), .sum({ \level_1_sums[14][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[103] [4:0] }), .sum({ \level_1_sums[14][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[14][51] [5:0] }),
     .b({ \level_1_sums[14][50] [5:0] }), .sum({ \level_2_sums[14][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[14][25] [6:0] }), .b({ \level_2_sums[14][24] [6:0] }), .sum({ \level_3_sums[14][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[105] [4:0] }), .sum({ \level_1_sums[14][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[107] [4:0] }), .sum({ \level_1_sums[14][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[14][53] [5:0] }),
     .b({ \level_1_sums[14][52] [5:0] }), .sum({ \level_2_sums[14][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[109] [4:0] }), .sum({ \level_1_sums[14][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[111] [4:0] }), .sum({ \level_1_sums[14][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[14][55] [5:0] }),
     .b({ \level_1_sums[14][54] [5:0] }), .sum({ \level_2_sums[14][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[14][27] [6:0] }), .b({ \level_2_sums[14][26] [6:0] }), .sum({ \level_3_sums[14][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[14][13] [7:0] }),
     .b({ \level_3_sums[14][12] [7:0] }), .sum({ \level_4_sums[14][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[113] [4:0] }), .sum({ \level_1_sums[14][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[115] [4:0] }), .sum({ \level_1_sums[14][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[14][57] [5:0] }),
     .b({ \level_1_sums[14][56] [5:0] }), .sum({ \level_2_sums[14][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[117] [4:0] }), .sum({ \level_1_sums[14][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[119] [4:0] }), .sum({ \level_1_sums[14][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[14][59] [5:0] }),
     .b({ \level_1_sums[14][58] [5:0] }), .sum({ \level_2_sums[14][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[14][29] [6:0] }), .b({ \level_2_sums[14][28] [6:0] }), .sum({ \level_3_sums[14][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[121] [4:0] }), .sum({ \level_1_sums[14][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[123] [4:0] }), .sum({ \level_1_sums[14][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[14][61] [5:0] }),
     .b({ \level_1_sums[14][60] [5:0] }), .sum({ \level_2_sums[14][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[125] [4:0] }), .sum({ \level_1_sums[14][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[127] [4:0] }), .sum({ \level_1_sums[14][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[14][63] [5:0] }),
     .b({ \level_1_sums[14][62] [5:0] }), .sum({ \level_2_sums[14][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[14][31] [6:0] }), .b({ \level_2_sums[14][30] [6:0] }), .sum({ \level_3_sums[14][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[14][15] [7:0] }),
     .b({ \level_3_sums[14][14] [7:0] }), .sum({ \level_4_sums[14][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[14][7] [8:0] }),
     .b({ \level_4_sums[14][6] [8:0] }), .sum({ \level_5_sums[14][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[14][3] [9:0] }),
     .b({ \level_5_sums[14][2] [9:0] }), .sum({ \level_6_sums[14][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[14][1] [9:0] }),
     .b({ \level_6_sums[14][0] [9:0] }), .sum({ \level_7_sums[14][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[129] [4:0] }), .sum({ \level_1_sums[14][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[131] [4:0] }), .sum({ \level_1_sums[14][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[14][65] [5:0] }),
     .b({ \level_1_sums[14][64] [5:0] }), .sum({ \level_2_sums[14][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[133] [4:0] }), .sum({ \level_1_sums[14][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[135] [4:0] }), .sum({ \level_1_sums[14][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[14][67] [5:0] }),
     .b({ \level_1_sums[14][66] [5:0] }), .sum({ \level_2_sums[14][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[14][33] [6:0] }), .b({ \level_2_sums[14][32] [6:0] }), .sum({ \level_3_sums[14][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[137] [4:0] }), .sum({ \level_1_sums[14][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[139] [4:0] }), .sum({ \level_1_sums[14][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[14][69] [5:0] }),
     .b({ \level_1_sums[14][68] [5:0] }), .sum({ \level_2_sums[14][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[141] [4:0] }), .sum({ \level_1_sums[14][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[143] [4:0] }), .sum({ \level_1_sums[14][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[14][71] [5:0] }),
     .b({ \level_1_sums[14][70] [5:0] }), .sum({ \level_2_sums[14][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[14][35] [6:0] }), .b({ \level_2_sums[14][34] [6:0] }), .sum({ \level_3_sums[14][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[14][17] [7:0] }),
     .b({ \level_3_sums[14][16] [7:0] }), .sum({ \level_4_sums[14][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[145] [4:0] }), .sum({ \level_1_sums[14][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[147] [4:0] }), .sum({ \level_1_sums[14][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[14][73] [5:0] }),
     .b({ \level_1_sums[14][72] [5:0] }), .sum({ \level_2_sums[14][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[149] [4:0] }), .sum({ \level_1_sums[14][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[151] [4:0] }), .sum({ \level_1_sums[14][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[14][75] [5:0] }),
     .b({ \level_1_sums[14][74] [5:0] }), .sum({ \level_2_sums[14][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[14][37] [6:0] }), .b({ \level_2_sums[14][36] [6:0] }), .sum({ \level_3_sums[14][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[153] [4:0] }), .sum({ \level_1_sums[14][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[155] [4:0] }), .sum({ \level_1_sums[14][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[14][77] [5:0] }),
     .b({ \level_1_sums[14][76] [5:0] }), .sum({ \level_2_sums[14][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[157] [4:0] }), .sum({ \level_1_sums[14][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[159] [4:0] }), .sum({ \level_1_sums[14][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[14][79] [5:0] }),
     .b({ \level_1_sums[14][78] [5:0] }), .sum({ \level_2_sums[14][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[14][39] [6:0] }), .b({ \level_2_sums[14][38] [6:0] }), .sum({ \level_3_sums[14][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[14][19] [7:0] }),
     .b({ \level_3_sums[14][18] [7:0] }), .sum({ \level_4_sums[14][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[14][9] [8:0] }),
     .b({ \level_4_sums[14][8] [8:0] }), .sum({ \level_5_sums[14][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[161] [4:0] }), .sum({ \level_1_sums[14][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[163] [4:0] }), .sum({ \level_1_sums[14][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[14][81] [5:0] }),
     .b({ \level_1_sums[14][80] [5:0] }), .sum({ \level_2_sums[14][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[165] [4:0] }), .sum({ \level_1_sums[14][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[167] [4:0] }), .sum({ \level_1_sums[14][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[14][83] [5:0] }),
     .b({ \level_1_sums[14][82] [5:0] }), .sum({ \level_2_sums[14][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[14][41] [6:0] }), .b({ \level_2_sums[14][40] [6:0] }), .sum({ \level_3_sums[14][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[169] [4:0] }), .sum({ \level_1_sums[14][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[171] [4:0] }), .sum({ \level_1_sums[14][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[14][85] [5:0] }),
     .b({ \level_1_sums[14][84] [5:0] }), .sum({ \level_2_sums[14][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[173] [4:0] }), .sum({ \level_1_sums[14][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[175] [4:0] }), .sum({ \level_1_sums[14][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[14][87] [5:0] }),
     .b({ \level_1_sums[14][86] [5:0] }), .sum({ \level_2_sums[14][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[14][43] [6:0] }), .b({ \level_2_sums[14][42] [6:0] }), .sum({ \level_3_sums[14][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[14][21] [7:0] }),
     .b({ \level_3_sums[14][20] [7:0] }), .sum({ \level_4_sums[14][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[177] [4:0] }), .sum({ \level_1_sums[14][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[179] [4:0] }), .sum({ \level_1_sums[14][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[14][89] [5:0] }),
     .b({ \level_1_sums[14][88] [5:0] }), .sum({ \level_2_sums[14][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[181] [4:0] }), .sum({ \level_1_sums[14][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[183] [4:0] }), .sum({ \level_1_sums[14][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[14][91] [5:0] }),
     .b({ \level_1_sums[14][90] [5:0] }), .sum({ \level_2_sums[14][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[14][45] [6:0] }), .b({ \level_2_sums[14][44] [6:0] }), .sum({ \level_3_sums[14][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[185] [4:0] }), .sum({ \level_1_sums[14][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[187] [4:0] }), .sum({ \level_1_sums[14][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[14][93] [5:0] }),
     .b({ \level_1_sums[14][92] [5:0] }), .sum({ \level_2_sums[14][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[189] [4:0] }), .sum({ \level_1_sums[14][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[191] [4:0] }), .sum({ \level_1_sums[14][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[14][95] [5:0] }),
     .b({ \level_1_sums[14][94] [5:0] }), .sum({ \level_2_sums[14][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[14][47] [6:0] }), .b({ \level_2_sums[14][46] [6:0] }), .sum({ \level_3_sums[14][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[14][23] [7:0] }),
     .b({ \level_3_sums[14][22] [7:0] }), .sum({ \level_4_sums[14][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[14][11] [8:0] }),
     .b({ \level_4_sums[14][10] [8:0] }), .sum({ \level_5_sums[14][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[14][5] [9:0] }),
     .b({ \level_5_sums[14][4] [9:0] }), .sum({ \level_6_sums[14][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[193] [4:0] }), .sum({ \level_1_sums[14][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[195] [4:0] }), .sum({ \level_1_sums[14][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[14][97] [5:0] }),
     .b({ \level_1_sums[14][96] [5:0] }), .sum({ \level_2_sums[14][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[197] [4:0] }), .sum({ \level_1_sums[14][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[199] [4:0] }), .sum({ \level_1_sums[14][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[14][99] [5:0] }),
     .b({ \level_1_sums[14][98] [5:0] }), .sum({ \level_2_sums[14][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[14][49] [6:0] }), .b({ \level_2_sums[14][48] [6:0] }), .sum({ \level_3_sums[14][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[201] [4:0] }), .sum({ \level_1_sums[14][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[203] [4:0] }), .sum({ \level_1_sums[14][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[14][101] [5:0] }),
     .b({ \level_1_sums[14][100] [5:0] }), .sum({ \level_2_sums[14][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[205] [4:0] }), .sum({ \level_1_sums[14][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[207] [4:0] }), .sum({ \level_1_sums[14][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[14][103] [5:0] }),
     .b({ \level_1_sums[14][102] [5:0] }), .sum({ \level_2_sums[14][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[14][51] [6:0] }), .b({ \level_2_sums[14][50] [6:0] }), .sum({ \level_3_sums[14][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[14][25] [7:0] }),
     .b({ \level_3_sums[14][24] [7:0] }), .sum({ \level_4_sums[14][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[209] [4:0] }), .sum({ \level_1_sums[14][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[211] [4:0] }), .sum({ \level_1_sums[14][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[14][105] [5:0] }),
     .b({ \level_1_sums[14][104] [5:0] }), .sum({ \level_2_sums[14][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[213] [4:0] }), .sum({ \level_1_sums[14][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[215] [4:0] }), .sum({ \level_1_sums[14][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[14][107] [5:0] }),
     .b({ \level_1_sums[14][106] [5:0] }), .sum({ \level_2_sums[14][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[14][53] [6:0] }), .b({ \level_2_sums[14][52] [6:0] }), .sum({ \level_3_sums[14][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[217] [4:0] }), .sum({ \level_1_sums[14][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[219] [4:0] }), .sum({ \level_1_sums[14][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[14][109] [5:0] }),
     .b({ \level_1_sums[14][108] [5:0] }), .sum({ \level_2_sums[14][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[221] [4:0] }), .sum({ \level_1_sums[14][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[223] [4:0] }), .sum({ \level_1_sums[14][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[14][111] [5:0] }),
     .b({ \level_1_sums[14][110] [5:0] }), .sum({ \level_2_sums[14][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[14][55] [6:0] }), .b({ \level_2_sums[14][54] [6:0] }), .sum({ \level_3_sums[14][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[14][27] [7:0] }),
     .b({ \level_3_sums[14][26] [7:0] }), .sum({ \level_4_sums[14][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[14][13] [8:0] }),
     .b({ \level_4_sums[14][12] [8:0] }), .sum({ \level_5_sums[14][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[225] [4:0] }), .sum({ \level_1_sums[14][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[227] [4:0] }), .sum({ \level_1_sums[14][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[14][113] [5:0] }),
     .b({ \level_1_sums[14][112] [5:0] }), .sum({ \level_2_sums[14][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[229] [4:0] }), .sum({ \level_1_sums[14][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[231] [4:0] }), .sum({ \level_1_sums[14][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[14][115] [5:0] }),
     .b({ \level_1_sums[14][114] [5:0] }), .sum({ \level_2_sums[14][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[14][57] [6:0] }), .b({ \level_2_sums[14][56] [6:0] }), .sum({ \level_3_sums[14][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[233] [4:0] }), .sum({ \level_1_sums[14][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[235] [4:0] }), .sum({ \level_1_sums[14][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[14][117] [5:0] }),
     .b({ \level_1_sums[14][116] [5:0] }), .sum({ \level_2_sums[14][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[237] [4:0] }), .sum({ \level_1_sums[14][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[239] [4:0] }), .sum({ \level_1_sums[14][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[14][119] [5:0] }),
     .b({ \level_1_sums[14][118] [5:0] }), .sum({ \level_2_sums[14][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[14][59] [6:0] }), .b({ \level_2_sums[14][58] [6:0] }), .sum({ \level_3_sums[14][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[14][29] [7:0] }),
     .b({ \level_3_sums[14][28] [7:0] }), .sum({ \level_4_sums[14][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[241] [4:0] }), .sum({ \level_1_sums[14][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[243] [4:0] }), .sum({ \level_1_sums[14][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[14][121] [5:0] }),
     .b({ \level_1_sums[14][120] [5:0] }), .sum({ \level_2_sums[14][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[245] [4:0] }), .sum({ \level_1_sums[14][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[247] [4:0] }), .sum({ \level_1_sums[14][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[14][123] [5:0] }),
     .b({ \level_1_sums[14][122] [5:0] }), .sum({ \level_2_sums[14][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[14][61] [6:0] }), .b({ \level_2_sums[14][60] [6:0] }), .sum({ \level_3_sums[14][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[249] [4:0] }), .sum({ \level_1_sums[14][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[251] [4:0] }), .sum({ \level_1_sums[14][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[14][125] [5:0] }),
     .b({ \level_1_sums[14][124] [5:0] }), .sum({ \level_2_sums[14][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[253] [4:0] }), .sum({ \level_1_sums[14][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[14].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[14].product_terms[255] [4:0] }), .sum({ \level_1_sums[14][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[14][127] [5:0] }),
     .b({ \level_1_sums[14][126] [5:0] }), .sum({ \level_2_sums[14][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[14][63] [6:0] }), .b({ \level_2_sums[14][62] [6:0] }), .sum({ \level_3_sums[14][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[14][31] [7:0] }),
     .b({ \level_3_sums[14][30] [7:0] }), .sum({ \level_4_sums[14][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[14][15] [8:0] }),
     .b({ \level_4_sums[14][14] [8:0] }), .sum({ \level_5_sums[14][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[14][7] [9:0] }),
     .b({ \level_5_sums[14][6] [9:0] }), .sum({ \level_6_sums[14][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[14][3] [9:0] }),
     .b({ \level_6_sums[14][2] [9:0] }), .sum({ \level_7_sums[14][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[14].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[14][0] [9:0] }),
     .b({ \level_7_sums[14][1] [9:0] }), .sum({ \level_8_sums[14] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[15].relu_inst (.in_data({ \final_sums[15] [9:0] }), .out_data({ \out_sig[15] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[1] [4:0] }), .sum({ \level_1_sums[15][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[3] [4:0] }), .sum({ \level_1_sums[15][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[15][1] [5:0] }),
     .b({ \level_1_sums[15][0] [5:0] }), .sum({ \level_2_sums[15][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[5] [4:0] }), .sum({ \level_1_sums[15][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[7] [4:0] }), .sum({ \level_1_sums[15][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[15][3] [5:0] }),
     .b({ \level_1_sums[15][2] [5:0] }), .sum({ \level_2_sums[15][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[15][1] [6:0] }),
     .b({ \level_2_sums[15][0] [6:0] }), .sum({ \level_3_sums[15][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[9] [4:0] }), .sum({ \level_1_sums[15][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[11] [4:0] }), .sum({ \level_1_sums[15][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[15][5] [5:0] }),
     .b({ \level_1_sums[15][4] [5:0] }), .sum({ \level_2_sums[15][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[13] [4:0] }), .sum({ \level_1_sums[15][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[15] [4:0] }), .sum({ \level_1_sums[15][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[15][7] [5:0] }),
     .b({ \level_1_sums[15][6] [5:0] }), .sum({ \level_2_sums[15][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[15][3] [6:0] }),
     .b({ \level_2_sums[15][2] [6:0] }), .sum({ \level_3_sums[15][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[15][1] [7:0] }),
     .b({ \level_3_sums[15][0] [7:0] }), .sum({ \level_4_sums[15][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[17] [4:0] }), .sum({ \level_1_sums[15][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[19] [4:0] }), .sum({ \level_1_sums[15][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[15][9] [5:0] }),
     .b({ \level_1_sums[15][8] [5:0] }), .sum({ \level_2_sums[15][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[21] [4:0] }), .sum({ \level_1_sums[15][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[23] [4:0] }), .sum({ \level_1_sums[15][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[15][11] [5:0] }),
     .b({ \level_1_sums[15][10] [5:0] }), .sum({ \level_2_sums[15][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[15][5] [6:0] }),
     .b({ \level_2_sums[15][4] [6:0] }), .sum({ \level_3_sums[15][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[25] [4:0] }), .sum({ \level_1_sums[15][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[27] [4:0] }), .sum({ \level_1_sums[15][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[15][13] [5:0] }),
     .b({ \level_1_sums[15][12] [5:0] }), .sum({ \level_2_sums[15][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[29] [4:0] }), .sum({ \level_1_sums[15][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[31] [4:0] }), .sum({ \level_1_sums[15][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[15][15] [5:0] }),
     .b({ \level_1_sums[15][14] [5:0] }), .sum({ \level_2_sums[15][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[15][7] [6:0] }),
     .b({ \level_2_sums[15][6] [6:0] }), .sum({ \level_3_sums[15][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[15][3] [7:0] }),
     .b({ \level_3_sums[15][2] [7:0] }), .sum({ \level_4_sums[15][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[15][1] [8:0] }),
     .b({ \level_4_sums[15][0] [8:0] }), .sum({ \level_5_sums[15][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[33] [4:0] }), .sum({ \level_1_sums[15][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[35] [4:0] }), .sum({ \level_1_sums[15][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[15][17] [5:0] }),
     .b({ \level_1_sums[15][16] [5:0] }), .sum({ \level_2_sums[15][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[37] [4:0] }), .sum({ \level_1_sums[15][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[39] [4:0] }), .sum({ \level_1_sums[15][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[15][19] [5:0] }),
     .b({ \level_1_sums[15][18] [5:0] }), .sum({ \level_2_sums[15][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[15][9] [6:0] }),
     .b({ \level_2_sums[15][8] [6:0] }), .sum({ \level_3_sums[15][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[41] [4:0] }), .sum({ \level_1_sums[15][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[43] [4:0] }), .sum({ \level_1_sums[15][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[15][21] [5:0] }),
     .b({ \level_1_sums[15][20] [5:0] }), .sum({ \level_2_sums[15][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[45] [4:0] }), .sum({ \level_1_sums[15][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[47] [4:0] }), .sum({ \level_1_sums[15][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[15][23] [5:0] }),
     .b({ \level_1_sums[15][22] [5:0] }), .sum({ \level_2_sums[15][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[15][11] [6:0] }),
     .b({ \level_2_sums[15][10] [6:0] }), .sum({ \level_3_sums[15][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[15][5] [7:0] }),
     .b({ \level_3_sums[15][4] [7:0] }), .sum({ \level_4_sums[15][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[49] [4:0] }), .sum({ \level_1_sums[15][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[51] [4:0] }), .sum({ \level_1_sums[15][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[15][25] [5:0] }),
     .b({ \level_1_sums[15][24] [5:0] }), .sum({ \level_2_sums[15][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[53] [4:0] }), .sum({ \level_1_sums[15][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[55] [4:0] }), .sum({ \level_1_sums[15][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[15][27] [5:0] }),
     .b({ \level_1_sums[15][26] [5:0] }), .sum({ \level_2_sums[15][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[15][13] [6:0] }),
     .b({ \level_2_sums[15][12] [6:0] }), .sum({ \level_3_sums[15][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[57] [4:0] }), .sum({ \level_1_sums[15][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[59] [4:0] }), .sum({ \level_1_sums[15][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[15][29] [5:0] }),
     .b({ \level_1_sums[15][28] [5:0] }), .sum({ \level_2_sums[15][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[61] [4:0] }), .sum({ \level_1_sums[15][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[63] [4:0] }), .sum({ \level_1_sums[15][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[15][31] [5:0] }),
     .b({ \level_1_sums[15][30] [5:0] }), .sum({ \level_2_sums[15][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[15][15] [6:0] }),
     .b({ \level_2_sums[15][14] [6:0] }), .sum({ \level_3_sums[15][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[15][7] [7:0] }),
     .b({ \level_3_sums[15][6] [7:0] }), .sum({ \level_4_sums[15][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[15][3] [8:0] }),
     .b({ \level_4_sums[15][2] [8:0] }), .sum({ \level_5_sums[15][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[15][1] [9:0] }),
     .b({ \level_5_sums[15][0] [9:0] }), .sum({ \level_6_sums[15][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[65] [4:0] }), .sum({ \level_1_sums[15][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[67] [4:0] }), .sum({ \level_1_sums[15][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[15][33] [5:0] }),
     .b({ \level_1_sums[15][32] [5:0] }), .sum({ \level_2_sums[15][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[69] [4:0] }), .sum({ \level_1_sums[15][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[71] [4:0] }), .sum({ \level_1_sums[15][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[15][35] [5:0] }),
     .b({ \level_1_sums[15][34] [5:0] }), .sum({ \level_2_sums[15][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[15][17] [6:0] }),
     .b({ \level_2_sums[15][16] [6:0] }), .sum({ \level_3_sums[15][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[73] [4:0] }), .sum({ \level_1_sums[15][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[75] [4:0] }), .sum({ \level_1_sums[15][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[15][37] [5:0] }),
     .b({ \level_1_sums[15][36] [5:0] }), .sum({ \level_2_sums[15][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[77] [4:0] }), .sum({ \level_1_sums[15][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[79] [4:0] }), .sum({ \level_1_sums[15][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[15][39] [5:0] }),
     .b({ \level_1_sums[15][38] [5:0] }), .sum({ \level_2_sums[15][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[15][19] [6:0] }),
     .b({ \level_2_sums[15][18] [6:0] }), .sum({ \level_3_sums[15][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[15][9] [7:0] }),
     .b({ \level_3_sums[15][8] [7:0] }), .sum({ \level_4_sums[15][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[81] [4:0] }), .sum({ \level_1_sums[15][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[83] [4:0] }), .sum({ \level_1_sums[15][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[15][41] [5:0] }),
     .b({ \level_1_sums[15][40] [5:0] }), .sum({ \level_2_sums[15][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[85] [4:0] }), .sum({ \level_1_sums[15][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[87] [4:0] }), .sum({ \level_1_sums[15][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[15][43] [5:0] }),
     .b({ \level_1_sums[15][42] [5:0] }), .sum({ \level_2_sums[15][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[15][21] [6:0] }),
     .b({ \level_2_sums[15][20] [6:0] }), .sum({ \level_3_sums[15][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[89] [4:0] }), .sum({ \level_1_sums[15][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[91] [4:0] }), .sum({ \level_1_sums[15][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[15][45] [5:0] }),
     .b({ \level_1_sums[15][44] [5:0] }), .sum({ \level_2_sums[15][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[93] [4:0] }), .sum({ \level_1_sums[15][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[95] [4:0] }), .sum({ \level_1_sums[15][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[15][47] [5:0] }),
     .b({ \level_1_sums[15][46] [5:0] }), .sum({ \level_2_sums[15][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[15][23] [6:0] }),
     .b({ \level_2_sums[15][22] [6:0] }), .sum({ \level_3_sums[15][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[15][11] [7:0] }),
     .b({ \level_3_sums[15][10] [7:0] }), .sum({ \level_4_sums[15][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[15][5] [8:0] }),
     .b({ \level_4_sums[15][4] [8:0] }), .sum({ \level_5_sums[15][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[97] [4:0] }), .sum({ \level_1_sums[15][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[99] [4:0] }), .sum({ \level_1_sums[15][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[15][49] [5:0] }),
     .b({ \level_1_sums[15][48] [5:0] }), .sum({ \level_2_sums[15][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[101] [4:0] }), .sum({ \level_1_sums[15][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[103] [4:0] }), .sum({ \level_1_sums[15][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[15][51] [5:0] }),
     .b({ \level_1_sums[15][50] [5:0] }), .sum({ \level_2_sums[15][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[15][25] [6:0] }), .b({ \level_2_sums[15][24] [6:0] }), .sum({ \level_3_sums[15][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[105] [4:0] }), .sum({ \level_1_sums[15][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[107] [4:0] }), .sum({ \level_1_sums[15][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[15][53] [5:0] }),
     .b({ \level_1_sums[15][52] [5:0] }), .sum({ \level_2_sums[15][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[109] [4:0] }), .sum({ \level_1_sums[15][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[111] [4:0] }), .sum({ \level_1_sums[15][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[15][55] [5:0] }),
     .b({ \level_1_sums[15][54] [5:0] }), .sum({ \level_2_sums[15][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[15][27] [6:0] }), .b({ \level_2_sums[15][26] [6:0] }), .sum({ \level_3_sums[15][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[15][13] [7:0] }),
     .b({ \level_3_sums[15][12] [7:0] }), .sum({ \level_4_sums[15][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[113] [4:0] }), .sum({ \level_1_sums[15][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[115] [4:0] }), .sum({ \level_1_sums[15][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[15][57] [5:0] }),
     .b({ \level_1_sums[15][56] [5:0] }), .sum({ \level_2_sums[15][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[117] [4:0] }), .sum({ \level_1_sums[15][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[119] [4:0] }), .sum({ \level_1_sums[15][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[15][59] [5:0] }),
     .b({ \level_1_sums[15][58] [5:0] }), .sum({ \level_2_sums[15][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[15][29] [6:0] }), .b({ \level_2_sums[15][28] [6:0] }), .sum({ \level_3_sums[15][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[121] [4:0] }), .sum({ \level_1_sums[15][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[123] [4:0] }), .sum({ \level_1_sums[15][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[15][61] [5:0] }),
     .b({ \level_1_sums[15][60] [5:0] }), .sum({ \level_2_sums[15][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[125] [4:0] }), .sum({ \level_1_sums[15][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[127] [4:0] }), .sum({ \level_1_sums[15][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[15][63] [5:0] }),
     .b({ \level_1_sums[15][62] [5:0] }), .sum({ \level_2_sums[15][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[15][31] [6:0] }), .b({ \level_2_sums[15][30] [6:0] }), .sum({ \level_3_sums[15][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[15][15] [7:0] }),
     .b({ \level_3_sums[15][14] [7:0] }), .sum({ \level_4_sums[15][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[15][7] [8:0] }),
     .b({ \level_4_sums[15][6] [8:0] }), .sum({ \level_5_sums[15][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[15][3] [9:0] }),
     .b({ \level_5_sums[15][2] [9:0] }), .sum({ \level_6_sums[15][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[15][1] [9:0] }),
     .b({ \level_6_sums[15][0] [9:0] }), .sum({ \level_7_sums[15][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[129] [4:0] }), .sum({ \level_1_sums[15][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[131] [4:0] }), .sum({ \level_1_sums[15][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[15][65] [5:0] }),
     .b({ \level_1_sums[15][64] [5:0] }), .sum({ \level_2_sums[15][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[133] [4:0] }), .sum({ \level_1_sums[15][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[135] [4:0] }), .sum({ \level_1_sums[15][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[15][67] [5:0] }),
     .b({ \level_1_sums[15][66] [5:0] }), .sum({ \level_2_sums[15][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[15][33] [6:0] }), .b({ \level_2_sums[15][32] [6:0] }), .sum({ \level_3_sums[15][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[137] [4:0] }), .sum({ \level_1_sums[15][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[139] [4:0] }), .sum({ \level_1_sums[15][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[15][69] [5:0] }),
     .b({ \level_1_sums[15][68] [5:0] }), .sum({ \level_2_sums[15][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[141] [4:0] }), .sum({ \level_1_sums[15][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[143] [4:0] }), .sum({ \level_1_sums[15][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[15][71] [5:0] }),
     .b({ \level_1_sums[15][70] [5:0] }), .sum({ \level_2_sums[15][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[15][35] [6:0] }), .b({ \level_2_sums[15][34] [6:0] }), .sum({ \level_3_sums[15][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[15][17] [7:0] }),
     .b({ \level_3_sums[15][16] [7:0] }), .sum({ \level_4_sums[15][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[145] [4:0] }), .sum({ \level_1_sums[15][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[147] [4:0] }), .sum({ \level_1_sums[15][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[15][73] [5:0] }),
     .b({ \level_1_sums[15][72] [5:0] }), .sum({ \level_2_sums[15][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[149] [4:0] }), .sum({ \level_1_sums[15][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[151] [4:0] }), .sum({ \level_1_sums[15][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[15][75] [5:0] }),
     .b({ \level_1_sums[15][74] [5:0] }), .sum({ \level_2_sums[15][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[15][37] [6:0] }), .b({ \level_2_sums[15][36] [6:0] }), .sum({ \level_3_sums[15][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[153] [4:0] }), .sum({ \level_1_sums[15][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[155] [4:0] }), .sum({ \level_1_sums[15][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[15][77] [5:0] }),
     .b({ \level_1_sums[15][76] [5:0] }), .sum({ \level_2_sums[15][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[157] [4:0] }), .sum({ \level_1_sums[15][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[159] [4:0] }), .sum({ \level_1_sums[15][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[15][79] [5:0] }),
     .b({ \level_1_sums[15][78] [5:0] }), .sum({ \level_2_sums[15][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[15][39] [6:0] }), .b({ \level_2_sums[15][38] [6:0] }), .sum({ \level_3_sums[15][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[15][19] [7:0] }),
     .b({ \level_3_sums[15][18] [7:0] }), .sum({ \level_4_sums[15][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[15][9] [8:0] }),
     .b({ \level_4_sums[15][8] [8:0] }), .sum({ \level_5_sums[15][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[161] [4:0] }), .sum({ \level_1_sums[15][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[163] [4:0] }), .sum({ \level_1_sums[15][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[15][81] [5:0] }),
     .b({ \level_1_sums[15][80] [5:0] }), .sum({ \level_2_sums[15][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[165] [4:0] }), .sum({ \level_1_sums[15][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[167] [4:0] }), .sum({ \level_1_sums[15][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[15][83] [5:0] }),
     .b({ \level_1_sums[15][82] [5:0] }), .sum({ \level_2_sums[15][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[15][41] [6:0] }), .b({ \level_2_sums[15][40] [6:0] }), .sum({ \level_3_sums[15][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[169] [4:0] }), .sum({ \level_1_sums[15][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[171] [4:0] }), .sum({ \level_1_sums[15][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[15][85] [5:0] }),
     .b({ \level_1_sums[15][84] [5:0] }), .sum({ \level_2_sums[15][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[173] [4:0] }), .sum({ \level_1_sums[15][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[175] [4:0] }), .sum({ \level_1_sums[15][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[15][87] [5:0] }),
     .b({ \level_1_sums[15][86] [5:0] }), .sum({ \level_2_sums[15][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[15][43] [6:0] }), .b({ \level_2_sums[15][42] [6:0] }), .sum({ \level_3_sums[15][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[15][21] [7:0] }),
     .b({ \level_3_sums[15][20] [7:0] }), .sum({ \level_4_sums[15][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[177] [4:0] }), .sum({ \level_1_sums[15][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[179] [4:0] }), .sum({ \level_1_sums[15][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[15][89] [5:0] }),
     .b({ \level_1_sums[15][88] [5:0] }), .sum({ \level_2_sums[15][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[181] [4:0] }), .sum({ \level_1_sums[15][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[183] [4:0] }), .sum({ \level_1_sums[15][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[15][91] [5:0] }),
     .b({ \level_1_sums[15][90] [5:0] }), .sum({ \level_2_sums[15][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[15][45] [6:0] }), .b({ \level_2_sums[15][44] [6:0] }), .sum({ \level_3_sums[15][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[185] [4:0] }), .sum({ \level_1_sums[15][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[187] [4:0] }), .sum({ \level_1_sums[15][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[15][93] [5:0] }),
     .b({ \level_1_sums[15][92] [5:0] }), .sum({ \level_2_sums[15][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[189] [4:0] }), .sum({ \level_1_sums[15][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[191] [4:0] }), .sum({ \level_1_sums[15][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[15][95] [5:0] }),
     .b({ \level_1_sums[15][94] [5:0] }), .sum({ \level_2_sums[15][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[15][47] [6:0] }), .b({ \level_2_sums[15][46] [6:0] }), .sum({ \level_3_sums[15][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[15][23] [7:0] }),
     .b({ \level_3_sums[15][22] [7:0] }), .sum({ \level_4_sums[15][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[15][11] [8:0] }),
     .b({ \level_4_sums[15][10] [8:0] }), .sum({ \level_5_sums[15][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[15][5] [9:0] }),
     .b({ \level_5_sums[15][4] [9:0] }), .sum({ \level_6_sums[15][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[193] [4:0] }), .sum({ \level_1_sums[15][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[195] [4:0] }), .sum({ \level_1_sums[15][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[15][97] [5:0] }),
     .b({ \level_1_sums[15][96] [5:0] }), .sum({ \level_2_sums[15][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[197] [4:0] }), .sum({ \level_1_sums[15][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[199] [4:0] }), .sum({ \level_1_sums[15][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[15][99] [5:0] }),
     .b({ \level_1_sums[15][98] [5:0] }), .sum({ \level_2_sums[15][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[15][49] [6:0] }), .b({ \level_2_sums[15][48] [6:0] }), .sum({ \level_3_sums[15][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[201] [4:0] }), .sum({ \level_1_sums[15][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[203] [4:0] }), .sum({ \level_1_sums[15][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[15][101] [5:0] }),
     .b({ \level_1_sums[15][100] [5:0] }), .sum({ \level_2_sums[15][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[205] [4:0] }), .sum({ \level_1_sums[15][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[207] [4:0] }), .sum({ \level_1_sums[15][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[15][103] [5:0] }),
     .b({ \level_1_sums[15][102] [5:0] }), .sum({ \level_2_sums[15][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[15][51] [6:0] }), .b({ \level_2_sums[15][50] [6:0] }), .sum({ \level_3_sums[15][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[15][25] [7:0] }),
     .b({ \level_3_sums[15][24] [7:0] }), .sum({ \level_4_sums[15][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[209] [4:0] }), .sum({ \level_1_sums[15][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[211] [4:0] }), .sum({ \level_1_sums[15][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[15][105] [5:0] }),
     .b({ \level_1_sums[15][104] [5:0] }), .sum({ \level_2_sums[15][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[213] [4:0] }), .sum({ \level_1_sums[15][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[215] [4:0] }), .sum({ \level_1_sums[15][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[15][107] [5:0] }),
     .b({ \level_1_sums[15][106] [5:0] }), .sum({ \level_2_sums[15][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[15][53] [6:0] }), .b({ \level_2_sums[15][52] [6:0] }), .sum({ \level_3_sums[15][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[217] [4:0] }), .sum({ \level_1_sums[15][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[219] [4:0] }), .sum({ \level_1_sums[15][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[15][109] [5:0] }),
     .b({ \level_1_sums[15][108] [5:0] }), .sum({ \level_2_sums[15][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[221] [4:0] }), .sum({ \level_1_sums[15][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[223] [4:0] }), .sum({ \level_1_sums[15][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[15][111] [5:0] }),
     .b({ \level_1_sums[15][110] [5:0] }), .sum({ \level_2_sums[15][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[15][55] [6:0] }), .b({ \level_2_sums[15][54] [6:0] }), .sum({ \level_3_sums[15][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[15][27] [7:0] }),
     .b({ \level_3_sums[15][26] [7:0] }), .sum({ \level_4_sums[15][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[15][13] [8:0] }),
     .b({ \level_4_sums[15][12] [8:0] }), .sum({ \level_5_sums[15][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[225] [4:0] }), .sum({ \level_1_sums[15][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[227] [4:0] }), .sum({ \level_1_sums[15][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[15][113] [5:0] }),
     .b({ \level_1_sums[15][112] [5:0] }), .sum({ \level_2_sums[15][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[229] [4:0] }), .sum({ \level_1_sums[15][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[231] [4:0] }), .sum({ \level_1_sums[15][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[15][115] [5:0] }),
     .b({ \level_1_sums[15][114] [5:0] }), .sum({ \level_2_sums[15][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[15][57] [6:0] }), .b({ \level_2_sums[15][56] [6:0] }), .sum({ \level_3_sums[15][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[233] [4:0] }), .sum({ \level_1_sums[15][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[235] [4:0] }), .sum({ \level_1_sums[15][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[15][117] [5:0] }),
     .b({ \level_1_sums[15][116] [5:0] }), .sum({ \level_2_sums[15][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[237] [4:0] }), .sum({ \level_1_sums[15][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[239] [4:0] }), .sum({ \level_1_sums[15][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[15][119] [5:0] }),
     .b({ \level_1_sums[15][118] [5:0] }), .sum({ \level_2_sums[15][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[15][59] [6:0] }), .b({ \level_2_sums[15][58] [6:0] }), .sum({ \level_3_sums[15][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[15][29] [7:0] }),
     .b({ \level_3_sums[15][28] [7:0] }), .sum({ \level_4_sums[15][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[241] [4:0] }), .sum({ \level_1_sums[15][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[243] [4:0] }), .sum({ \level_1_sums[15][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[15][121] [5:0] }),
     .b({ \level_1_sums[15][120] [5:0] }), .sum({ \level_2_sums[15][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[245] [4:0] }), .sum({ \level_1_sums[15][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[247] [4:0] }), .sum({ \level_1_sums[15][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[15][123] [5:0] }),
     .b({ \level_1_sums[15][122] [5:0] }), .sum({ \level_2_sums[15][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[15][61] [6:0] }), .b({ \level_2_sums[15][60] [6:0] }), .sum({ \level_3_sums[15][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[249] [4:0] }), .sum({ \level_1_sums[15][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[251] [4:0] }), .sum({ \level_1_sums[15][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[15][125] [5:0] }),
     .b({ \level_1_sums[15][124] [5:0] }), .sum({ \level_2_sums[15][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[253] [4:0] }), .sum({ \level_1_sums[15][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[15].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[15].product_terms[255] [4:0] }), .sum({ \level_1_sums[15][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[15][127] [5:0] }),
     .b({ \level_1_sums[15][126] [5:0] }), .sum({ \level_2_sums[15][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[15][63] [6:0] }), .b({ \level_2_sums[15][62] [6:0] }), .sum({ \level_3_sums[15][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[15][31] [7:0] }),
     .b({ \level_3_sums[15][30] [7:0] }), .sum({ \level_4_sums[15][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[15][15] [8:0] }),
     .b({ \level_4_sums[15][14] [8:0] }), .sum({ \level_5_sums[15][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[15][7] [9:0] }),
     .b({ \level_5_sums[15][6] [9:0] }), .sum({ \level_6_sums[15][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[15][3] [9:0] }),
     .b({ \level_6_sums[15][2] [9:0] }), .sum({ \level_7_sums[15][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[15].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[15][0] [9:0] }),
     .b({ \level_7_sums[15][1] [9:0] }), .sum({ \level_8_sums[15] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[16].relu_inst (.in_data({ \final_sums[16] [9:0] }), .out_data({ \out_sig[16] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[1] [4:0] }), .sum({ \level_1_sums[16][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[3] [4:0] }), .sum({ \level_1_sums[16][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[16][1] [5:0] }),
     .b({ \level_1_sums[16][0] [5:0] }), .sum({ \level_2_sums[16][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[5] [4:0] }), .sum({ \level_1_sums[16][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[7] [4:0] }), .sum({ \level_1_sums[16][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[16][3] [5:0] }),
     .b({ \level_1_sums[16][2] [5:0] }), .sum({ \level_2_sums[16][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[16][1] [6:0] }),
     .b({ \level_2_sums[16][0] [6:0] }), .sum({ \level_3_sums[16][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[9] [4:0] }), .sum({ \level_1_sums[16][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[11] [4:0] }), .sum({ \level_1_sums[16][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[16][5] [5:0] }),
     .b({ \level_1_sums[16][4] [5:0] }), .sum({ \level_2_sums[16][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[13] [4:0] }), .sum({ \level_1_sums[16][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[15] [4:0] }), .sum({ \level_1_sums[16][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[16][7] [5:0] }),
     .b({ \level_1_sums[16][6] [5:0] }), .sum({ \level_2_sums[16][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[16][3] [6:0] }),
     .b({ \level_2_sums[16][2] [6:0] }), .sum({ \level_3_sums[16][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[16][1] [7:0] }),
     .b({ \level_3_sums[16][0] [7:0] }), .sum({ \level_4_sums[16][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[17] [4:0] }), .sum({ \level_1_sums[16][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[19] [4:0] }), .sum({ \level_1_sums[16][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[16][9] [5:0] }),
     .b({ \level_1_sums[16][8] [5:0] }), .sum({ \level_2_sums[16][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[21] [4:0] }), .sum({ \level_1_sums[16][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[23] [4:0] }), .sum({ \level_1_sums[16][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[16][11] [5:0] }),
     .b({ \level_1_sums[16][10] [5:0] }), .sum({ \level_2_sums[16][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[16][5] [6:0] }),
     .b({ \level_2_sums[16][4] [6:0] }), .sum({ \level_3_sums[16][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[25] [4:0] }), .sum({ \level_1_sums[16][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[27] [4:0] }), .sum({ \level_1_sums[16][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[16][13] [5:0] }),
     .b({ \level_1_sums[16][12] [5:0] }), .sum({ \level_2_sums[16][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[29] [4:0] }), .sum({ \level_1_sums[16][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[31] [4:0] }), .sum({ \level_1_sums[16][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[16][15] [5:0] }),
     .b({ \level_1_sums[16][14] [5:0] }), .sum({ \level_2_sums[16][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[16][7] [6:0] }),
     .b({ \level_2_sums[16][6] [6:0] }), .sum({ \level_3_sums[16][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[16][3] [7:0] }),
     .b({ \level_3_sums[16][2] [7:0] }), .sum({ \level_4_sums[16][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[16][1] [8:0] }),
     .b({ \level_4_sums[16][0] [8:0] }), .sum({ \level_5_sums[16][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[33] [4:0] }), .sum({ \level_1_sums[16][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[35] [4:0] }), .sum({ \level_1_sums[16][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[16][17] [5:0] }),
     .b({ \level_1_sums[16][16] [5:0] }), .sum({ \level_2_sums[16][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[37] [4:0] }), .sum({ \level_1_sums[16][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[39] [4:0] }), .sum({ \level_1_sums[16][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[16][19] [5:0] }),
     .b({ \level_1_sums[16][18] [5:0] }), .sum({ \level_2_sums[16][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[16][9] [6:0] }),
     .b({ \level_2_sums[16][8] [6:0] }), .sum({ \level_3_sums[16][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[41] [4:0] }), .sum({ \level_1_sums[16][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[43] [4:0] }), .sum({ \level_1_sums[16][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[16][21] [5:0] }),
     .b({ \level_1_sums[16][20] [5:0] }), .sum({ \level_2_sums[16][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[45] [4:0] }), .sum({ \level_1_sums[16][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[47] [4:0] }), .sum({ \level_1_sums[16][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[16][23] [5:0] }),
     .b({ \level_1_sums[16][22] [5:0] }), .sum({ \level_2_sums[16][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[16][11] [6:0] }),
     .b({ \level_2_sums[16][10] [6:0] }), .sum({ \level_3_sums[16][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[16][5] [7:0] }),
     .b({ \level_3_sums[16][4] [7:0] }), .sum({ \level_4_sums[16][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[49] [4:0] }), .sum({ \level_1_sums[16][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[51] [4:0] }), .sum({ \level_1_sums[16][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[16][25] [5:0] }),
     .b({ \level_1_sums[16][24] [5:0] }), .sum({ \level_2_sums[16][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[53] [4:0] }), .sum({ \level_1_sums[16][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[55] [4:0] }), .sum({ \level_1_sums[16][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[16][27] [5:0] }),
     .b({ \level_1_sums[16][26] [5:0] }), .sum({ \level_2_sums[16][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[16][13] [6:0] }),
     .b({ \level_2_sums[16][12] [6:0] }), .sum({ \level_3_sums[16][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[57] [4:0] }), .sum({ \level_1_sums[16][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[59] [4:0] }), .sum({ \level_1_sums[16][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[16][29] [5:0] }),
     .b({ \level_1_sums[16][28] [5:0] }), .sum({ \level_2_sums[16][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[61] [4:0] }), .sum({ \level_1_sums[16][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[63] [4:0] }), .sum({ \level_1_sums[16][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[16][31] [5:0] }),
     .b({ \level_1_sums[16][30] [5:0] }), .sum({ \level_2_sums[16][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[16][15] [6:0] }),
     .b({ \level_2_sums[16][14] [6:0] }), .sum({ \level_3_sums[16][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[16][7] [7:0] }),
     .b({ \level_3_sums[16][6] [7:0] }), .sum({ \level_4_sums[16][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[16][3] [8:0] }),
     .b({ \level_4_sums[16][2] [8:0] }), .sum({ \level_5_sums[16][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[16][1] [9:0] }),
     .b({ \level_5_sums[16][0] [9:0] }), .sum({ \level_6_sums[16][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[65] [4:0] }), .sum({ \level_1_sums[16][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[67] [4:0] }), .sum({ \level_1_sums[16][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[16][33] [5:0] }),
     .b({ \level_1_sums[16][32] [5:0] }), .sum({ \level_2_sums[16][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[69] [4:0] }), .sum({ \level_1_sums[16][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[71] [4:0] }), .sum({ \level_1_sums[16][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[16][35] [5:0] }),
     .b({ \level_1_sums[16][34] [5:0] }), .sum({ \level_2_sums[16][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[16][17] [6:0] }),
     .b({ \level_2_sums[16][16] [6:0] }), .sum({ \level_3_sums[16][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[73] [4:0] }), .sum({ \level_1_sums[16][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[75] [4:0] }), .sum({ \level_1_sums[16][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[16][37] [5:0] }),
     .b({ \level_1_sums[16][36] [5:0] }), .sum({ \level_2_sums[16][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[77] [4:0] }), .sum({ \level_1_sums[16][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[79] [4:0] }), .sum({ \level_1_sums[16][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[16][39] [5:0] }),
     .b({ \level_1_sums[16][38] [5:0] }), .sum({ \level_2_sums[16][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[16][19] [6:0] }),
     .b({ \level_2_sums[16][18] [6:0] }), .sum({ \level_3_sums[16][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[16][9] [7:0] }),
     .b({ \level_3_sums[16][8] [7:0] }), .sum({ \level_4_sums[16][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[81] [4:0] }), .sum({ \level_1_sums[16][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[83] [4:0] }), .sum({ \level_1_sums[16][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[16][41] [5:0] }),
     .b({ \level_1_sums[16][40] [5:0] }), .sum({ \level_2_sums[16][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[85] [4:0] }), .sum({ \level_1_sums[16][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[87] [4:0] }), .sum({ \level_1_sums[16][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[16][43] [5:0] }),
     .b({ \level_1_sums[16][42] [5:0] }), .sum({ \level_2_sums[16][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[16][21] [6:0] }),
     .b({ \level_2_sums[16][20] [6:0] }), .sum({ \level_3_sums[16][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[89] [4:0] }), .sum({ \level_1_sums[16][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[91] [4:0] }), .sum({ \level_1_sums[16][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[16][45] [5:0] }),
     .b({ \level_1_sums[16][44] [5:0] }), .sum({ \level_2_sums[16][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[93] [4:0] }), .sum({ \level_1_sums[16][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[95] [4:0] }), .sum({ \level_1_sums[16][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[16][47] [5:0] }),
     .b({ \level_1_sums[16][46] [5:0] }), .sum({ \level_2_sums[16][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[16][23] [6:0] }),
     .b({ \level_2_sums[16][22] [6:0] }), .sum({ \level_3_sums[16][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[16][11] [7:0] }),
     .b({ \level_3_sums[16][10] [7:0] }), .sum({ \level_4_sums[16][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[16][5] [8:0] }),
     .b({ \level_4_sums[16][4] [8:0] }), .sum({ \level_5_sums[16][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[97] [4:0] }), .sum({ \level_1_sums[16][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[99] [4:0] }), .sum({ \level_1_sums[16][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[16][49] [5:0] }),
     .b({ \level_1_sums[16][48] [5:0] }), .sum({ \level_2_sums[16][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[101] [4:0] }), .sum({ \level_1_sums[16][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[103] [4:0] }), .sum({ \level_1_sums[16][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[16][51] [5:0] }),
     .b({ \level_1_sums[16][50] [5:0] }), .sum({ \level_2_sums[16][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[16][25] [6:0] }), .b({ \level_2_sums[16][24] [6:0] }), .sum({ \level_3_sums[16][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[105] [4:0] }), .sum({ \level_1_sums[16][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[107] [4:0] }), .sum({ \level_1_sums[16][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[16][53] [5:0] }),
     .b({ \level_1_sums[16][52] [5:0] }), .sum({ \level_2_sums[16][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[109] [4:0] }), .sum({ \level_1_sums[16][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[111] [4:0] }), .sum({ \level_1_sums[16][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[16][55] [5:0] }),
     .b({ \level_1_sums[16][54] [5:0] }), .sum({ \level_2_sums[16][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[16][27] [6:0] }), .b({ \level_2_sums[16][26] [6:0] }), .sum({ \level_3_sums[16][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[16][13] [7:0] }),
     .b({ \level_3_sums[16][12] [7:0] }), .sum({ \level_4_sums[16][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[113] [4:0] }), .sum({ \level_1_sums[16][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[115] [4:0] }), .sum({ \level_1_sums[16][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[16][57] [5:0] }),
     .b({ \level_1_sums[16][56] [5:0] }), .sum({ \level_2_sums[16][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[117] [4:0] }), .sum({ \level_1_sums[16][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[119] [4:0] }), .sum({ \level_1_sums[16][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[16][59] [5:0] }),
     .b({ \level_1_sums[16][58] [5:0] }), .sum({ \level_2_sums[16][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[16][29] [6:0] }), .b({ \level_2_sums[16][28] [6:0] }), .sum({ \level_3_sums[16][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[121] [4:0] }), .sum({ \level_1_sums[16][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[123] [4:0] }), .sum({ \level_1_sums[16][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[16][61] [5:0] }),
     .b({ \level_1_sums[16][60] [5:0] }), .sum({ \level_2_sums[16][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[125] [4:0] }), .sum({ \level_1_sums[16][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[127] [4:0] }), .sum({ \level_1_sums[16][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[16][63] [5:0] }),
     .b({ \level_1_sums[16][62] [5:0] }), .sum({ \level_2_sums[16][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[16][31] [6:0] }), .b({ \level_2_sums[16][30] [6:0] }), .sum({ \level_3_sums[16][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[16][15] [7:0] }),
     .b({ \level_3_sums[16][14] [7:0] }), .sum({ \level_4_sums[16][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[16][7] [8:0] }),
     .b({ \level_4_sums[16][6] [8:0] }), .sum({ \level_5_sums[16][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[16][3] [9:0] }),
     .b({ \level_5_sums[16][2] [9:0] }), .sum({ \level_6_sums[16][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[16][1] [9:0] }),
     .b({ \level_6_sums[16][0] [9:0] }), .sum({ \level_7_sums[16][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[129] [4:0] }), .sum({ \level_1_sums[16][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[131] [4:0] }), .sum({ \level_1_sums[16][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[16][65] [5:0] }),
     .b({ \level_1_sums[16][64] [5:0] }), .sum({ \level_2_sums[16][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[133] [4:0] }), .sum({ \level_1_sums[16][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[135] [4:0] }), .sum({ \level_1_sums[16][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[16][67] [5:0] }),
     .b({ \level_1_sums[16][66] [5:0] }), .sum({ \level_2_sums[16][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[16][33] [6:0] }), .b({ \level_2_sums[16][32] [6:0] }), .sum({ \level_3_sums[16][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[137] [4:0] }), .sum({ \level_1_sums[16][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[139] [4:0] }), .sum({ \level_1_sums[16][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[16][69] [5:0] }),
     .b({ \level_1_sums[16][68] [5:0] }), .sum({ \level_2_sums[16][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[141] [4:0] }), .sum({ \level_1_sums[16][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[143] [4:0] }), .sum({ \level_1_sums[16][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[16][71] [5:0] }),
     .b({ \level_1_sums[16][70] [5:0] }), .sum({ \level_2_sums[16][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[16][35] [6:0] }), .b({ \level_2_sums[16][34] [6:0] }), .sum({ \level_3_sums[16][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[16][17] [7:0] }),
     .b({ \level_3_sums[16][16] [7:0] }), .sum({ \level_4_sums[16][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[145] [4:0] }), .sum({ \level_1_sums[16][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[147] [4:0] }), .sum({ \level_1_sums[16][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[16][73] [5:0] }),
     .b({ \level_1_sums[16][72] [5:0] }), .sum({ \level_2_sums[16][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[149] [4:0] }), .sum({ \level_1_sums[16][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[151] [4:0] }), .sum({ \level_1_sums[16][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[16][75] [5:0] }),
     .b({ \level_1_sums[16][74] [5:0] }), .sum({ \level_2_sums[16][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[16][37] [6:0] }), .b({ \level_2_sums[16][36] [6:0] }), .sum({ \level_3_sums[16][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[153] [4:0] }), .sum({ \level_1_sums[16][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[155] [4:0] }), .sum({ \level_1_sums[16][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[16][77] [5:0] }),
     .b({ \level_1_sums[16][76] [5:0] }), .sum({ \level_2_sums[16][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[157] [4:0] }), .sum({ \level_1_sums[16][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[159] [4:0] }), .sum({ \level_1_sums[16][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[16][79] [5:0] }),
     .b({ \level_1_sums[16][78] [5:0] }), .sum({ \level_2_sums[16][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[16][39] [6:0] }), .b({ \level_2_sums[16][38] [6:0] }), .sum({ \level_3_sums[16][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[16][19] [7:0] }),
     .b({ \level_3_sums[16][18] [7:0] }), .sum({ \level_4_sums[16][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[16][9] [8:0] }),
     .b({ \level_4_sums[16][8] [8:0] }), .sum({ \level_5_sums[16][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[161] [4:0] }), .sum({ \level_1_sums[16][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[163] [4:0] }), .sum({ \level_1_sums[16][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[16][81] [5:0] }),
     .b({ \level_1_sums[16][80] [5:0] }), .sum({ \level_2_sums[16][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[165] [4:0] }), .sum({ \level_1_sums[16][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[167] [4:0] }), .sum({ \level_1_sums[16][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[16][83] [5:0] }),
     .b({ \level_1_sums[16][82] [5:0] }), .sum({ \level_2_sums[16][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[16][41] [6:0] }), .b({ \level_2_sums[16][40] [6:0] }), .sum({ \level_3_sums[16][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[169] [4:0] }), .sum({ \level_1_sums[16][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[171] [4:0] }), .sum({ \level_1_sums[16][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[16][85] [5:0] }),
     .b({ \level_1_sums[16][84] [5:0] }), .sum({ \level_2_sums[16][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[173] [4:0] }), .sum({ \level_1_sums[16][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[175] [4:0] }), .sum({ \level_1_sums[16][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[16][87] [5:0] }),
     .b({ \level_1_sums[16][86] [5:0] }), .sum({ \level_2_sums[16][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[16][43] [6:0] }), .b({ \level_2_sums[16][42] [6:0] }), .sum({ \level_3_sums[16][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[16][21] [7:0] }),
     .b({ \level_3_sums[16][20] [7:0] }), .sum({ \level_4_sums[16][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[177] [4:0] }), .sum({ \level_1_sums[16][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[179] [4:0] }), .sum({ \level_1_sums[16][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[16][89] [5:0] }),
     .b({ \level_1_sums[16][88] [5:0] }), .sum({ \level_2_sums[16][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[181] [4:0] }), .sum({ \level_1_sums[16][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[183] [4:0] }), .sum({ \level_1_sums[16][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[16][91] [5:0] }),
     .b({ \level_1_sums[16][90] [5:0] }), .sum({ \level_2_sums[16][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[16][45] [6:0] }), .b({ \level_2_sums[16][44] [6:0] }), .sum({ \level_3_sums[16][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[185] [4:0] }), .sum({ \level_1_sums[16][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[187] [4:0] }), .sum({ \level_1_sums[16][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[16][93] [5:0] }),
     .b({ \level_1_sums[16][92] [5:0] }), .sum({ \level_2_sums[16][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[189] [4:0] }), .sum({ \level_1_sums[16][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[191] [4:0] }), .sum({ \level_1_sums[16][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[16][95] [5:0] }),
     .b({ \level_1_sums[16][94] [5:0] }), .sum({ \level_2_sums[16][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[16][47] [6:0] }), .b({ \level_2_sums[16][46] [6:0] }), .sum({ \level_3_sums[16][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[16][23] [7:0] }),
     .b({ \level_3_sums[16][22] [7:0] }), .sum({ \level_4_sums[16][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[16][11] [8:0] }),
     .b({ \level_4_sums[16][10] [8:0] }), .sum({ \level_5_sums[16][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[16][5] [9:0] }),
     .b({ \level_5_sums[16][4] [9:0] }), .sum({ \level_6_sums[16][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[193] [4:0] }), .sum({ \level_1_sums[16][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[195] [4:0] }), .sum({ \level_1_sums[16][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[16][97] [5:0] }),
     .b({ \level_1_sums[16][96] [5:0] }), .sum({ \level_2_sums[16][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[197] [4:0] }), .sum({ \level_1_sums[16][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[199] [4:0] }), .sum({ \level_1_sums[16][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[16][99] [5:0] }),
     .b({ \level_1_sums[16][98] [5:0] }), .sum({ \level_2_sums[16][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[16][49] [6:0] }), .b({ \level_2_sums[16][48] [6:0] }), .sum({ \level_3_sums[16][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[201] [4:0] }), .sum({ \level_1_sums[16][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[203] [4:0] }), .sum({ \level_1_sums[16][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[16][101] [5:0] }),
     .b({ \level_1_sums[16][100] [5:0] }), .sum({ \level_2_sums[16][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[205] [4:0] }), .sum({ \level_1_sums[16][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[207] [4:0] }), .sum({ \level_1_sums[16][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[16][103] [5:0] }),
     .b({ \level_1_sums[16][102] [5:0] }), .sum({ \level_2_sums[16][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[16][51] [6:0] }), .b({ \level_2_sums[16][50] [6:0] }), .sum({ \level_3_sums[16][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[16][25] [7:0] }),
     .b({ \level_3_sums[16][24] [7:0] }), .sum({ \level_4_sums[16][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[209] [4:0] }), .sum({ \level_1_sums[16][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[211] [4:0] }), .sum({ \level_1_sums[16][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[16][105] [5:0] }),
     .b({ \level_1_sums[16][104] [5:0] }), .sum({ \level_2_sums[16][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[213] [4:0] }), .sum({ \level_1_sums[16][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[215] [4:0] }), .sum({ \level_1_sums[16][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[16][107] [5:0] }),
     .b({ \level_1_sums[16][106] [5:0] }), .sum({ \level_2_sums[16][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[16][53] [6:0] }), .b({ \level_2_sums[16][52] [6:0] }), .sum({ \level_3_sums[16][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[217] [4:0] }), .sum({ \level_1_sums[16][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[219] [4:0] }), .sum({ \level_1_sums[16][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[16][109] [5:0] }),
     .b({ \level_1_sums[16][108] [5:0] }), .sum({ \level_2_sums[16][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[221] [4:0] }), .sum({ \level_1_sums[16][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[223] [4:0] }), .sum({ \level_1_sums[16][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[16][111] [5:0] }),
     .b({ \level_1_sums[16][110] [5:0] }), .sum({ \level_2_sums[16][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[16][55] [6:0] }), .b({ \level_2_sums[16][54] [6:0] }), .sum({ \level_3_sums[16][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[16][27] [7:0] }),
     .b({ \level_3_sums[16][26] [7:0] }), .sum({ \level_4_sums[16][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[16][13] [8:0] }),
     .b({ \level_4_sums[16][12] [8:0] }), .sum({ \level_5_sums[16][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[225] [4:0] }), .sum({ \level_1_sums[16][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[227] [4:0] }), .sum({ \level_1_sums[16][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[16][113] [5:0] }),
     .b({ \level_1_sums[16][112] [5:0] }), .sum({ \level_2_sums[16][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[229] [4:0] }), .sum({ \level_1_sums[16][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[231] [4:0] }), .sum({ \level_1_sums[16][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[16][115] [5:0] }),
     .b({ \level_1_sums[16][114] [5:0] }), .sum({ \level_2_sums[16][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[16][57] [6:0] }), .b({ \level_2_sums[16][56] [6:0] }), .sum({ \level_3_sums[16][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[233] [4:0] }), .sum({ \level_1_sums[16][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[235] [4:0] }), .sum({ \level_1_sums[16][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[16][117] [5:0] }),
     .b({ \level_1_sums[16][116] [5:0] }), .sum({ \level_2_sums[16][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[237] [4:0] }), .sum({ \level_1_sums[16][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[239] [4:0] }), .sum({ \level_1_sums[16][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[16][119] [5:0] }),
     .b({ \level_1_sums[16][118] [5:0] }), .sum({ \level_2_sums[16][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[16][59] [6:0] }), .b({ \level_2_sums[16][58] [6:0] }), .sum({ \level_3_sums[16][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[16][29] [7:0] }),
     .b({ \level_3_sums[16][28] [7:0] }), .sum({ \level_4_sums[16][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[241] [4:0] }), .sum({ \level_1_sums[16][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[243] [4:0] }), .sum({ \level_1_sums[16][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[16][121] [5:0] }),
     .b({ \level_1_sums[16][120] [5:0] }), .sum({ \level_2_sums[16][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[245] [4:0] }), .sum({ \level_1_sums[16][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[247] [4:0] }), .sum({ \level_1_sums[16][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[16][123] [5:0] }),
     .b({ \level_1_sums[16][122] [5:0] }), .sum({ \level_2_sums[16][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[16][61] [6:0] }), .b({ \level_2_sums[16][60] [6:0] }), .sum({ \level_3_sums[16][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[249] [4:0] }), .sum({ \level_1_sums[16][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[251] [4:0] }), .sum({ \level_1_sums[16][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[16][125] [5:0] }),
     .b({ \level_1_sums[16][124] [5:0] }), .sum({ \level_2_sums[16][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[253] [4:0] }), .sum({ \level_1_sums[16][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[16].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[16].product_terms[255] [4:0] }), .sum({ \level_1_sums[16][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[16][127] [5:0] }),
     .b({ \level_1_sums[16][126] [5:0] }), .sum({ \level_2_sums[16][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[16][63] [6:0] }), .b({ \level_2_sums[16][62] [6:0] }), .sum({ \level_3_sums[16][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[16][31] [7:0] }),
     .b({ \level_3_sums[16][30] [7:0] }), .sum({ \level_4_sums[16][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[16][15] [8:0] }),
     .b({ \level_4_sums[16][14] [8:0] }), .sum({ \level_5_sums[16][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[16][7] [9:0] }),
     .b({ \level_5_sums[16][6] [9:0] }), .sum({ \level_6_sums[16][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[16][3] [9:0] }),
     .b({ \level_6_sums[16][2] [9:0] }), .sum({ \level_7_sums[16][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[16].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[16][0] [9:0] }),
     .b({ \level_7_sums[16][1] [9:0] }), .sum({ \level_8_sums[16] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[17].relu_inst (.in_data({ \final_sums[17] [9:0] }), .out_data({ \out_sig[17] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[1] [4:0] }), .sum({ \level_1_sums[17][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[3] [4:0] }), .sum({ \level_1_sums[17][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[17][1] [5:0] }),
     .b({ \level_1_sums[17][0] [5:0] }), .sum({ \level_2_sums[17][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[5] [4:0] }), .sum({ \level_1_sums[17][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[7] [4:0] }), .sum({ \level_1_sums[17][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[17][3] [5:0] }),
     .b({ \level_1_sums[17][2] [5:0] }), .sum({ \level_2_sums[17][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[17][1] [6:0] }),
     .b({ \level_2_sums[17][0] [6:0] }), .sum({ \level_3_sums[17][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[9] [4:0] }), .sum({ \level_1_sums[17][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[11] [4:0] }), .sum({ \level_1_sums[17][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[17][5] [5:0] }),
     .b({ \level_1_sums[17][4] [5:0] }), .sum({ \level_2_sums[17][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[13] [4:0] }), .sum({ \level_1_sums[17][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[15] [4:0] }), .sum({ \level_1_sums[17][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[17][7] [5:0] }),
     .b({ \level_1_sums[17][6] [5:0] }), .sum({ \level_2_sums[17][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[17][3] [6:0] }),
     .b({ \level_2_sums[17][2] [6:0] }), .sum({ \level_3_sums[17][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[17][1] [7:0] }),
     .b({ \level_3_sums[17][0] [7:0] }), .sum({ \level_4_sums[17][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[17] [4:0] }), .sum({ \level_1_sums[17][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[19] [4:0] }), .sum({ \level_1_sums[17][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[17][9] [5:0] }),
     .b({ \level_1_sums[17][8] [5:0] }), .sum({ \level_2_sums[17][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[21] [4:0] }), .sum({ \level_1_sums[17][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[23] [4:0] }), .sum({ \level_1_sums[17][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[17][11] [5:0] }),
     .b({ \level_1_sums[17][10] [5:0] }), .sum({ \level_2_sums[17][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[17][5] [6:0] }),
     .b({ \level_2_sums[17][4] [6:0] }), .sum({ \level_3_sums[17][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[25] [4:0] }), .sum({ \level_1_sums[17][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[27] [4:0] }), .sum({ \level_1_sums[17][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[17][13] [5:0] }),
     .b({ \level_1_sums[17][12] [5:0] }), .sum({ \level_2_sums[17][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[29] [4:0] }), .sum({ \level_1_sums[17][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[31] [4:0] }), .sum({ \level_1_sums[17][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[17][15] [5:0] }),
     .b({ \level_1_sums[17][14] [5:0] }), .sum({ \level_2_sums[17][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[17][7] [6:0] }),
     .b({ \level_2_sums[17][6] [6:0] }), .sum({ \level_3_sums[17][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[17][3] [7:0] }),
     .b({ \level_3_sums[17][2] [7:0] }), .sum({ \level_4_sums[17][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[17][1] [8:0] }),
     .b({ \level_4_sums[17][0] [8:0] }), .sum({ \level_5_sums[17][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[33] [4:0] }), .sum({ \level_1_sums[17][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[35] [4:0] }), .sum({ \level_1_sums[17][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[17][17] [5:0] }),
     .b({ \level_1_sums[17][16] [5:0] }), .sum({ \level_2_sums[17][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[37] [4:0] }), .sum({ \level_1_sums[17][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[39] [4:0] }), .sum({ \level_1_sums[17][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[17][19] [5:0] }),
     .b({ \level_1_sums[17][18] [5:0] }), .sum({ \level_2_sums[17][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[17][9] [6:0] }),
     .b({ \level_2_sums[17][8] [6:0] }), .sum({ \level_3_sums[17][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[41] [4:0] }), .sum({ \level_1_sums[17][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[43] [4:0] }), .sum({ \level_1_sums[17][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[17][21] [5:0] }),
     .b({ \level_1_sums[17][20] [5:0] }), .sum({ \level_2_sums[17][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[45] [4:0] }), .sum({ \level_1_sums[17][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[47] [4:0] }), .sum({ \level_1_sums[17][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[17][23] [5:0] }),
     .b({ \level_1_sums[17][22] [5:0] }), .sum({ \level_2_sums[17][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[17][11] [6:0] }),
     .b({ \level_2_sums[17][10] [6:0] }), .sum({ \level_3_sums[17][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[17][5] [7:0] }),
     .b({ \level_3_sums[17][4] [7:0] }), .sum({ \level_4_sums[17][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[49] [4:0] }), .sum({ \level_1_sums[17][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[51] [4:0] }), .sum({ \level_1_sums[17][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[17][25] [5:0] }),
     .b({ \level_1_sums[17][24] [5:0] }), .sum({ \level_2_sums[17][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[53] [4:0] }), .sum({ \level_1_sums[17][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[55] [4:0] }), .sum({ \level_1_sums[17][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[17][27] [5:0] }),
     .b({ \level_1_sums[17][26] [5:0] }), .sum({ \level_2_sums[17][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[17][13] [6:0] }),
     .b({ \level_2_sums[17][12] [6:0] }), .sum({ \level_3_sums[17][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[57] [4:0] }), .sum({ \level_1_sums[17][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[59] [4:0] }), .sum({ \level_1_sums[17][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[17][29] [5:0] }),
     .b({ \level_1_sums[17][28] [5:0] }), .sum({ \level_2_sums[17][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[61] [4:0] }), .sum({ \level_1_sums[17][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[63] [4:0] }), .sum({ \level_1_sums[17][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[17][31] [5:0] }),
     .b({ \level_1_sums[17][30] [5:0] }), .sum({ \level_2_sums[17][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[17][15] [6:0] }),
     .b({ \level_2_sums[17][14] [6:0] }), .sum({ \level_3_sums[17][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[17][7] [7:0] }),
     .b({ \level_3_sums[17][6] [7:0] }), .sum({ \level_4_sums[17][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[17][3] [8:0] }),
     .b({ \level_4_sums[17][2] [8:0] }), .sum({ \level_5_sums[17][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[17][1] [9:0] }),
     .b({ \level_5_sums[17][0] [9:0] }), .sum({ \level_6_sums[17][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[65] [4:0] }), .sum({ \level_1_sums[17][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[67] [4:0] }), .sum({ \level_1_sums[17][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[17][33] [5:0] }),
     .b({ \level_1_sums[17][32] [5:0] }), .sum({ \level_2_sums[17][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[69] [4:0] }), .sum({ \level_1_sums[17][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[71] [4:0] }), .sum({ \level_1_sums[17][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[17][35] [5:0] }),
     .b({ \level_1_sums[17][34] [5:0] }), .sum({ \level_2_sums[17][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[17][17] [6:0] }),
     .b({ \level_2_sums[17][16] [6:0] }), .sum({ \level_3_sums[17][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[73] [4:0] }), .sum({ \level_1_sums[17][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[75] [4:0] }), .sum({ \level_1_sums[17][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[17][37] [5:0] }),
     .b({ \level_1_sums[17][36] [5:0] }), .sum({ \level_2_sums[17][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[77] [4:0] }), .sum({ \level_1_sums[17][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[79] [4:0] }), .sum({ \level_1_sums[17][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[17][39] [5:0] }),
     .b({ \level_1_sums[17][38] [5:0] }), .sum({ \level_2_sums[17][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[17][19] [6:0] }),
     .b({ \level_2_sums[17][18] [6:0] }), .sum({ \level_3_sums[17][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[17][9] [7:0] }),
     .b({ \level_3_sums[17][8] [7:0] }), .sum({ \level_4_sums[17][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[81] [4:0] }), .sum({ \level_1_sums[17][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[83] [4:0] }), .sum({ \level_1_sums[17][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[17][41] [5:0] }),
     .b({ \level_1_sums[17][40] [5:0] }), .sum({ \level_2_sums[17][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[85] [4:0] }), .sum({ \level_1_sums[17][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[87] [4:0] }), .sum({ \level_1_sums[17][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[17][43] [5:0] }),
     .b({ \level_1_sums[17][42] [5:0] }), .sum({ \level_2_sums[17][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[17][21] [6:0] }),
     .b({ \level_2_sums[17][20] [6:0] }), .sum({ \level_3_sums[17][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[89] [4:0] }), .sum({ \level_1_sums[17][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[91] [4:0] }), .sum({ \level_1_sums[17][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[17][45] [5:0] }),
     .b({ \level_1_sums[17][44] [5:0] }), .sum({ \level_2_sums[17][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[93] [4:0] }), .sum({ \level_1_sums[17][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[95] [4:0] }), .sum({ \level_1_sums[17][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[17][47] [5:0] }),
     .b({ \level_1_sums[17][46] [5:0] }), .sum({ \level_2_sums[17][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[17][23] [6:0] }),
     .b({ \level_2_sums[17][22] [6:0] }), .sum({ \level_3_sums[17][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[17][11] [7:0] }),
     .b({ \level_3_sums[17][10] [7:0] }), .sum({ \level_4_sums[17][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[17][5] [8:0] }),
     .b({ \level_4_sums[17][4] [8:0] }), .sum({ \level_5_sums[17][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[97] [4:0] }), .sum({ \level_1_sums[17][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[99] [4:0] }), .sum({ \level_1_sums[17][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[17][49] [5:0] }),
     .b({ \level_1_sums[17][48] [5:0] }), .sum({ \level_2_sums[17][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[101] [4:0] }), .sum({ \level_1_sums[17][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[103] [4:0] }), .sum({ \level_1_sums[17][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[17][51] [5:0] }),
     .b({ \level_1_sums[17][50] [5:0] }), .sum({ \level_2_sums[17][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[17][25] [6:0] }), .b({ \level_2_sums[17][24] [6:0] }), .sum({ \level_3_sums[17][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[105] [4:0] }), .sum({ \level_1_sums[17][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[107] [4:0] }), .sum({ \level_1_sums[17][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[17][53] [5:0] }),
     .b({ \level_1_sums[17][52] [5:0] }), .sum({ \level_2_sums[17][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[109] [4:0] }), .sum({ \level_1_sums[17][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[111] [4:0] }), .sum({ \level_1_sums[17][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[17][55] [5:0] }),
     .b({ \level_1_sums[17][54] [5:0] }), .sum({ \level_2_sums[17][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[17][27] [6:0] }), .b({ \level_2_sums[17][26] [6:0] }), .sum({ \level_3_sums[17][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[17][13] [7:0] }),
     .b({ \level_3_sums[17][12] [7:0] }), .sum({ \level_4_sums[17][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[113] [4:0] }), .sum({ \level_1_sums[17][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[115] [4:0] }), .sum({ \level_1_sums[17][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[17][57] [5:0] }),
     .b({ \level_1_sums[17][56] [5:0] }), .sum({ \level_2_sums[17][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[117] [4:0] }), .sum({ \level_1_sums[17][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[119] [4:0] }), .sum({ \level_1_sums[17][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[17][59] [5:0] }),
     .b({ \level_1_sums[17][58] [5:0] }), .sum({ \level_2_sums[17][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[17][29] [6:0] }), .b({ \level_2_sums[17][28] [6:0] }), .sum({ \level_3_sums[17][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[121] [4:0] }), .sum({ \level_1_sums[17][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[123] [4:0] }), .sum({ \level_1_sums[17][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[17][61] [5:0] }),
     .b({ \level_1_sums[17][60] [5:0] }), .sum({ \level_2_sums[17][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[125] [4:0] }), .sum({ \level_1_sums[17][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[127] [4:0] }), .sum({ \level_1_sums[17][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[17][63] [5:0] }),
     .b({ \level_1_sums[17][62] [5:0] }), .sum({ \level_2_sums[17][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[17][31] [6:0] }), .b({ \level_2_sums[17][30] [6:0] }), .sum({ \level_3_sums[17][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[17][15] [7:0] }),
     .b({ \level_3_sums[17][14] [7:0] }), .sum({ \level_4_sums[17][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[17][7] [8:0] }),
     .b({ \level_4_sums[17][6] [8:0] }), .sum({ \level_5_sums[17][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[17][3] [9:0] }),
     .b({ \level_5_sums[17][2] [9:0] }), .sum({ \level_6_sums[17][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[17][1] [9:0] }),
     .b({ \level_6_sums[17][0] [9:0] }), .sum({ \level_7_sums[17][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[129] [4:0] }), .sum({ \level_1_sums[17][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[131] [4:0] }), .sum({ \level_1_sums[17][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[17][65] [5:0] }),
     .b({ \level_1_sums[17][64] [5:0] }), .sum({ \level_2_sums[17][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[133] [4:0] }), .sum({ \level_1_sums[17][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[135] [4:0] }), .sum({ \level_1_sums[17][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[17][67] [5:0] }),
     .b({ \level_1_sums[17][66] [5:0] }), .sum({ \level_2_sums[17][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[17][33] [6:0] }), .b({ \level_2_sums[17][32] [6:0] }), .sum({ \level_3_sums[17][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[137] [4:0] }), .sum({ \level_1_sums[17][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[139] [4:0] }), .sum({ \level_1_sums[17][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[17][69] [5:0] }),
     .b({ \level_1_sums[17][68] [5:0] }), .sum({ \level_2_sums[17][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[141] [4:0] }), .sum({ \level_1_sums[17][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[143] [4:0] }), .sum({ \level_1_sums[17][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[17][71] [5:0] }),
     .b({ \level_1_sums[17][70] [5:0] }), .sum({ \level_2_sums[17][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[17][35] [6:0] }), .b({ \level_2_sums[17][34] [6:0] }), .sum({ \level_3_sums[17][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[17][17] [7:0] }),
     .b({ \level_3_sums[17][16] [7:0] }), .sum({ \level_4_sums[17][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[145] [4:0] }), .sum({ \level_1_sums[17][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[147] [4:0] }), .sum({ \level_1_sums[17][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[17][73] [5:0] }),
     .b({ \level_1_sums[17][72] [5:0] }), .sum({ \level_2_sums[17][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[149] [4:0] }), .sum({ \level_1_sums[17][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[151] [4:0] }), .sum({ \level_1_sums[17][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[17][75] [5:0] }),
     .b({ \level_1_sums[17][74] [5:0] }), .sum({ \level_2_sums[17][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[17][37] [6:0] }), .b({ \level_2_sums[17][36] [6:0] }), .sum({ \level_3_sums[17][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[153] [4:0] }), .sum({ \level_1_sums[17][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[155] [4:0] }), .sum({ \level_1_sums[17][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[17][77] [5:0] }),
     .b({ \level_1_sums[17][76] [5:0] }), .sum({ \level_2_sums[17][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[157] [4:0] }), .sum({ \level_1_sums[17][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[159] [4:0] }), .sum({ \level_1_sums[17][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[17][79] [5:0] }),
     .b({ \level_1_sums[17][78] [5:0] }), .sum({ \level_2_sums[17][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[17][39] [6:0] }), .b({ \level_2_sums[17][38] [6:0] }), .sum({ \level_3_sums[17][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[17][19] [7:0] }),
     .b({ \level_3_sums[17][18] [7:0] }), .sum({ \level_4_sums[17][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[17][9] [8:0] }),
     .b({ \level_4_sums[17][8] [8:0] }), .sum({ \level_5_sums[17][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[161] [4:0] }), .sum({ \level_1_sums[17][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[163] [4:0] }), .sum({ \level_1_sums[17][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[17][81] [5:0] }),
     .b({ \level_1_sums[17][80] [5:0] }), .sum({ \level_2_sums[17][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[165] [4:0] }), .sum({ \level_1_sums[17][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[167] [4:0] }), .sum({ \level_1_sums[17][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[17][83] [5:0] }),
     .b({ \level_1_sums[17][82] [5:0] }), .sum({ \level_2_sums[17][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[17][41] [6:0] }), .b({ \level_2_sums[17][40] [6:0] }), .sum({ \level_3_sums[17][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[169] [4:0] }), .sum({ \level_1_sums[17][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[171] [4:0] }), .sum({ \level_1_sums[17][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[17][85] [5:0] }),
     .b({ \level_1_sums[17][84] [5:0] }), .sum({ \level_2_sums[17][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[173] [4:0] }), .sum({ \level_1_sums[17][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[175] [4:0] }), .sum({ \level_1_sums[17][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[17][87] [5:0] }),
     .b({ \level_1_sums[17][86] [5:0] }), .sum({ \level_2_sums[17][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[17][43] [6:0] }), .b({ \level_2_sums[17][42] [6:0] }), .sum({ \level_3_sums[17][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[17][21] [7:0] }),
     .b({ \level_3_sums[17][20] [7:0] }), .sum({ \level_4_sums[17][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[177] [4:0] }), .sum({ \level_1_sums[17][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[179] [4:0] }), .sum({ \level_1_sums[17][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[17][89] [5:0] }),
     .b({ \level_1_sums[17][88] [5:0] }), .sum({ \level_2_sums[17][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[181] [4:0] }), .sum({ \level_1_sums[17][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[183] [4:0] }), .sum({ \level_1_sums[17][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[17][91] [5:0] }),
     .b({ \level_1_sums[17][90] [5:0] }), .sum({ \level_2_sums[17][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[17][45] [6:0] }), .b({ \level_2_sums[17][44] [6:0] }), .sum({ \level_3_sums[17][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[185] [4:0] }), .sum({ \level_1_sums[17][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[187] [4:0] }), .sum({ \level_1_sums[17][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[17][93] [5:0] }),
     .b({ \level_1_sums[17][92] [5:0] }), .sum({ \level_2_sums[17][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[189] [4:0] }), .sum({ \level_1_sums[17][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[191] [4:0] }), .sum({ \level_1_sums[17][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[17][95] [5:0] }),
     .b({ \level_1_sums[17][94] [5:0] }), .sum({ \level_2_sums[17][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[17][47] [6:0] }), .b({ \level_2_sums[17][46] [6:0] }), .sum({ \level_3_sums[17][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[17][23] [7:0] }),
     .b({ \level_3_sums[17][22] [7:0] }), .sum({ \level_4_sums[17][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[17][11] [8:0] }),
     .b({ \level_4_sums[17][10] [8:0] }), .sum({ \level_5_sums[17][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[17][5] [9:0] }),
     .b({ \level_5_sums[17][4] [9:0] }), .sum({ \level_6_sums[17][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[193] [4:0] }), .sum({ \level_1_sums[17][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[195] [4:0] }), .sum({ \level_1_sums[17][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[17][97] [5:0] }),
     .b({ \level_1_sums[17][96] [5:0] }), .sum({ \level_2_sums[17][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[197] [4:0] }), .sum({ \level_1_sums[17][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[199] [4:0] }), .sum({ \level_1_sums[17][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[17][99] [5:0] }),
     .b({ \level_1_sums[17][98] [5:0] }), .sum({ \level_2_sums[17][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[17][49] [6:0] }), .b({ \level_2_sums[17][48] [6:0] }), .sum({ \level_3_sums[17][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[201] [4:0] }), .sum({ \level_1_sums[17][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[203] [4:0] }), .sum({ \level_1_sums[17][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[17][101] [5:0] }),
     .b({ \level_1_sums[17][100] [5:0] }), .sum({ \level_2_sums[17][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[205] [4:0] }), .sum({ \level_1_sums[17][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[207] [4:0] }), .sum({ \level_1_sums[17][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[17][103] [5:0] }),
     .b({ \level_1_sums[17][102] [5:0] }), .sum({ \level_2_sums[17][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[17][51] [6:0] }), .b({ \level_2_sums[17][50] [6:0] }), .sum({ \level_3_sums[17][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[17][25] [7:0] }),
     .b({ \level_3_sums[17][24] [7:0] }), .sum({ \level_4_sums[17][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[209] [4:0] }), .sum({ \level_1_sums[17][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[211] [4:0] }), .sum({ \level_1_sums[17][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[17][105] [5:0] }),
     .b({ \level_1_sums[17][104] [5:0] }), .sum({ \level_2_sums[17][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[213] [4:0] }), .sum({ \level_1_sums[17][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[215] [4:0] }), .sum({ \level_1_sums[17][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[17][107] [5:0] }),
     .b({ \level_1_sums[17][106] [5:0] }), .sum({ \level_2_sums[17][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[17][53] [6:0] }), .b({ \level_2_sums[17][52] [6:0] }), .sum({ \level_3_sums[17][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[217] [4:0] }), .sum({ \level_1_sums[17][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[219] [4:0] }), .sum({ \level_1_sums[17][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[17][109] [5:0] }),
     .b({ \level_1_sums[17][108] [5:0] }), .sum({ \level_2_sums[17][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[221] [4:0] }), .sum({ \level_1_sums[17][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[223] [4:0] }), .sum({ \level_1_sums[17][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[17][111] [5:0] }),
     .b({ \level_1_sums[17][110] [5:0] }), .sum({ \level_2_sums[17][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[17][55] [6:0] }), .b({ \level_2_sums[17][54] [6:0] }), .sum({ \level_3_sums[17][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[17][27] [7:0] }),
     .b({ \level_3_sums[17][26] [7:0] }), .sum({ \level_4_sums[17][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[17][13] [8:0] }),
     .b({ \level_4_sums[17][12] [8:0] }), .sum({ \level_5_sums[17][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[225] [4:0] }), .sum({ \level_1_sums[17][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[227] [4:0] }), .sum({ \level_1_sums[17][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[17][113] [5:0] }),
     .b({ \level_1_sums[17][112] [5:0] }), .sum({ \level_2_sums[17][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[229] [4:0] }), .sum({ \level_1_sums[17][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[231] [4:0] }), .sum({ \level_1_sums[17][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[17][115] [5:0] }),
     .b({ \level_1_sums[17][114] [5:0] }), .sum({ \level_2_sums[17][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[17][57] [6:0] }), .b({ \level_2_sums[17][56] [6:0] }), .sum({ \level_3_sums[17][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[233] [4:0] }), .sum({ \level_1_sums[17][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[235] [4:0] }), .sum({ \level_1_sums[17][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[17][117] [5:0] }),
     .b({ \level_1_sums[17][116] [5:0] }), .sum({ \level_2_sums[17][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[237] [4:0] }), .sum({ \level_1_sums[17][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[239] [4:0] }), .sum({ \level_1_sums[17][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[17][119] [5:0] }),
     .b({ \level_1_sums[17][118] [5:0] }), .sum({ \level_2_sums[17][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[17][59] [6:0] }), .b({ \level_2_sums[17][58] [6:0] }), .sum({ \level_3_sums[17][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[17][29] [7:0] }),
     .b({ \level_3_sums[17][28] [7:0] }), .sum({ \level_4_sums[17][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[241] [4:0] }), .sum({ \level_1_sums[17][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[243] [4:0] }), .sum({ \level_1_sums[17][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[17][121] [5:0] }),
     .b({ \level_1_sums[17][120] [5:0] }), .sum({ \level_2_sums[17][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[245] [4:0] }), .sum({ \level_1_sums[17][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[247] [4:0] }), .sum({ \level_1_sums[17][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[17][123] [5:0] }),
     .b({ \level_1_sums[17][122] [5:0] }), .sum({ \level_2_sums[17][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[17][61] [6:0] }), .b({ \level_2_sums[17][60] [6:0] }), .sum({ \level_3_sums[17][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[249] [4:0] }), .sum({ \level_1_sums[17][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[251] [4:0] }), .sum({ \level_1_sums[17][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[17][125] [5:0] }),
     .b({ \level_1_sums[17][124] [5:0] }), .sum({ \level_2_sums[17][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[253] [4:0] }), .sum({ \level_1_sums[17][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[17].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[17].product_terms[255] [4:0] }), .sum({ \level_1_sums[17][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[17][127] [5:0] }),
     .b({ \level_1_sums[17][126] [5:0] }), .sum({ \level_2_sums[17][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[17][63] [6:0] }), .b({ \level_2_sums[17][62] [6:0] }), .sum({ \level_3_sums[17][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[17][31] [7:0] }),
     .b({ \level_3_sums[17][30] [7:0] }), .sum({ \level_4_sums[17][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[17][15] [8:0] }),
     .b({ \level_4_sums[17][14] [8:0] }), .sum({ \level_5_sums[17][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[17][7] [9:0] }),
     .b({ \level_5_sums[17][6] [9:0] }), .sum({ \level_6_sums[17][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[17][3] [9:0] }),
     .b({ \level_6_sums[17][2] [9:0] }), .sum({ \level_7_sums[17][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[17].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[17][0] [9:0] }),
     .b({ \level_7_sums[17][1] [9:0] }), .sum({ \level_8_sums[17] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[18].relu_inst (.in_data({ \final_sums[18] [9:0] }), .out_data({ \out_sig[18] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[1] [4:0] }), .sum({ \level_1_sums[18][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[3] [4:0] }), .sum({ \level_1_sums[18][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[18][1] [5:0] }),
     .b({ \level_1_sums[18][0] [5:0] }), .sum({ \level_2_sums[18][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[5] [4:0] }), .sum({ \level_1_sums[18][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[7] [4:0] }), .sum({ \level_1_sums[18][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[18][3] [5:0] }),
     .b({ \level_1_sums[18][2] [5:0] }), .sum({ \level_2_sums[18][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[18][1] [6:0] }),
     .b({ \level_2_sums[18][0] [6:0] }), .sum({ \level_3_sums[18][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[9] [4:0] }), .sum({ \level_1_sums[18][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[11] [4:0] }), .sum({ \level_1_sums[18][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[18][5] [5:0] }),
     .b({ \level_1_sums[18][4] [5:0] }), .sum({ \level_2_sums[18][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[13] [4:0] }), .sum({ \level_1_sums[18][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[15] [4:0] }), .sum({ \level_1_sums[18][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[18][7] [5:0] }),
     .b({ \level_1_sums[18][6] [5:0] }), .sum({ \level_2_sums[18][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[18][3] [6:0] }),
     .b({ \level_2_sums[18][2] [6:0] }), .sum({ \level_3_sums[18][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[18][1] [7:0] }),
     .b({ \level_3_sums[18][0] [7:0] }), .sum({ \level_4_sums[18][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[17] [4:0] }), .sum({ \level_1_sums[18][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[19] [4:0] }), .sum({ \level_1_sums[18][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[18][9] [5:0] }),
     .b({ \level_1_sums[18][8] [5:0] }), .sum({ \level_2_sums[18][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[21] [4:0] }), .sum({ \level_1_sums[18][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[23] [4:0] }), .sum({ \level_1_sums[18][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[18][11] [5:0] }),
     .b({ \level_1_sums[18][10] [5:0] }), .sum({ \level_2_sums[18][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[18][5] [6:0] }),
     .b({ \level_2_sums[18][4] [6:0] }), .sum({ \level_3_sums[18][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[25] [4:0] }), .sum({ \level_1_sums[18][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[27] [4:0] }), .sum({ \level_1_sums[18][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[18][13] [5:0] }),
     .b({ \level_1_sums[18][12] [5:0] }), .sum({ \level_2_sums[18][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[29] [4:0] }), .sum({ \level_1_sums[18][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[31] [4:0] }), .sum({ \level_1_sums[18][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[18][15] [5:0] }),
     .b({ \level_1_sums[18][14] [5:0] }), .sum({ \level_2_sums[18][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[18][7] [6:0] }),
     .b({ \level_2_sums[18][6] [6:0] }), .sum({ \level_3_sums[18][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[18][3] [7:0] }),
     .b({ \level_3_sums[18][2] [7:0] }), .sum({ \level_4_sums[18][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[18][1] [8:0] }),
     .b({ \level_4_sums[18][0] [8:0] }), .sum({ \level_5_sums[18][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[33] [4:0] }), .sum({ \level_1_sums[18][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[35] [4:0] }), .sum({ \level_1_sums[18][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[18][17] [5:0] }),
     .b({ \level_1_sums[18][16] [5:0] }), .sum({ \level_2_sums[18][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[37] [4:0] }), .sum({ \level_1_sums[18][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[39] [4:0] }), .sum({ \level_1_sums[18][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[18][19] [5:0] }),
     .b({ \level_1_sums[18][18] [5:0] }), .sum({ \level_2_sums[18][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[18][9] [6:0] }),
     .b({ \level_2_sums[18][8] [6:0] }), .sum({ \level_3_sums[18][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[41] [4:0] }), .sum({ \level_1_sums[18][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[43] [4:0] }), .sum({ \level_1_sums[18][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[18][21] [5:0] }),
     .b({ \level_1_sums[18][20] [5:0] }), .sum({ \level_2_sums[18][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[45] [4:0] }), .sum({ \level_1_sums[18][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[47] [4:0] }), .sum({ \level_1_sums[18][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[18][23] [5:0] }),
     .b({ \level_1_sums[18][22] [5:0] }), .sum({ \level_2_sums[18][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[18][11] [6:0] }),
     .b({ \level_2_sums[18][10] [6:0] }), .sum({ \level_3_sums[18][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[18][5] [7:0] }),
     .b({ \level_3_sums[18][4] [7:0] }), .sum({ \level_4_sums[18][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[49] [4:0] }), .sum({ \level_1_sums[18][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[51] [4:0] }), .sum({ \level_1_sums[18][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[18][25] [5:0] }),
     .b({ \level_1_sums[18][24] [5:0] }), .sum({ \level_2_sums[18][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[53] [4:0] }), .sum({ \level_1_sums[18][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[55] [4:0] }), .sum({ \level_1_sums[18][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[18][27] [5:0] }),
     .b({ \level_1_sums[18][26] [5:0] }), .sum({ \level_2_sums[18][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[18][13] [6:0] }),
     .b({ \level_2_sums[18][12] [6:0] }), .sum({ \level_3_sums[18][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[57] [4:0] }), .sum({ \level_1_sums[18][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[59] [4:0] }), .sum({ \level_1_sums[18][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[18][29] [5:0] }),
     .b({ \level_1_sums[18][28] [5:0] }), .sum({ \level_2_sums[18][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[61] [4:0] }), .sum({ \level_1_sums[18][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[63] [4:0] }), .sum({ \level_1_sums[18][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[18][31] [5:0] }),
     .b({ \level_1_sums[18][30] [5:0] }), .sum({ \level_2_sums[18][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[18][15] [6:0] }),
     .b({ \level_2_sums[18][14] [6:0] }), .sum({ \level_3_sums[18][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[18][7] [7:0] }),
     .b({ \level_3_sums[18][6] [7:0] }), .sum({ \level_4_sums[18][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[18][3] [8:0] }),
     .b({ \level_4_sums[18][2] [8:0] }), .sum({ \level_5_sums[18][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[18][1] [9:0] }),
     .b({ \level_5_sums[18][0] [9:0] }), .sum({ \level_6_sums[18][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[65] [4:0] }), .sum({ \level_1_sums[18][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[67] [4:0] }), .sum({ \level_1_sums[18][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[18][33] [5:0] }),
     .b({ \level_1_sums[18][32] [5:0] }), .sum({ \level_2_sums[18][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[69] [4:0] }), .sum({ \level_1_sums[18][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[71] [4:0] }), .sum({ \level_1_sums[18][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[18][35] [5:0] }),
     .b({ \level_1_sums[18][34] [5:0] }), .sum({ \level_2_sums[18][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[18][17] [6:0] }),
     .b({ \level_2_sums[18][16] [6:0] }), .sum({ \level_3_sums[18][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[73] [4:0] }), .sum({ \level_1_sums[18][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[75] [4:0] }), .sum({ \level_1_sums[18][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[18][37] [5:0] }),
     .b({ \level_1_sums[18][36] [5:0] }), .sum({ \level_2_sums[18][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[77] [4:0] }), .sum({ \level_1_sums[18][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[79] [4:0] }), .sum({ \level_1_sums[18][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[18][39] [5:0] }),
     .b({ \level_1_sums[18][38] [5:0] }), .sum({ \level_2_sums[18][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[18][19] [6:0] }),
     .b({ \level_2_sums[18][18] [6:0] }), .sum({ \level_3_sums[18][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[18][9] [7:0] }),
     .b({ \level_3_sums[18][8] [7:0] }), .sum({ \level_4_sums[18][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[81] [4:0] }), .sum({ \level_1_sums[18][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[83] [4:0] }), .sum({ \level_1_sums[18][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[18][41] [5:0] }),
     .b({ \level_1_sums[18][40] [5:0] }), .sum({ \level_2_sums[18][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[85] [4:0] }), .sum({ \level_1_sums[18][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[87] [4:0] }), .sum({ \level_1_sums[18][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[18][43] [5:0] }),
     .b({ \level_1_sums[18][42] [5:0] }), .sum({ \level_2_sums[18][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[18][21] [6:0] }),
     .b({ \level_2_sums[18][20] [6:0] }), .sum({ \level_3_sums[18][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[89] [4:0] }), .sum({ \level_1_sums[18][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[91] [4:0] }), .sum({ \level_1_sums[18][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[18][45] [5:0] }),
     .b({ \level_1_sums[18][44] [5:0] }), .sum({ \level_2_sums[18][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[93] [4:0] }), .sum({ \level_1_sums[18][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[95] [4:0] }), .sum({ \level_1_sums[18][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[18][47] [5:0] }),
     .b({ \level_1_sums[18][46] [5:0] }), .sum({ \level_2_sums[18][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[18][23] [6:0] }),
     .b({ \level_2_sums[18][22] [6:0] }), .sum({ \level_3_sums[18][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[18][11] [7:0] }),
     .b({ \level_3_sums[18][10] [7:0] }), .sum({ \level_4_sums[18][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[18][5] [8:0] }),
     .b({ \level_4_sums[18][4] [8:0] }), .sum({ \level_5_sums[18][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[97] [4:0] }), .sum({ \level_1_sums[18][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[99] [4:0] }), .sum({ \level_1_sums[18][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[18][49] [5:0] }),
     .b({ \level_1_sums[18][48] [5:0] }), .sum({ \level_2_sums[18][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[101] [4:0] }), .sum({ \level_1_sums[18][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[103] [4:0] }), .sum({ \level_1_sums[18][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[18][51] [5:0] }),
     .b({ \level_1_sums[18][50] [5:0] }), .sum({ \level_2_sums[18][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[18][25] [6:0] }), .b({ \level_2_sums[18][24] [6:0] }), .sum({ \level_3_sums[18][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[105] [4:0] }), .sum({ \level_1_sums[18][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[107] [4:0] }), .sum({ \level_1_sums[18][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[18][53] [5:0] }),
     .b({ \level_1_sums[18][52] [5:0] }), .sum({ \level_2_sums[18][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[109] [4:0] }), .sum({ \level_1_sums[18][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[111] [4:0] }), .sum({ \level_1_sums[18][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[18][55] [5:0] }),
     .b({ \level_1_sums[18][54] [5:0] }), .sum({ \level_2_sums[18][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[18][27] [6:0] }), .b({ \level_2_sums[18][26] [6:0] }), .sum({ \level_3_sums[18][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[18][13] [7:0] }),
     .b({ \level_3_sums[18][12] [7:0] }), .sum({ \level_4_sums[18][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[113] [4:0] }), .sum({ \level_1_sums[18][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[115] [4:0] }), .sum({ \level_1_sums[18][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[18][57] [5:0] }),
     .b({ \level_1_sums[18][56] [5:0] }), .sum({ \level_2_sums[18][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[117] [4:0] }), .sum({ \level_1_sums[18][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[119] [4:0] }), .sum({ \level_1_sums[18][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[18][59] [5:0] }),
     .b({ \level_1_sums[18][58] [5:0] }), .sum({ \level_2_sums[18][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[18][29] [6:0] }), .b({ \level_2_sums[18][28] [6:0] }), .sum({ \level_3_sums[18][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[121] [4:0] }), .sum({ \level_1_sums[18][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[123] [4:0] }), .sum({ \level_1_sums[18][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[18][61] [5:0] }),
     .b({ \level_1_sums[18][60] [5:0] }), .sum({ \level_2_sums[18][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[125] [4:0] }), .sum({ \level_1_sums[18][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[127] [4:0] }), .sum({ \level_1_sums[18][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[18][63] [5:0] }),
     .b({ \level_1_sums[18][62] [5:0] }), .sum({ \level_2_sums[18][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[18][31] [6:0] }), .b({ \level_2_sums[18][30] [6:0] }), .sum({ \level_3_sums[18][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[18][15] [7:0] }),
     .b({ \level_3_sums[18][14] [7:0] }), .sum({ \level_4_sums[18][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[18][7] [8:0] }),
     .b({ \level_4_sums[18][6] [8:0] }), .sum({ \level_5_sums[18][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[18][3] [9:0] }),
     .b({ \level_5_sums[18][2] [9:0] }), .sum({ \level_6_sums[18][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[18][1] [9:0] }),
     .b({ \level_6_sums[18][0] [9:0] }), .sum({ \level_7_sums[18][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[129] [4:0] }), .sum({ \level_1_sums[18][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[131] [4:0] }), .sum({ \level_1_sums[18][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[18][65] [5:0] }),
     .b({ \level_1_sums[18][64] [5:0] }), .sum({ \level_2_sums[18][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[133] [4:0] }), .sum({ \level_1_sums[18][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[135] [4:0] }), .sum({ \level_1_sums[18][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[18][67] [5:0] }),
     .b({ \level_1_sums[18][66] [5:0] }), .sum({ \level_2_sums[18][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[18][33] [6:0] }), .b({ \level_2_sums[18][32] [6:0] }), .sum({ \level_3_sums[18][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[137] [4:0] }), .sum({ \level_1_sums[18][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[139] [4:0] }), .sum({ \level_1_sums[18][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[18][69] [5:0] }),
     .b({ \level_1_sums[18][68] [5:0] }), .sum({ \level_2_sums[18][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[141] [4:0] }), .sum({ \level_1_sums[18][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[143] [4:0] }), .sum({ \level_1_sums[18][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[18][71] [5:0] }),
     .b({ \level_1_sums[18][70] [5:0] }), .sum({ \level_2_sums[18][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[18][35] [6:0] }), .b({ \level_2_sums[18][34] [6:0] }), .sum({ \level_3_sums[18][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[18][17] [7:0] }),
     .b({ \level_3_sums[18][16] [7:0] }), .sum({ \level_4_sums[18][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[145] [4:0] }), .sum({ \level_1_sums[18][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[147] [4:0] }), .sum({ \level_1_sums[18][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[18][73] [5:0] }),
     .b({ \level_1_sums[18][72] [5:0] }), .sum({ \level_2_sums[18][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[149] [4:0] }), .sum({ \level_1_sums[18][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[151] [4:0] }), .sum({ \level_1_sums[18][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[18][75] [5:0] }),
     .b({ \level_1_sums[18][74] [5:0] }), .sum({ \level_2_sums[18][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[18][37] [6:0] }), .b({ \level_2_sums[18][36] [6:0] }), .sum({ \level_3_sums[18][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[153] [4:0] }), .sum({ \level_1_sums[18][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[155] [4:0] }), .sum({ \level_1_sums[18][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[18][77] [5:0] }),
     .b({ \level_1_sums[18][76] [5:0] }), .sum({ \level_2_sums[18][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[157] [4:0] }), .sum({ \level_1_sums[18][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[159] [4:0] }), .sum({ \level_1_sums[18][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[18][79] [5:0] }),
     .b({ \level_1_sums[18][78] [5:0] }), .sum({ \level_2_sums[18][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[18][39] [6:0] }), .b({ \level_2_sums[18][38] [6:0] }), .sum({ \level_3_sums[18][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[18][19] [7:0] }),
     .b({ \level_3_sums[18][18] [7:0] }), .sum({ \level_4_sums[18][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[18][9] [8:0] }),
     .b({ \level_4_sums[18][8] [8:0] }), .sum({ \level_5_sums[18][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[161] [4:0] }), .sum({ \level_1_sums[18][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[163] [4:0] }), .sum({ \level_1_sums[18][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[18][81] [5:0] }),
     .b({ \level_1_sums[18][80] [5:0] }), .sum({ \level_2_sums[18][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[165] [4:0] }), .sum({ \level_1_sums[18][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[167] [4:0] }), .sum({ \level_1_sums[18][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[18][83] [5:0] }),
     .b({ \level_1_sums[18][82] [5:0] }), .sum({ \level_2_sums[18][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[18][41] [6:0] }), .b({ \level_2_sums[18][40] [6:0] }), .sum({ \level_3_sums[18][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[169] [4:0] }), .sum({ \level_1_sums[18][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[171] [4:0] }), .sum({ \level_1_sums[18][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[18][85] [5:0] }),
     .b({ \level_1_sums[18][84] [5:0] }), .sum({ \level_2_sums[18][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[173] [4:0] }), .sum({ \level_1_sums[18][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[175] [4:0] }), .sum({ \level_1_sums[18][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[18][87] [5:0] }),
     .b({ \level_1_sums[18][86] [5:0] }), .sum({ \level_2_sums[18][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[18][43] [6:0] }), .b({ \level_2_sums[18][42] [6:0] }), .sum({ \level_3_sums[18][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[18][21] [7:0] }),
     .b({ \level_3_sums[18][20] [7:0] }), .sum({ \level_4_sums[18][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[177] [4:0] }), .sum({ \level_1_sums[18][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[179] [4:0] }), .sum({ \level_1_sums[18][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[18][89] [5:0] }),
     .b({ \level_1_sums[18][88] [5:0] }), .sum({ \level_2_sums[18][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[181] [4:0] }), .sum({ \level_1_sums[18][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[183] [4:0] }), .sum({ \level_1_sums[18][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[18][91] [5:0] }),
     .b({ \level_1_sums[18][90] [5:0] }), .sum({ \level_2_sums[18][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[18][45] [6:0] }), .b({ \level_2_sums[18][44] [6:0] }), .sum({ \level_3_sums[18][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[185] [4:0] }), .sum({ \level_1_sums[18][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[187] [4:0] }), .sum({ \level_1_sums[18][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[18][93] [5:0] }),
     .b({ \level_1_sums[18][92] [5:0] }), .sum({ \level_2_sums[18][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[189] [4:0] }), .sum({ \level_1_sums[18][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[191] [4:0] }), .sum({ \level_1_sums[18][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[18][95] [5:0] }),
     .b({ \level_1_sums[18][94] [5:0] }), .sum({ \level_2_sums[18][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[18][47] [6:0] }), .b({ \level_2_sums[18][46] [6:0] }), .sum({ \level_3_sums[18][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[18][23] [7:0] }),
     .b({ \level_3_sums[18][22] [7:0] }), .sum({ \level_4_sums[18][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[18][11] [8:0] }),
     .b({ \level_4_sums[18][10] [8:0] }), .sum({ \level_5_sums[18][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[18][5] [9:0] }),
     .b({ \level_5_sums[18][4] [9:0] }), .sum({ \level_6_sums[18][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[193] [4:0] }), .sum({ \level_1_sums[18][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[195] [4:0] }), .sum({ \level_1_sums[18][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[18][97] [5:0] }),
     .b({ \level_1_sums[18][96] [5:0] }), .sum({ \level_2_sums[18][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[197] [4:0] }), .sum({ \level_1_sums[18][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[199] [4:0] }), .sum({ \level_1_sums[18][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[18][99] [5:0] }),
     .b({ \level_1_sums[18][98] [5:0] }), .sum({ \level_2_sums[18][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[18][49] [6:0] }), .b({ \level_2_sums[18][48] [6:0] }), .sum({ \level_3_sums[18][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[201] [4:0] }), .sum({ \level_1_sums[18][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[203] [4:0] }), .sum({ \level_1_sums[18][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[18][101] [5:0] }),
     .b({ \level_1_sums[18][100] [5:0] }), .sum({ \level_2_sums[18][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[205] [4:0] }), .sum({ \level_1_sums[18][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[207] [4:0] }), .sum({ \level_1_sums[18][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[18][103] [5:0] }),
     .b({ \level_1_sums[18][102] [5:0] }), .sum({ \level_2_sums[18][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[18][51] [6:0] }), .b({ \level_2_sums[18][50] [6:0] }), .sum({ \level_3_sums[18][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[18][25] [7:0] }),
     .b({ \level_3_sums[18][24] [7:0] }), .sum({ \level_4_sums[18][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[209] [4:0] }), .sum({ \level_1_sums[18][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[211] [4:0] }), .sum({ \level_1_sums[18][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[18][105] [5:0] }),
     .b({ \level_1_sums[18][104] [5:0] }), .sum({ \level_2_sums[18][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[213] [4:0] }), .sum({ \level_1_sums[18][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[215] [4:0] }), .sum({ \level_1_sums[18][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[18][107] [5:0] }),
     .b({ \level_1_sums[18][106] [5:0] }), .sum({ \level_2_sums[18][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[18][53] [6:0] }), .b({ \level_2_sums[18][52] [6:0] }), .sum({ \level_3_sums[18][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[217] [4:0] }), .sum({ \level_1_sums[18][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[219] [4:0] }), .sum({ \level_1_sums[18][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[18][109] [5:0] }),
     .b({ \level_1_sums[18][108] [5:0] }), .sum({ \level_2_sums[18][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[221] [4:0] }), .sum({ \level_1_sums[18][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[223] [4:0] }), .sum({ \level_1_sums[18][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[18][111] [5:0] }),
     .b({ \level_1_sums[18][110] [5:0] }), .sum({ \level_2_sums[18][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[18][55] [6:0] }), .b({ \level_2_sums[18][54] [6:0] }), .sum({ \level_3_sums[18][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[18][27] [7:0] }),
     .b({ \level_3_sums[18][26] [7:0] }), .sum({ \level_4_sums[18][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[18][13] [8:0] }),
     .b({ \level_4_sums[18][12] [8:0] }), .sum({ \level_5_sums[18][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[225] [4:0] }), .sum({ \level_1_sums[18][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[227] [4:0] }), .sum({ \level_1_sums[18][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[18][113] [5:0] }),
     .b({ \level_1_sums[18][112] [5:0] }), .sum({ \level_2_sums[18][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[229] [4:0] }), .sum({ \level_1_sums[18][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[231] [4:0] }), .sum({ \level_1_sums[18][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[18][115] [5:0] }),
     .b({ \level_1_sums[18][114] [5:0] }), .sum({ \level_2_sums[18][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[18][57] [6:0] }), .b({ \level_2_sums[18][56] [6:0] }), .sum({ \level_3_sums[18][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[233] [4:0] }), .sum({ \level_1_sums[18][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[235] [4:0] }), .sum({ \level_1_sums[18][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[18][117] [5:0] }),
     .b({ \level_1_sums[18][116] [5:0] }), .sum({ \level_2_sums[18][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[237] [4:0] }), .sum({ \level_1_sums[18][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[239] [4:0] }), .sum({ \level_1_sums[18][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[18][119] [5:0] }),
     .b({ \level_1_sums[18][118] [5:0] }), .sum({ \level_2_sums[18][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[18][59] [6:0] }), .b({ \level_2_sums[18][58] [6:0] }), .sum({ \level_3_sums[18][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[18][29] [7:0] }),
     .b({ \level_3_sums[18][28] [7:0] }), .sum({ \level_4_sums[18][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[241] [4:0] }), .sum({ \level_1_sums[18][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[243] [4:0] }), .sum({ \level_1_sums[18][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[18][121] [5:0] }),
     .b({ \level_1_sums[18][120] [5:0] }), .sum({ \level_2_sums[18][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[245] [4:0] }), .sum({ \level_1_sums[18][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[247] [4:0] }), .sum({ \level_1_sums[18][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[18][123] [5:0] }),
     .b({ \level_1_sums[18][122] [5:0] }), .sum({ \level_2_sums[18][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[18][61] [6:0] }), .b({ \level_2_sums[18][60] [6:0] }), .sum({ \level_3_sums[18][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[249] [4:0] }), .sum({ \level_1_sums[18][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[251] [4:0] }), .sum({ \level_1_sums[18][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[18][125] [5:0] }),
     .b({ \level_1_sums[18][124] [5:0] }), .sum({ \level_2_sums[18][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[253] [4:0] }), .sum({ \level_1_sums[18][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[18].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[18].product_terms[255] [4:0] }), .sum({ \level_1_sums[18][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[18][127] [5:0] }),
     .b({ \level_1_sums[18][126] [5:0] }), .sum({ \level_2_sums[18][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[18][63] [6:0] }), .b({ \level_2_sums[18][62] [6:0] }), .sum({ \level_3_sums[18][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[18][31] [7:0] }),
     .b({ \level_3_sums[18][30] [7:0] }), .sum({ \level_4_sums[18][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[18][15] [8:0] }),
     .b({ \level_4_sums[18][14] [8:0] }), .sum({ \level_5_sums[18][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[18][7] [9:0] }),
     .b({ \level_5_sums[18][6] [9:0] }), .sum({ \level_6_sums[18][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[18][3] [9:0] }),
     .b({ \level_6_sums[18][2] [9:0] }), .sum({ \level_7_sums[18][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[18].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[18][0] [9:0] }),
     .b({ \level_7_sums[18][1] [9:0] }), .sum({ \level_8_sums[18] [9:0] }));
  ReLU_10bit \dot_product_and_ReLU[19].relu_inst (.in_data({ \final_sums[19] [9:0] }), .out_data({ \out_sig[19] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[1].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[0] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[1] [4:0] }), .sum({ \level_1_sums[19][0] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[3].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[2] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[3] [4:0] }), .sum({ \level_1_sums[19][1] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[3].adder_quads.adder_inst (.a({ \level_1_sums[19][1] [5:0] }),
     .b({ \level_1_sums[19][0] [5:0] }), .sum({ \level_2_sums[19][0] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[5].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[4] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[5] [4:0] }), .sum({ \level_1_sums[19][2] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[7].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[6] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[7] [4:0] }), .sum({ \level_1_sums[19][3] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[7].adder_quads.adder_inst (.a({ \level_1_sums[19][3] [5:0] }),
     .b({ \level_1_sums[19][2] [5:0] }), .sum({ \level_2_sums[19][1] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[7].adder_octets.adder_inst (.a({ \level_2_sums[19][1] [6:0] }),
     .b({ \level_2_sums[19][0] [6:0] }), .sum({ \level_3_sums[19][0] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[9].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[8] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[9] [4:0] }), .sum({ \level_1_sums[19][4] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[11].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[10] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[11] [4:0] }), .sum({ \level_1_sums[19][5] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[11].adder_quads.adder_inst (.a({ \level_1_sums[19][5] [5:0] }),
     .b({ \level_1_sums[19][4] [5:0] }), .sum({ \level_2_sums[19][2] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[13].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[12] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[13] [4:0] }), .sum({ \level_1_sums[19][6] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[15].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[14] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[15] [4:0] }), .sum({ \level_1_sums[19][7] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[15].adder_quads.adder_inst (.a({ \level_1_sums[19][7] [5:0] }),
     .b({ \level_1_sums[19][6] [5:0] }), .sum({ \level_2_sums[19][3] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[15].adder_octets.adder_inst (.a({ \level_2_sums[19][3] [6:0] }),
     .b({ \level_2_sums[19][2] [6:0] }), .sum({ \level_3_sums[19][1] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[15].adder_16s.adder_inst (.a({ \level_3_sums[19][1] [7:0] }),
     .b({ \level_3_sums[19][0] [7:0] }), .sum({ \level_4_sums[19][0] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[17].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[16] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[17] [4:0] }), .sum({ \level_1_sums[19][8] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[19].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[18] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[19] [4:0] }), .sum({ \level_1_sums[19][9] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[19].adder_quads.adder_inst (.a({ \level_1_sums[19][9] [5:0] }),
     .b({ \level_1_sums[19][8] [5:0] }), .sum({ \level_2_sums[19][4] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[21].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[20] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[21] [4:0] }), .sum({ \level_1_sums[19][10] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[23].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[22] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[23] [4:0] }), .sum({ \level_1_sums[19][11] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[23].adder_quads.adder_inst (.a({ \level_1_sums[19][11] [5:0] }),
     .b({ \level_1_sums[19][10] [5:0] }), .sum({ \level_2_sums[19][5] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[23].adder_octets.adder_inst (.a({ \level_2_sums[19][5] [6:0] }),
     .b({ \level_2_sums[19][4] [6:0] }), .sum({ \level_3_sums[19][2] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[25].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[24] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[25] [4:0] }), .sum({ \level_1_sums[19][12] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[27].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[26] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[27] [4:0] }), .sum({ \level_1_sums[19][13] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[27].adder_quads.adder_inst (.a({ \level_1_sums[19][13] [5:0] }),
     .b({ \level_1_sums[19][12] [5:0] }), .sum({ \level_2_sums[19][6] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[29].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[28] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[29] [4:0] }), .sum({ \level_1_sums[19][14] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[31].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[30] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[31] [4:0] }), .sum({ \level_1_sums[19][15] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[31].adder_quads.adder_inst (.a({ \level_1_sums[19][15] [5:0] }),
     .b({ \level_1_sums[19][14] [5:0] }), .sum({ \level_2_sums[19][7] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[31].adder_octets.adder_inst (.a({ \level_2_sums[19][7] [6:0] }),
     .b({ \level_2_sums[19][6] [6:0] }), .sum({ \level_3_sums[19][3] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[31].adder_16s.adder_inst (.a({ \level_3_sums[19][3] [7:0] }),
     .b({ \level_3_sums[19][2] [7:0] }), .sum({ \level_4_sums[19][1] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[31].adder_32s.adder_inst (.a({ \level_4_sums[19][1] [8:0] }),
     .b({ \level_4_sums[19][0] [8:0] }), .sum({ \level_5_sums[19][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[33].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[32] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[33] [4:0] }), .sum({ \level_1_sums[19][16] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[35].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[34] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[35] [4:0] }), .sum({ \level_1_sums[19][17] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[35].adder_quads.adder_inst (.a({ \level_1_sums[19][17] [5:0] }),
     .b({ \level_1_sums[19][16] [5:0] }), .sum({ \level_2_sums[19][8] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[37].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[36] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[37] [4:0] }), .sum({ \level_1_sums[19][18] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[39].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[38] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[39] [4:0] }), .sum({ \level_1_sums[19][19] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[39].adder_quads.adder_inst (.a({ \level_1_sums[19][19] [5:0] }),
     .b({ \level_1_sums[19][18] [5:0] }), .sum({ \level_2_sums[19][9] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[39].adder_octets.adder_inst (.a({ \level_2_sums[19][9] [6:0] }),
     .b({ \level_2_sums[19][8] [6:0] }), .sum({ \level_3_sums[19][4] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[41].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[40] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[41] [4:0] }), .sum({ \level_1_sums[19][20] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[43].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[42] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[43] [4:0] }), .sum({ \level_1_sums[19][21] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[43].adder_quads.adder_inst (.a({ \level_1_sums[19][21] [5:0] }),
     .b({ \level_1_sums[19][20] [5:0] }), .sum({ \level_2_sums[19][10] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[45].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[44] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[45] [4:0] }), .sum({ \level_1_sums[19][22] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[47].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[46] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[47] [4:0] }), .sum({ \level_1_sums[19][23] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[47].adder_quads.adder_inst (.a({ \level_1_sums[19][23] [5:0] }),
     .b({ \level_1_sums[19][22] [5:0] }), .sum({ \level_2_sums[19][11] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[47].adder_octets.adder_inst (.a({ \level_2_sums[19][11] [6:0] }),
     .b({ \level_2_sums[19][10] [6:0] }), .sum({ \level_3_sums[19][5] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[47].adder_16s.adder_inst (.a({ \level_3_sums[19][5] [7:0] }),
     .b({ \level_3_sums[19][4] [7:0] }), .sum({ \level_4_sums[19][2] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[49].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[48] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[49] [4:0] }), .sum({ \level_1_sums[19][24] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[51].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[50] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[51] [4:0] }), .sum({ \level_1_sums[19][25] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[51].adder_quads.adder_inst (.a({ \level_1_sums[19][25] [5:0] }),
     .b({ \level_1_sums[19][24] [5:0] }), .sum({ \level_2_sums[19][12] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[53].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[52] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[53] [4:0] }), .sum({ \level_1_sums[19][26] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[55].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[54] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[55] [4:0] }), .sum({ \level_1_sums[19][27] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[55].adder_quads.adder_inst (.a({ \level_1_sums[19][27] [5:0] }),
     .b({ \level_1_sums[19][26] [5:0] }), .sum({ \level_2_sums[19][13] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[55].adder_octets.adder_inst (.a({ \level_2_sums[19][13] [6:0] }),
     .b({ \level_2_sums[19][12] [6:0] }), .sum({ \level_3_sums[19][6] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[57].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[56] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[57] [4:0] }), .sum({ \level_1_sums[19][28] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[59].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[58] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[59] [4:0] }), .sum({ \level_1_sums[19][29] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[59].adder_quads.adder_inst (.a({ \level_1_sums[19][29] [5:0] }),
     .b({ \level_1_sums[19][28] [5:0] }), .sum({ \level_2_sums[19][14] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[61].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[60] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[61] [4:0] }), .sum({ \level_1_sums[19][30] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[62] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[63] [4:0] }), .sum({ \level_1_sums[19][31] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_quads.adder_inst (.a({ \level_1_sums[19][31] [5:0] }),
     .b({ \level_1_sums[19][30] [5:0] }), .sum({ \level_2_sums[19][15] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_octets.adder_inst (.a({ \level_2_sums[19][15] [6:0] }),
     .b({ \level_2_sums[19][14] [6:0] }), .sum({ \level_3_sums[19][7] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_16s.adder_inst (.a({ \level_3_sums[19][7] [7:0] }),
     .b({ \level_3_sums[19][6] [7:0] }), .sum({ \level_4_sums[19][3] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_32s.adder_inst (.a({ \level_4_sums[19][3] [8:0] }),
     .b({ \level_4_sums[19][2] [8:0] }), .sum({ \level_5_sums[19][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[63].adder_64s.adder_inst (.a({ \level_5_sums[19][1] [9:0] }),
     .b({ \level_5_sums[19][0] [9:0] }), .sum({ \level_6_sums[19][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[65].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[64] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[65] [4:0] }), .sum({ \level_1_sums[19][32] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[67].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[66] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[67] [4:0] }), .sum({ \level_1_sums[19][33] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[67].adder_quads.adder_inst (.a({ \level_1_sums[19][33] [5:0] }),
     .b({ \level_1_sums[19][32] [5:0] }), .sum({ \level_2_sums[19][16] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[69].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[68] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[69] [4:0] }), .sum({ \level_1_sums[19][34] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[71].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[70] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[71] [4:0] }), .sum({ \level_1_sums[19][35] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[71].adder_quads.adder_inst (.a({ \level_1_sums[19][35] [5:0] }),
     .b({ \level_1_sums[19][34] [5:0] }), .sum({ \level_2_sums[19][17] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[71].adder_octets.adder_inst (.a({ \level_2_sums[19][17] [6:0] }),
     .b({ \level_2_sums[19][16] [6:0] }), .sum({ \level_3_sums[19][8] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[73].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[72] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[73] [4:0] }), .sum({ \level_1_sums[19][36] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[75].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[74] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[75] [4:0] }), .sum({ \level_1_sums[19][37] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[75].adder_quads.adder_inst (.a({ \level_1_sums[19][37] [5:0] }),
     .b({ \level_1_sums[19][36] [5:0] }), .sum({ \level_2_sums[19][18] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[77].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[76] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[77] [4:0] }), .sum({ \level_1_sums[19][38] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[79].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[78] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[79] [4:0] }), .sum({ \level_1_sums[19][39] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[79].adder_quads.adder_inst (.a({ \level_1_sums[19][39] [5:0] }),
     .b({ \level_1_sums[19][38] [5:0] }), .sum({ \level_2_sums[19][19] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[79].adder_octets.adder_inst (.a({ \level_2_sums[19][19] [6:0] }),
     .b({ \level_2_sums[19][18] [6:0] }), .sum({ \level_3_sums[19][9] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[79].adder_16s.adder_inst (.a({ \level_3_sums[19][9] [7:0] }),
     .b({ \level_3_sums[19][8] [7:0] }), .sum({ \level_4_sums[19][4] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[81].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[80] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[81] [4:0] }), .sum({ \level_1_sums[19][40] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[83].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[82] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[83] [4:0] }), .sum({ \level_1_sums[19][41] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[83].adder_quads.adder_inst (.a({ \level_1_sums[19][41] [5:0] }),
     .b({ \level_1_sums[19][40] [5:0] }), .sum({ \level_2_sums[19][20] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[85].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[84] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[85] [4:0] }), .sum({ \level_1_sums[19][42] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[87].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[86] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[87] [4:0] }), .sum({ \level_1_sums[19][43] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[87].adder_quads.adder_inst (.a({ \level_1_sums[19][43] [5:0] }),
     .b({ \level_1_sums[19][42] [5:0] }), .sum({ \level_2_sums[19][21] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[87].adder_octets.adder_inst (.a({ \level_2_sums[19][21] [6:0] }),
     .b({ \level_2_sums[19][20] [6:0] }), .sum({ \level_3_sums[19][10] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[89].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[88] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[89] [4:0] }), .sum({ \level_1_sums[19][44] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[91].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[90] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[91] [4:0] }), .sum({ \level_1_sums[19][45] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[91].adder_quads.adder_inst (.a({ \level_1_sums[19][45] [5:0] }),
     .b({ \level_1_sums[19][44] [5:0] }), .sum({ \level_2_sums[19][22] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[93].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[92] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[93] [4:0] }), .sum({ \level_1_sums[19][46] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[95].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[94] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[95] [4:0] }), .sum({ \level_1_sums[19][47] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[95].adder_quads.adder_inst (.a({ \level_1_sums[19][47] [5:0] }),
     .b({ \level_1_sums[19][46] [5:0] }), .sum({ \level_2_sums[19][23] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[95].adder_octets.adder_inst (.a({ \level_2_sums[19][23] [6:0] }),
     .b({ \level_2_sums[19][22] [6:0] }), .sum({ \level_3_sums[19][11] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[95].adder_16s.adder_inst (.a({ \level_3_sums[19][11] [7:0] }),
     .b({ \level_3_sums[19][10] [7:0] }), .sum({ \level_4_sums[19][5] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[95].adder_32s.adder_inst (.a({ \level_4_sums[19][5] [8:0] }),
     .b({ \level_4_sums[19][4] [8:0] }), .sum({ \level_5_sums[19][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[97].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[96] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[97] [4:0] }), .sum({ \level_1_sums[19][48] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[99].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[98] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[99] [4:0] }), .sum({ \level_1_sums[19][49] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[99].adder_quads.adder_inst (.a({ \level_1_sums[19][49] [5:0] }),
     .b({ \level_1_sums[19][48] [5:0] }), .sum({ \level_2_sums[19][24] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[101].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[100] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[101] [4:0] }), .sum({ \level_1_sums[19][50] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[103].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[102] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[103] [4:0] }), .sum({ \level_1_sums[19][51] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[103].adder_quads.adder_inst (.a({ \level_1_sums[19][51] [5:0] }),
     .b({ \level_1_sums[19][50] [5:0] }), .sum({ \level_2_sums[19][25] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[103].adder_octets.adder_inst (
    .a({ \level_2_sums[19][25] [6:0] }), .b({ \level_2_sums[19][24] [6:0] }), .sum({ \level_3_sums[19][12] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[105].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[104] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[105] [4:0] }), .sum({ \level_1_sums[19][52] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[107].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[106] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[107] [4:0] }), .sum({ \level_1_sums[19][53] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[107].adder_quads.adder_inst (.a({ \level_1_sums[19][53] [5:0] }),
     .b({ \level_1_sums[19][52] [5:0] }), .sum({ \level_2_sums[19][26] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[109].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[108] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[109] [4:0] }), .sum({ \level_1_sums[19][54] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[111].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[110] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[111] [4:0] }), .sum({ \level_1_sums[19][55] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[111].adder_quads.adder_inst (.a({ \level_1_sums[19][55] [5:0] }),
     .b({ \level_1_sums[19][54] [5:0] }), .sum({ \level_2_sums[19][27] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[111].adder_octets.adder_inst (
    .a({ \level_2_sums[19][27] [6:0] }), .b({ \level_2_sums[19][26] [6:0] }), .sum({ \level_3_sums[19][13] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[111].adder_16s.adder_inst (.a({ \level_3_sums[19][13] [7:0] }),
     .b({ \level_3_sums[19][12] [7:0] }), .sum({ \level_4_sums[19][6] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[113].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[112] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[113] [4:0] }), .sum({ \level_1_sums[19][56] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[115].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[114] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[115] [4:0] }), .sum({ \level_1_sums[19][57] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[115].adder_quads.adder_inst (.a({ \level_1_sums[19][57] [5:0] }),
     .b({ \level_1_sums[19][56] [5:0] }), .sum({ \level_2_sums[19][28] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[117].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[116] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[117] [4:0] }), .sum({ \level_1_sums[19][58] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[119].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[118] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[119] [4:0] }), .sum({ \level_1_sums[19][59] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[119].adder_quads.adder_inst (.a({ \level_1_sums[19][59] [5:0] }),
     .b({ \level_1_sums[19][58] [5:0] }), .sum({ \level_2_sums[19][29] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[119].adder_octets.adder_inst (
    .a({ \level_2_sums[19][29] [6:0] }), .b({ \level_2_sums[19][28] [6:0] }), .sum({ \level_3_sums[19][14] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[121].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[120] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[121] [4:0] }), .sum({ \level_1_sums[19][60] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[123].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[122] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[123] [4:0] }), .sum({ \level_1_sums[19][61] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[123].adder_quads.adder_inst (.a({ \level_1_sums[19][61] [5:0] }),
     .b({ \level_1_sums[19][60] [5:0] }), .sum({ \level_2_sums[19][30] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[125].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[124] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[125] [4:0] }), .sum({ \level_1_sums[19][62] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[126] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[127] [4:0] }), .sum({ \level_1_sums[19][63] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_quads.adder_inst (.a({ \level_1_sums[19][63] [5:0] }),
     .b({ \level_1_sums[19][62] [5:0] }), .sum({ \level_2_sums[19][31] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_octets.adder_inst (
    .a({ \level_2_sums[19][31] [6:0] }), .b({ \level_2_sums[19][30] [6:0] }), .sum({ \level_3_sums[19][15] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_16s.adder_inst (.a({ \level_3_sums[19][15] [7:0] }),
     .b({ \level_3_sums[19][14] [7:0] }), .sum({ \level_4_sums[19][7] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_32s.adder_inst (.a({ \level_4_sums[19][7] [8:0] }),
     .b({ \level_4_sums[19][6] [8:0] }), .sum({ \level_5_sums[19][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_64s.adder_inst (.a({ \level_5_sums[19][3] [9:0] }),
     .b({ \level_5_sums[19][2] [9:0] }), .sum({ \level_6_sums[19][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[127].adder_128s.adder_inst (.a({ \level_6_sums[19][1] [9:0] }),
     .b({ \level_6_sums[19][0] [9:0] }), .sum({ \level_7_sums[19][0] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[129].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[128] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[129] [4:0] }), .sum({ \level_1_sums[19][64] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[131].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[130] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[131] [4:0] }), .sum({ \level_1_sums[19][65] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[131].adder_quads.adder_inst (.a({ \level_1_sums[19][65] [5:0] }),
     .b({ \level_1_sums[19][64] [5:0] }), .sum({ \level_2_sums[19][32] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[133].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[132] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[133] [4:0] }), .sum({ \level_1_sums[19][66] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[135].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[134] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[135] [4:0] }), .sum({ \level_1_sums[19][67] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[135].adder_quads.adder_inst (.a({ \level_1_sums[19][67] [5:0] }),
     .b({ \level_1_sums[19][66] [5:0] }), .sum({ \level_2_sums[19][33] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[135].adder_octets.adder_inst (
    .a({ \level_2_sums[19][33] [6:0] }), .b({ \level_2_sums[19][32] [6:0] }), .sum({ \level_3_sums[19][16] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[137].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[136] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[137] [4:0] }), .sum({ \level_1_sums[19][68] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[139].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[138] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[139] [4:0] }), .sum({ \level_1_sums[19][69] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[139].adder_quads.adder_inst (.a({ \level_1_sums[19][69] [5:0] }),
     .b({ \level_1_sums[19][68] [5:0] }), .sum({ \level_2_sums[19][34] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[141].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[140] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[141] [4:0] }), .sum({ \level_1_sums[19][70] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[143].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[142] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[143] [4:0] }), .sum({ \level_1_sums[19][71] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[143].adder_quads.adder_inst (.a({ \level_1_sums[19][71] [5:0] }),
     .b({ \level_1_sums[19][70] [5:0] }), .sum({ \level_2_sums[19][35] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[143].adder_octets.adder_inst (
    .a({ \level_2_sums[19][35] [6:0] }), .b({ \level_2_sums[19][34] [6:0] }), .sum({ \level_3_sums[19][17] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[143].adder_16s.adder_inst (.a({ \level_3_sums[19][17] [7:0] }),
     .b({ \level_3_sums[19][16] [7:0] }), .sum({ \level_4_sums[19][8] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[145].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[144] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[145] [4:0] }), .sum({ \level_1_sums[19][72] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[147].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[146] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[147] [4:0] }), .sum({ \level_1_sums[19][73] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[147].adder_quads.adder_inst (.a({ \level_1_sums[19][73] [5:0] }),
     .b({ \level_1_sums[19][72] [5:0] }), .sum({ \level_2_sums[19][36] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[149].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[148] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[149] [4:0] }), .sum({ \level_1_sums[19][74] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[151].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[150] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[151] [4:0] }), .sum({ \level_1_sums[19][75] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[151].adder_quads.adder_inst (.a({ \level_1_sums[19][75] [5:0] }),
     .b({ \level_1_sums[19][74] [5:0] }), .sum({ \level_2_sums[19][37] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[151].adder_octets.adder_inst (
    .a({ \level_2_sums[19][37] [6:0] }), .b({ \level_2_sums[19][36] [6:0] }), .sum({ \level_3_sums[19][18] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[153].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[152] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[153] [4:0] }), .sum({ \level_1_sums[19][76] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[155].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[154] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[155] [4:0] }), .sum({ \level_1_sums[19][77] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[155].adder_quads.adder_inst (.a({ \level_1_sums[19][77] [5:0] }),
     .b({ \level_1_sums[19][76] [5:0] }), .sum({ \level_2_sums[19][38] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[157].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[156] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[157] [4:0] }), .sum({ \level_1_sums[19][78] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[159].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[158] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[159] [4:0] }), .sum({ \level_1_sums[19][79] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[159].adder_quads.adder_inst (.a({ \level_1_sums[19][79] [5:0] }),
     .b({ \level_1_sums[19][78] [5:0] }), .sum({ \level_2_sums[19][39] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[159].adder_octets.adder_inst (
    .a({ \level_2_sums[19][39] [6:0] }), .b({ \level_2_sums[19][38] [6:0] }), .sum({ \level_3_sums[19][19] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[159].adder_16s.adder_inst (.a({ \level_3_sums[19][19] [7:0] }),
     .b({ \level_3_sums[19][18] [7:0] }), .sum({ \level_4_sums[19][9] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[159].adder_32s.adder_inst (.a({ \level_4_sums[19][9] [8:0] }),
     .b({ \level_4_sums[19][8] [8:0] }), .sum({ \level_5_sums[19][4] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[161].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[160] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[161] [4:0] }), .sum({ \level_1_sums[19][80] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[163].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[162] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[163] [4:0] }), .sum({ \level_1_sums[19][81] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[163].adder_quads.adder_inst (.a({ \level_1_sums[19][81] [5:0] }),
     .b({ \level_1_sums[19][80] [5:0] }), .sum({ \level_2_sums[19][40] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[165].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[164] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[165] [4:0] }), .sum({ \level_1_sums[19][82] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[167].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[166] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[167] [4:0] }), .sum({ \level_1_sums[19][83] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[167].adder_quads.adder_inst (.a({ \level_1_sums[19][83] [5:0] }),
     .b({ \level_1_sums[19][82] [5:0] }), .sum({ \level_2_sums[19][41] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[167].adder_octets.adder_inst (
    .a({ \level_2_sums[19][41] [6:0] }), .b({ \level_2_sums[19][40] [6:0] }), .sum({ \level_3_sums[19][20] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[169].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[168] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[169] [4:0] }), .sum({ \level_1_sums[19][84] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[171].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[170] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[171] [4:0] }), .sum({ \level_1_sums[19][85] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[171].adder_quads.adder_inst (.a({ \level_1_sums[19][85] [5:0] }),
     .b({ \level_1_sums[19][84] [5:0] }), .sum({ \level_2_sums[19][42] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[173].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[172] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[173] [4:0] }), .sum({ \level_1_sums[19][86] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[175].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[174] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[175] [4:0] }), .sum({ \level_1_sums[19][87] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[175].adder_quads.adder_inst (.a({ \level_1_sums[19][87] [5:0] }),
     .b({ \level_1_sums[19][86] [5:0] }), .sum({ \level_2_sums[19][43] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[175].adder_octets.adder_inst (
    .a({ \level_2_sums[19][43] [6:0] }), .b({ \level_2_sums[19][42] [6:0] }), .sum({ \level_3_sums[19][21] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[175].adder_16s.adder_inst (.a({ \level_3_sums[19][21] [7:0] }),
     .b({ \level_3_sums[19][20] [7:0] }), .sum({ \level_4_sums[19][10] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[177].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[176] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[177] [4:0] }), .sum({ \level_1_sums[19][88] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[179].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[178] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[179] [4:0] }), .sum({ \level_1_sums[19][89] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[179].adder_quads.adder_inst (.a({ \level_1_sums[19][89] [5:0] }),
     .b({ \level_1_sums[19][88] [5:0] }), .sum({ \level_2_sums[19][44] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[181].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[180] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[181] [4:0] }), .sum({ \level_1_sums[19][90] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[183].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[182] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[183] [4:0] }), .sum({ \level_1_sums[19][91] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[183].adder_quads.adder_inst (.a({ \level_1_sums[19][91] [5:0] }),
     .b({ \level_1_sums[19][90] [5:0] }), .sum({ \level_2_sums[19][45] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[183].adder_octets.adder_inst (
    .a({ \level_2_sums[19][45] [6:0] }), .b({ \level_2_sums[19][44] [6:0] }), .sum({ \level_3_sums[19][22] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[185].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[184] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[185] [4:0] }), .sum({ \level_1_sums[19][92] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[187].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[186] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[187] [4:0] }), .sum({ \level_1_sums[19][93] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[187].adder_quads.adder_inst (.a({ \level_1_sums[19][93] [5:0] }),
     .b({ \level_1_sums[19][92] [5:0] }), .sum({ \level_2_sums[19][46] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[189].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[188] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[189] [4:0] }), .sum({ \level_1_sums[19][94] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[190] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[191] [4:0] }), .sum({ \level_1_sums[19][95] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_quads.adder_inst (.a({ \level_1_sums[19][95] [5:0] }),
     .b({ \level_1_sums[19][94] [5:0] }), .sum({ \level_2_sums[19][47] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_octets.adder_inst (
    .a({ \level_2_sums[19][47] [6:0] }), .b({ \level_2_sums[19][46] [6:0] }), .sum({ \level_3_sums[19][23] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_16s.adder_inst (.a({ \level_3_sums[19][23] [7:0] }),
     .b({ \level_3_sums[19][22] [7:0] }), .sum({ \level_4_sums[19][11] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_32s.adder_inst (.a({ \level_4_sums[19][11] [8:0] }),
     .b({ \level_4_sums[19][10] [8:0] }), .sum({ \level_5_sums[19][5] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[191].adder_64s.adder_inst (.a({ \level_5_sums[19][5] [9:0] }),
     .b({ \level_5_sums[19][4] [9:0] }), .sum({ \level_6_sums[19][2] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[193].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[192] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[193] [4:0] }), .sum({ \level_1_sums[19][96] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[195].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[194] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[195] [4:0] }), .sum({ \level_1_sums[19][97] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[195].adder_quads.adder_inst (.a({ \level_1_sums[19][97] [5:0] }),
     .b({ \level_1_sums[19][96] [5:0] }), .sum({ \level_2_sums[19][48] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[197].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[196] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[197] [4:0] }), .sum({ \level_1_sums[19][98] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[199].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[198] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[199] [4:0] }), .sum({ \level_1_sums[19][99] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[199].adder_quads.adder_inst (.a({ \level_1_sums[19][99] [5:0] }),
     .b({ \level_1_sums[19][98] [5:0] }), .sum({ \level_2_sums[19][49] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[199].adder_octets.adder_inst (
    .a({ \level_2_sums[19][49] [6:0] }), .b({ \level_2_sums[19][48] [6:0] }), .sum({ \level_3_sums[19][24] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[201].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[200] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[201] [4:0] }), .sum({ \level_1_sums[19][100] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[203].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[202] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[203] [4:0] }), .sum({ \level_1_sums[19][101] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[203].adder_quads.adder_inst (.a({ \level_1_sums[19][101] [5:0] }),
     .b({ \level_1_sums[19][100] [5:0] }), .sum({ \level_2_sums[19][50] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[205].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[204] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[205] [4:0] }), .sum({ \level_1_sums[19][102] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[207].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[206] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[207] [4:0] }), .sum({ \level_1_sums[19][103] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[207].adder_quads.adder_inst (.a({ \level_1_sums[19][103] [5:0] }),
     .b({ \level_1_sums[19][102] [5:0] }), .sum({ \level_2_sums[19][51] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[207].adder_octets.adder_inst (
    .a({ \level_2_sums[19][51] [6:0] }), .b({ \level_2_sums[19][50] [6:0] }), .sum({ \level_3_sums[19][25] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[207].adder_16s.adder_inst (.a({ \level_3_sums[19][25] [7:0] }),
     .b({ \level_3_sums[19][24] [7:0] }), .sum({ \level_4_sums[19][12] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[209].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[208] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[209] [4:0] }), .sum({ \level_1_sums[19][104] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[211].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[210] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[211] [4:0] }), .sum({ \level_1_sums[19][105] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[211].adder_quads.adder_inst (.a({ \level_1_sums[19][105] [5:0] }),
     .b({ \level_1_sums[19][104] [5:0] }), .sum({ \level_2_sums[19][52] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[213].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[212] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[213] [4:0] }), .sum({ \level_1_sums[19][106] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[215].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[214] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[215] [4:0] }), .sum({ \level_1_sums[19][107] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[215].adder_quads.adder_inst (.a({ \level_1_sums[19][107] [5:0] }),
     .b({ \level_1_sums[19][106] [5:0] }), .sum({ \level_2_sums[19][53] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[215].adder_octets.adder_inst (
    .a({ \level_2_sums[19][53] [6:0] }), .b({ \level_2_sums[19][52] [6:0] }), .sum({ \level_3_sums[19][26] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[217].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[216] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[217] [4:0] }), .sum({ \level_1_sums[19][108] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[219].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[218] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[219] [4:0] }), .sum({ \level_1_sums[19][109] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[219].adder_quads.adder_inst (.a({ \level_1_sums[19][109] [5:0] }),
     .b({ \level_1_sums[19][108] [5:0] }), .sum({ \level_2_sums[19][54] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[221].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[220] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[221] [4:0] }), .sum({ \level_1_sums[19][110] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[223].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[222] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[223] [4:0] }), .sum({ \level_1_sums[19][111] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[223].adder_quads.adder_inst (.a({ \level_1_sums[19][111] [5:0] }),
     .b({ \level_1_sums[19][110] [5:0] }), .sum({ \level_2_sums[19][55] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[223].adder_octets.adder_inst (
    .a({ \level_2_sums[19][55] [6:0] }), .b({ \level_2_sums[19][54] [6:0] }), .sum({ \level_3_sums[19][27] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[223].adder_16s.adder_inst (.a({ \level_3_sums[19][27] [7:0] }),
     .b({ \level_3_sums[19][26] [7:0] }), .sum({ \level_4_sums[19][13] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[223].adder_32s.adder_inst (.a({ \level_4_sums[19][13] [8:0] }),
     .b({ \level_4_sums[19][12] [8:0] }), .sum({ \level_5_sums[19][6] [9:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[225].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[224] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[225] [4:0] }), .sum({ \level_1_sums[19][112] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[227].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[226] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[227] [4:0] }), .sum({ \level_1_sums[19][113] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[227].adder_quads.adder_inst (.a({ \level_1_sums[19][113] [5:0] }),
     .b({ \level_1_sums[19][112] [5:0] }), .sum({ \level_2_sums[19][56] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[229].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[228] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[229] [4:0] }), .sum({ \level_1_sums[19][114] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[231].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[230] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[231] [4:0] }), .sum({ \level_1_sums[19][115] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[231].adder_quads.adder_inst (.a({ \level_1_sums[19][115] [5:0] }),
     .b({ \level_1_sums[19][114] [5:0] }), .sum({ \level_2_sums[19][57] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[231].adder_octets.adder_inst (
    .a({ \level_2_sums[19][57] [6:0] }), .b({ \level_2_sums[19][56] [6:0] }), .sum({ \level_3_sums[19][28] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[233].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[232] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[233] [4:0] }), .sum({ \level_1_sums[19][116] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[235].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[234] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[235] [4:0] }), .sum({ \level_1_sums[19][117] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[235].adder_quads.adder_inst (.a({ \level_1_sums[19][117] [5:0] }),
     .b({ \level_1_sums[19][116] [5:0] }), .sum({ \level_2_sums[19][58] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[237].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[236] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[237] [4:0] }), .sum({ \level_1_sums[19][118] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[239].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[238] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[239] [4:0] }), .sum({ \level_1_sums[19][119] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[239].adder_quads.adder_inst (.a({ \level_1_sums[19][119] [5:0] }),
     .b({ \level_1_sums[19][118] [5:0] }), .sum({ \level_2_sums[19][59] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[239].adder_octets.adder_inst (
    .a({ \level_2_sums[19][59] [6:0] }), .b({ \level_2_sums[19][58] [6:0] }), .sum({ \level_3_sums[19][29] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[239].adder_16s.adder_inst (.a({ \level_3_sums[19][29] [7:0] }),
     .b({ \level_3_sums[19][28] [7:0] }), .sum({ \level_4_sums[19][14] [8:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[241].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[240] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[241] [4:0] }), .sum({ \level_1_sums[19][120] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[243].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[242] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[243] [4:0] }), .sum({ \level_1_sums[19][121] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[243].adder_quads.adder_inst (.a({ \level_1_sums[19][121] [5:0] }),
     .b({ \level_1_sums[19][120] [5:0] }), .sum({ \level_2_sums[19][60] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[245].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[244] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[245] [4:0] }), .sum({ \level_1_sums[19][122] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[247].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[246] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[247] [4:0] }), .sum({ \level_1_sums[19][123] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[247].adder_quads.adder_inst (.a({ \level_1_sums[19][123] [5:0] }),
     .b({ \level_1_sums[19][122] [5:0] }), .sum({ \level_2_sums[19][61] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[247].adder_octets.adder_inst (
    .a({ \level_2_sums[19][61] [6:0] }), .b({ \level_2_sums[19][60] [6:0] }), .sum({ \level_3_sums[19][30] [7:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[249].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[248] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[249] [4:0] }), .sum({ \level_1_sums[19][124] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[251].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[250] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[251] [4:0] }), .sum({ \level_1_sums[19][125] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[251].adder_quads.adder_inst (.a({ \level_1_sums[19][125] [5:0] }),
     .b({ \level_1_sums[19][124] [5:0] }), .sum({ \level_2_sums[19][62] [6:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[253].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[252] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[253] [4:0] }), .sum({ \level_1_sums[19][126] [5:0] }));
  adder_5to6 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_pairs.adder_inst (.a({ \dot_product_and_ReLU[19].product_terms[254] [4:0] }),
     .b({ \dot_product_and_ReLU[19].product_terms[255] [4:0] }), .sum({ \level_1_sums[19][127] [5:0] }));
  adder_6to7 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_quads.adder_inst (.a({ \level_1_sums[19][127] [5:0] }),
     .b({ \level_1_sums[19][126] [5:0] }), .sum({ \level_2_sums[19][63] [6:0] }));
  adder_7to8 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_octets.adder_inst (
    .a({ \level_2_sums[19][63] [6:0] }), .b({ \level_2_sums[19][62] [6:0] }), .sum({ \level_3_sums[19][31] [7:0] }));
  adder_8to9 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_16s.adder_inst (.a({ \level_3_sums[19][31] [7:0] }),
     .b({ \level_3_sums[19][30] [7:0] }), .sum({ \level_4_sums[19][15] [8:0] }));
  adder_9to10 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_32s.adder_inst (.a({ \level_4_sums[19][15] [8:0] }),
     .b({ \level_4_sums[19][14] [8:0] }), .sum({ \level_5_sums[19][7] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_64s.adder_inst (.a({ \level_5_sums[19][7] [9:0] }),
     .b({ \level_5_sums[19][6] [9:0] }), .sum({ \level_6_sums[19][3] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[255].adder_128s.adder_inst (.a({ \level_6_sums[19][3] [9:0] }),
     .b({ \level_6_sums[19][2] [9:0] }), .sum({ \level_7_sums[19][1] [9:0] }));
  adder_10to10 
    \dot_product_and_ReLU[19].product_terms_gen[255].final_adder.adder_inst (.a({ \level_7_sums[19][0] [9:0] }),
     .b({ \level_7_sums[19][1] [9:0] }), .sum({ \level_8_sums[19] [9:0] }));
endmodule

module VDW_ADD_19_1_0(SUM, A, B);
input   [18:0] A;
input   [18:0] B;
output  [18:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76, N$77, N$78, N$79, N$80, N$81, N$82, N$83, N$84, N$85, N$86, 
    N$87;
wire   [18:0] SUM;
wire   [18:0] B;
wire   [18:0] A;
  xor U$1(SUM[18], N$2, N$1);
  xor U$2(N$2, A[18], B[18]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[17], N$6);
  and U$5(N$4, B[17], N$6);
  and U$6(N$5, A[17], B[17]);
  xor U$7(SUM[17], N$7, N$6);
  xor U$8(N$7, A[17], B[17]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[16], N$11);
  and U$11(N$9, B[16], N$11);
  and U$12(N$10, A[16], B[16]);
  xor U$13(SUM[16], N$12, N$11);
  xor U$14(N$12, A[16], B[16]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[15], N$16);
  and U$17(N$14, B[15], N$16);
  and U$18(N$15, A[15], B[15]);
  xor U$19(SUM[15], N$17, N$16);
  xor U$20(N$17, A[15], B[15]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[14], N$21);
  and U$23(N$19, B[14], N$21);
  and U$24(N$20, A[14], B[14]);
  xor U$25(SUM[14], N$22, N$21);
  xor U$26(N$22, A[14], B[14]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[13], N$26);
  and U$29(N$24, B[13], N$26);
  and U$30(N$25, A[13], B[13]);
  xor U$31(SUM[13], N$27, N$26);
  xor U$32(N$27, A[13], B[13]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[12], N$31);
  and U$35(N$29, B[12], N$31);
  and U$36(N$30, A[12], B[12]);
  xor U$37(SUM[12], N$32, N$31);
  xor U$38(N$32, A[12], B[12]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[11], N$36);
  and U$41(N$34, B[11], N$36);
  and U$42(N$35, A[11], B[11]);
  xor U$43(SUM[11], N$37, N$36);
  xor U$44(N$37, A[11], B[11]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[10], N$41);
  and U$47(N$39, B[10], N$41);
  and U$48(N$40, A[10], B[10]);
  xor U$49(SUM[10], N$42, N$41);
  xor U$50(N$42, A[10], B[10]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[9], N$46);
  and U$53(N$44, B[9], N$46);
  and U$54(N$45, A[9], B[9]);
  xor U$55(SUM[9], N$47, N$46);
  xor U$56(N$47, A[9], B[9]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[8], N$51);
  and U$59(N$49, B[8], N$51);
  and U$60(N$50, A[8], B[8]);
  xor U$61(SUM[8], N$52, N$51);
  xor U$62(N$52, A[8], B[8]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[7], N$56);
  and U$65(N$54, B[7], N$56);
  and U$66(N$55, A[7], B[7]);
  xor U$67(SUM[7], N$57, N$56);
  xor U$68(N$57, A[7], B[7]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[6], N$61);
  and U$71(N$59, B[6], N$61);
  and U$72(N$60, A[6], B[6]);
  xor U$73(SUM[6], N$62, N$61);
  xor U$74(N$62, A[6], B[6]);
  or U$75(N$61, N$65, N$64, N$63);
  and U$76(N$63, A[5], N$66);
  and U$77(N$64, B[5], N$66);
  and U$78(N$65, A[5], B[5]);
  xor U$79(SUM[5], N$67, N$66);
  xor U$80(N$67, A[5], B[5]);
  or U$81(N$66, N$70, N$69, N$68);
  and U$82(N$68, A[4], N$71);
  and U$83(N$69, B[4], N$71);
  and U$84(N$70, A[4], B[4]);
  xor U$85(SUM[4], N$72, N$71);
  xor U$86(N$72, A[4], B[4]);
  or U$87(N$71, N$75, N$74, N$73);
  and U$88(N$73, A[3], N$76);
  and U$89(N$74, B[3], N$76);
  and U$90(N$75, A[3], B[3]);
  xor U$91(SUM[3], N$77, N$76);
  xor U$92(N$77, A[3], B[3]);
  or U$93(N$76, N$80, N$79, N$78);
  and U$94(N$78, A[2], N$81);
  and U$95(N$79, B[2], N$81);
  and U$96(N$80, A[2], B[2]);
  xor U$97(SUM[2], N$82, N$81);
  xor U$98(N$82, A[2], B[2]);
  or U$99(N$81, N$85, N$84, N$83);
  and U$100(N$83, A[1], N$86);
  and U$101(N$84, B[1], N$86);
  and U$102(N$85, A[1], B[1]);
  xor U$103(SUM[1], N$87, N$86);
  xor U$104(N$87, A[1], B[1]);
  and U$105(N$86, A[0], B[0]);
  xor U$106(SUM[0], A[0], B[0]);
endmodule

module VDW_ADD_18_1_0(SUM, A, B);
input   [17:0] A;
input   [17:0] B;
output  [17:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76, N$77, N$78, N$79, N$80, N$81, N$82;
wire   [17:0] SUM;
wire   [17:0] B;
wire   [17:0] A;
  xor U$1(SUM[17], N$2, N$1);
  xor U$2(N$2, A[17], B[17]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[16], N$6);
  and U$5(N$4, B[16], N$6);
  and U$6(N$5, A[16], B[16]);
  xor U$7(SUM[16], N$7, N$6);
  xor U$8(N$7, A[16], B[16]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[15], N$11);
  and U$11(N$9, B[15], N$11);
  and U$12(N$10, A[15], B[15]);
  xor U$13(SUM[15], N$12, N$11);
  xor U$14(N$12, A[15], B[15]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[14], N$16);
  and U$17(N$14, B[14], N$16);
  and U$18(N$15, A[14], B[14]);
  xor U$19(SUM[14], N$17, N$16);
  xor U$20(N$17, A[14], B[14]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[13], N$21);
  and U$23(N$19, B[13], N$21);
  and U$24(N$20, A[13], B[13]);
  xor U$25(SUM[13], N$22, N$21);
  xor U$26(N$22, A[13], B[13]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[12], N$26);
  and U$29(N$24, B[12], N$26);
  and U$30(N$25, A[12], B[12]);
  xor U$31(SUM[12], N$27, N$26);
  xor U$32(N$27, A[12], B[12]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[11], N$31);
  and U$35(N$29, B[11], N$31);
  and U$36(N$30, A[11], B[11]);
  xor U$37(SUM[11], N$32, N$31);
  xor U$38(N$32, A[11], B[11]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[10], N$36);
  and U$41(N$34, B[10], N$36);
  and U$42(N$35, A[10], B[10]);
  xor U$43(SUM[10], N$37, N$36);
  xor U$44(N$37, A[10], B[10]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[9], N$41);
  and U$47(N$39, B[9], N$41);
  and U$48(N$40, A[9], B[9]);
  xor U$49(SUM[9], N$42, N$41);
  xor U$50(N$42, A[9], B[9]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[8], N$46);
  and U$53(N$44, B[8], N$46);
  and U$54(N$45, A[8], B[8]);
  xor U$55(SUM[8], N$47, N$46);
  xor U$56(N$47, A[8], B[8]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[7], N$51);
  and U$59(N$49, B[7], N$51);
  and U$60(N$50, A[7], B[7]);
  xor U$61(SUM[7], N$52, N$51);
  xor U$62(N$52, A[7], B[7]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[6], N$56);
  and U$65(N$54, B[6], N$56);
  and U$66(N$55, A[6], B[6]);
  xor U$67(SUM[6], N$57, N$56);
  xor U$68(N$57, A[6], B[6]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[5], N$61);
  and U$71(N$59, B[5], N$61);
  and U$72(N$60, A[5], B[5]);
  xor U$73(SUM[5], N$62, N$61);
  xor U$74(N$62, A[5], B[5]);
  or U$75(N$61, N$65, N$64, N$63);
  and U$76(N$63, A[4], N$66);
  and U$77(N$64, B[4], N$66);
  and U$78(N$65, A[4], B[4]);
  xor U$79(SUM[4], N$67, N$66);
  xor U$80(N$67, A[4], B[4]);
  or U$81(N$66, N$70, N$69, N$68);
  and U$82(N$68, A[3], N$71);
  and U$83(N$69, B[3], N$71);
  and U$84(N$70, A[3], B[3]);
  xor U$85(SUM[3], N$72, N$71);
  xor U$86(N$72, A[3], B[3]);
  or U$87(N$71, N$75, N$74, N$73);
  and U$88(N$73, A[2], N$76);
  and U$89(N$74, B[2], N$76);
  and U$90(N$75, A[2], B[2]);
  xor U$91(SUM[2], N$77, N$76);
  xor U$92(N$77, A[2], B[2]);
  or U$93(N$76, N$80, N$79, N$78);
  and U$94(N$78, A[1], N$81);
  and U$95(N$79, B[1], N$81);
  and U$96(N$80, A[1], B[1]);
  xor U$97(SUM[1], N$82, N$81);
  xor U$98(N$82, A[1], B[1]);
  and U$99(N$81, A[0], B[0]);
  xor U$100(SUM[0], A[0], B[0]);
endmodule

module VDW_ADD_17_1_0(SUM, A, B);
input   [16:0] A;
input   [16:0] B;
output  [16:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76, N$77;
wire   [16:0] SUM;
wire   [16:0] B;
wire   [16:0] A;
  xor U$1(SUM[16], N$2, N$1);
  xor U$2(N$2, A[16], B[16]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[15], N$6);
  and U$5(N$4, B[15], N$6);
  and U$6(N$5, A[15], B[15]);
  xor U$7(SUM[15], N$7, N$6);
  xor U$8(N$7, A[15], B[15]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[14], N$11);
  and U$11(N$9, B[14], N$11);
  and U$12(N$10, A[14], B[14]);
  xor U$13(SUM[14], N$12, N$11);
  xor U$14(N$12, A[14], B[14]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[13], N$16);
  and U$17(N$14, B[13], N$16);
  and U$18(N$15, A[13], B[13]);
  xor U$19(SUM[13], N$17, N$16);
  xor U$20(N$17, A[13], B[13]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[12], N$21);
  and U$23(N$19, B[12], N$21);
  and U$24(N$20, A[12], B[12]);
  xor U$25(SUM[12], N$22, N$21);
  xor U$26(N$22, A[12], B[12]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[11], N$26);
  and U$29(N$24, B[11], N$26);
  and U$30(N$25, A[11], B[11]);
  xor U$31(SUM[11], N$27, N$26);
  xor U$32(N$27, A[11], B[11]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[10], N$31);
  and U$35(N$29, B[10], N$31);
  and U$36(N$30, A[10], B[10]);
  xor U$37(SUM[10], N$32, N$31);
  xor U$38(N$32, A[10], B[10]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[9], N$36);
  and U$41(N$34, B[9], N$36);
  and U$42(N$35, A[9], B[9]);
  xor U$43(SUM[9], N$37, N$36);
  xor U$44(N$37, A[9], B[9]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[8], N$41);
  and U$47(N$39, B[8], N$41);
  and U$48(N$40, A[8], B[8]);
  xor U$49(SUM[8], N$42, N$41);
  xor U$50(N$42, A[8], B[8]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[7], N$46);
  and U$53(N$44, B[7], N$46);
  and U$54(N$45, A[7], B[7]);
  xor U$55(SUM[7], N$47, N$46);
  xor U$56(N$47, A[7], B[7]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[6], N$51);
  and U$59(N$49, B[6], N$51);
  and U$60(N$50, A[6], B[6]);
  xor U$61(SUM[6], N$52, N$51);
  xor U$62(N$52, A[6], B[6]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[5], N$56);
  and U$65(N$54, B[5], N$56);
  and U$66(N$55, A[5], B[5]);
  xor U$67(SUM[5], N$57, N$56);
  xor U$68(N$57, A[5], B[5]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[4], N$61);
  and U$71(N$59, B[4], N$61);
  and U$72(N$60, A[4], B[4]);
  xor U$73(SUM[4], N$62, N$61);
  xor U$74(N$62, A[4], B[4]);
  or U$75(N$61, N$65, N$64, N$63);
  and U$76(N$63, A[3], N$66);
  and U$77(N$64, B[3], N$66);
  and U$78(N$65, A[3], B[3]);
  xor U$79(SUM[3], N$67, N$66);
  xor U$80(N$67, A[3], B[3]);
  or U$81(N$66, N$70, N$69, N$68);
  and U$82(N$68, A[2], N$71);
  and U$83(N$69, B[2], N$71);
  and U$84(N$70, A[2], B[2]);
  xor U$85(SUM[2], N$72, N$71);
  xor U$86(N$72, A[2], B[2]);
  or U$87(N$71, N$75, N$74, N$73);
  and U$88(N$73, A[1], N$76);
  and U$89(N$74, B[1], N$76);
  and U$90(N$75, A[1], B[1]);
  xor U$91(SUM[1], N$77, N$76);
  xor U$92(N$77, A[1], B[1]);
  and U$93(N$76, A[0], B[0]);
  xor U$94(SUM[0], A[0], B[0]);
endmodule

module VDW_ADD_16_1_0(SUM, A, B);
input   [15:0] A;
input   [15:0] B;
output  [15:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72;
wire   [15:0] SUM;
wire   [15:0] B;
wire   [15:0] A;
  xor U$1(SUM[15], N$2, N$1);
  xor U$2(N$2, A[15], B[15]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[14], N$6);
  and U$5(N$4, B[14], N$6);
  and U$6(N$5, A[14], B[14]);
  xor U$7(SUM[14], N$7, N$6);
  xor U$8(N$7, A[14], B[14]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[13], N$11);
  and U$11(N$9, B[13], N$11);
  and U$12(N$10, A[13], B[13]);
  xor U$13(SUM[13], N$12, N$11);
  xor U$14(N$12, A[13], B[13]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[12], N$16);
  and U$17(N$14, B[12], N$16);
  and U$18(N$15, A[12], B[12]);
  xor U$19(SUM[12], N$17, N$16);
  xor U$20(N$17, A[12], B[12]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[11], N$21);
  and U$23(N$19, B[11], N$21);
  and U$24(N$20, A[11], B[11]);
  xor U$25(SUM[11], N$22, N$21);
  xor U$26(N$22, A[11], B[11]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[10], N$26);
  and U$29(N$24, B[10], N$26);
  and U$30(N$25, A[10], B[10]);
  xor U$31(SUM[10], N$27, N$26);
  xor U$32(N$27, A[10], B[10]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[9], N$31);
  and U$35(N$29, B[9], N$31);
  and U$36(N$30, A[9], B[9]);
  xor U$37(SUM[9], N$32, N$31);
  xor U$38(N$32, A[9], B[9]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[8], N$36);
  and U$41(N$34, B[8], N$36);
  and U$42(N$35, A[8], B[8]);
  xor U$43(SUM[8], N$37, N$36);
  xor U$44(N$37, A[8], B[8]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[7], N$41);
  and U$47(N$39, B[7], N$41);
  and U$48(N$40, A[7], B[7]);
  xor U$49(SUM[7], N$42, N$41);
  xor U$50(N$42, A[7], B[7]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[6], N$46);
  and U$53(N$44, B[6], N$46);
  and U$54(N$45, A[6], B[6]);
  xor U$55(SUM[6], N$47, N$46);
  xor U$56(N$47, A[6], B[6]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[5], N$51);
  and U$59(N$49, B[5], N$51);
  and U$60(N$50, A[5], B[5]);
  xor U$61(SUM[5], N$52, N$51);
  xor U$62(N$52, A[5], B[5]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[4], N$56);
  and U$65(N$54, B[4], N$56);
  and U$66(N$55, A[4], B[4]);
  xor U$67(SUM[4], N$57, N$56);
  xor U$68(N$57, A[4], B[4]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[3], N$61);
  and U$71(N$59, B[3], N$61);
  and U$72(N$60, A[3], B[3]);
  xor U$73(SUM[3], N$62, N$61);
  xor U$74(N$62, A[3], B[3]);
  or U$75(N$61, N$65, N$64, N$63);
  and U$76(N$63, A[2], N$66);
  and U$77(N$64, B[2], N$66);
  and U$78(N$65, A[2], B[2]);
  xor U$79(SUM[2], N$67, N$66);
  xor U$80(N$67, A[2], B[2]);
  or U$81(N$66, N$70, N$69, N$68);
  and U$82(N$68, A[1], N$71);
  and U$83(N$69, B[1], N$71);
  and U$84(N$70, A[1], B[1]);
  xor U$85(SUM[1], N$72, N$71);
  xor U$86(N$72, A[1], B[1]);
  and U$87(N$71, A[0], B[0]);
  xor U$88(SUM[0], A[0], B[0]);
endmodule

module VDW_ADD_15_1_0(SUM, A, B);
input   [14:0] A;
input   [14:0] B;
output  [14:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67;
wire   [14:0] SUM;
wire   [14:0] B;
wire   [14:0] A;
  xor U$1(SUM[14], N$2, N$1);
  xor U$2(N$2, A[14], B[14]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[13], N$6);
  and U$5(N$4, B[13], N$6);
  and U$6(N$5, A[13], B[13]);
  xor U$7(SUM[13], N$7, N$6);
  xor U$8(N$7, A[13], B[13]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[12], N$11);
  and U$11(N$9, B[12], N$11);
  and U$12(N$10, A[12], B[12]);
  xor U$13(SUM[12], N$12, N$11);
  xor U$14(N$12, A[12], B[12]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[11], N$16);
  and U$17(N$14, B[11], N$16);
  and U$18(N$15, A[11], B[11]);
  xor U$19(SUM[11], N$17, N$16);
  xor U$20(N$17, A[11], B[11]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[10], N$21);
  and U$23(N$19, B[10], N$21);
  and U$24(N$20, A[10], B[10]);
  xor U$25(SUM[10], N$22, N$21);
  xor U$26(N$22, A[10], B[10]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[9], N$26);
  and U$29(N$24, B[9], N$26);
  and U$30(N$25, A[9], B[9]);
  xor U$31(SUM[9], N$27, N$26);
  xor U$32(N$27, A[9], B[9]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[8], N$31);
  and U$35(N$29, B[8], N$31);
  and U$36(N$30, A[8], B[8]);
  xor U$37(SUM[8], N$32, N$31);
  xor U$38(N$32, A[8], B[8]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[7], N$36);
  and U$41(N$34, B[7], N$36);
  and U$42(N$35, A[7], B[7]);
  xor U$43(SUM[7], N$37, N$36);
  xor U$44(N$37, A[7], B[7]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[6], N$41);
  and U$47(N$39, B[6], N$41);
  and U$48(N$40, A[6], B[6]);
  xor U$49(SUM[6], N$42, N$41);
  xor U$50(N$42, A[6], B[6]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[5], N$46);
  and U$53(N$44, B[5], N$46);
  and U$54(N$45, A[5], B[5]);
  xor U$55(SUM[5], N$47, N$46);
  xor U$56(N$47, A[5], B[5]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[4], N$51);
  and U$59(N$49, B[4], N$51);
  and U$60(N$50, A[4], B[4]);
  xor U$61(SUM[4], N$52, N$51);
  xor U$62(N$52, A[4], B[4]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[3], N$56);
  and U$65(N$54, B[3], N$56);
  and U$66(N$55, A[3], B[3]);
  xor U$67(SUM[3], N$57, N$56);
  xor U$68(N$57, A[3], B[3]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[2], N$61);
  and U$71(N$59, B[2], N$61);
  and U$72(N$60, A[2], B[2]);
  xor U$73(SUM[2], N$62, N$61);
  xor U$74(N$62, A[2], B[2]);
  or U$75(N$61, N$65, N$64, N$63);
  and U$76(N$63, A[1], N$66);
  and U$77(N$64, B[1], N$66);
  and U$78(N$65, A[1], B[1]);
  xor U$79(SUM[1], N$67, N$66);
  xor U$80(N$67, A[1], B[1]);
  and U$81(N$66, A[0], B[0]);
  xor U$82(SUM[0], A[0], B[0]);
endmodule

module VDW_WMUX18 (Z, A, B, S);
// conformal library_module
output [17:0] Z;
input [17:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module ReLU_19bit(in_data, out_data);
input   [18:0] in_data;
output  [17:0] out_data;
wire  n207;
wire   [17:0] out_data;
wire   [18:0] in_data;
  VDW_WMUX18 U$1(.Z({ out_data[17:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
    1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({ in_data[17:0] }), .S(n207));
  not U$2(n207, in_data[18]);
endmodule

module VDW_ADD_14_1_0(SUM, A, B);
input   [13:0] A;
input   [13:0] B;
output  [13:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62;
wire   [13:0] SUM;
wire   [13:0] B;
wire   [13:0] A;
  xor U$1(SUM[13], N$2, N$1);
  xor U$2(N$2, A[13], B[13]);
  or U$3(N$1, N$5, N$4, N$3);
  and U$4(N$3, A[12], N$6);
  and U$5(N$4, B[12], N$6);
  and U$6(N$5, A[12], B[12]);
  xor U$7(SUM[12], N$7, N$6);
  xor U$8(N$7, A[12], B[12]);
  or U$9(N$6, N$10, N$9, N$8);
  and U$10(N$8, A[11], N$11);
  and U$11(N$9, B[11], N$11);
  and U$12(N$10, A[11], B[11]);
  xor U$13(SUM[11], N$12, N$11);
  xor U$14(N$12, A[11], B[11]);
  or U$15(N$11, N$15, N$14, N$13);
  and U$16(N$13, A[10], N$16);
  and U$17(N$14, B[10], N$16);
  and U$18(N$15, A[10], B[10]);
  xor U$19(SUM[10], N$17, N$16);
  xor U$20(N$17, A[10], B[10]);
  or U$21(N$16, N$20, N$19, N$18);
  and U$22(N$18, A[9], N$21);
  and U$23(N$19, B[9], N$21);
  and U$24(N$20, A[9], B[9]);
  xor U$25(SUM[9], N$22, N$21);
  xor U$26(N$22, A[9], B[9]);
  or U$27(N$21, N$25, N$24, N$23);
  and U$28(N$23, A[8], N$26);
  and U$29(N$24, B[8], N$26);
  and U$30(N$25, A[8], B[8]);
  xor U$31(SUM[8], N$27, N$26);
  xor U$32(N$27, A[8], B[8]);
  or U$33(N$26, N$30, N$29, N$28);
  and U$34(N$28, A[7], N$31);
  and U$35(N$29, B[7], N$31);
  and U$36(N$30, A[7], B[7]);
  xor U$37(SUM[7], N$32, N$31);
  xor U$38(N$32, A[7], B[7]);
  or U$39(N$31, N$35, N$34, N$33);
  and U$40(N$33, A[6], N$36);
  and U$41(N$34, B[6], N$36);
  and U$42(N$35, A[6], B[6]);
  xor U$43(SUM[6], N$37, N$36);
  xor U$44(N$37, A[6], B[6]);
  or U$45(N$36, N$40, N$39, N$38);
  and U$46(N$38, A[5], N$41);
  and U$47(N$39, B[5], N$41);
  and U$48(N$40, A[5], B[5]);
  xor U$49(SUM[5], N$42, N$41);
  xor U$50(N$42, A[5], B[5]);
  or U$51(N$41, N$45, N$44, N$43);
  and U$52(N$43, A[4], N$46);
  and U$53(N$44, B[4], N$46);
  and U$54(N$45, A[4], B[4]);
  xor U$55(SUM[4], N$47, N$46);
  xor U$56(N$47, A[4], B[4]);
  or U$57(N$46, N$50, N$49, N$48);
  and U$58(N$48, A[3], N$51);
  and U$59(N$49, B[3], N$51);
  and U$60(N$50, A[3], B[3]);
  xor U$61(SUM[3], N$52, N$51);
  xor U$62(N$52, A[3], B[3]);
  or U$63(N$51, N$55, N$54, N$53);
  and U$64(N$53, A[2], N$56);
  and U$65(N$54, B[2], N$56);
  and U$66(N$55, A[2], B[2]);
  xor U$67(SUM[2], N$57, N$56);
  xor U$68(N$57, A[2], B[2]);
  or U$69(N$56, N$60, N$59, N$58);
  and U$70(N$58, A[1], N$61);
  and U$71(N$59, B[1], N$61);
  and U$72(N$60, A[1], B[1]);
  xor U$73(SUM[1], N$62, N$61);
  xor U$74(N$62, A[1], B[1]);
  and U$75(N$61, A[0], B[0]);
  xor U$76(SUM[0], A[0], B[0]);
endmodule

module VDW_SUB_14_1_0(SUM, A, B);
input   [13:0] A;
input   [13:0] B;
output  [13:0] SUM;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76;
wire   [13:0] SUM;
wire   [13:0] B;
wire   [13:0] A;
  xor U$1(SUM[13], N$2, N$1);
  xor U$2(N$2, A[13], N$3);
  not U$3(N$3, B[13]);
  or U$4(N$1, N$6, N$5, N$4);
  and U$5(N$4, A[12], N$7);
  and U$6(N$5, N$9, N$7);
  and U$7(N$6, A[12], N$9);
  xor U$8(SUM[12], N$8, N$7);
  xor U$9(N$8, A[12], N$9);
  not U$10(N$9, B[12]);
  or U$11(N$7, N$12, N$11, N$10);
  and U$12(N$10, A[11], N$13);
  and U$13(N$11, N$15, N$13);
  and U$14(N$12, A[11], N$15);
  xor U$15(SUM[11], N$14, N$13);
  xor U$16(N$14, A[11], N$15);
  not U$17(N$15, B[11]);
  or U$18(N$13, N$18, N$17, N$16);
  and U$19(N$16, A[10], N$19);
  and U$20(N$17, N$21, N$19);
  and U$21(N$18, A[10], N$21);
  xor U$22(SUM[10], N$20, N$19);
  xor U$23(N$20, A[10], N$21);
  not U$24(N$21, B[10]);
  or U$25(N$19, N$24, N$23, N$22);
  and U$26(N$22, A[9], N$25);
  and U$27(N$23, N$27, N$25);
  and U$28(N$24, A[9], N$27);
  xor U$29(SUM[9], N$26, N$25);
  xor U$30(N$26, A[9], N$27);
  not U$31(N$27, B[9]);
  or U$32(N$25, N$30, N$29, N$28);
  and U$33(N$28, A[8], N$31);
  and U$34(N$29, N$33, N$31);
  and U$35(N$30, A[8], N$33);
  xor U$36(SUM[8], N$32, N$31);
  xor U$37(N$32, A[8], N$33);
  not U$38(N$33, B[8]);
  or U$39(N$31, N$36, N$35, N$34);
  and U$40(N$34, A[7], N$37);
  and U$41(N$35, N$39, N$37);
  and U$42(N$36, A[7], N$39);
  xor U$43(SUM[7], N$38, N$37);
  xor U$44(N$38, A[7], N$39);
  not U$45(N$39, B[7]);
  or U$46(N$37, N$42, N$41, N$40);
  and U$47(N$40, A[6], N$43);
  and U$48(N$41, N$45, N$43);
  and U$49(N$42, A[6], N$45);
  xor U$50(SUM[6], N$44, N$43);
  xor U$51(N$44, A[6], N$45);
  not U$52(N$45, B[6]);
  or U$53(N$43, N$48, N$47, N$46);
  and U$54(N$46, A[5], N$49);
  and U$55(N$47, N$51, N$49);
  and U$56(N$48, A[5], N$51);
  xor U$57(SUM[5], N$50, N$49);
  xor U$58(N$50, A[5], N$51);
  not U$59(N$51, B[5]);
  or U$60(N$49, N$54, N$53, N$52);
  and U$61(N$52, A[4], N$55);
  and U$62(N$53, N$57, N$55);
  and U$63(N$54, A[4], N$57);
  xor U$64(SUM[4], N$56, N$55);
  xor U$65(N$56, A[4], N$57);
  not U$66(N$57, B[4]);
  or U$67(N$55, N$60, N$59, N$58);
  and U$68(N$58, A[3], N$61);
  and U$69(N$59, N$63, N$61);
  and U$70(N$60, A[3], N$63);
  xor U$71(SUM[3], N$62, N$61);
  xor U$72(N$62, A[3], N$63);
  not U$73(N$63, B[3]);
  or U$74(N$61, N$66, N$65, N$64);
  and U$75(N$64, A[2], N$67);
  and U$76(N$65, N$69, N$67);
  and U$77(N$66, A[2], N$69);
  xor U$78(SUM[2], N$68, N$67);
  xor U$79(N$68, A[2], N$69);
  not U$80(N$69, B[2]);
  or U$81(N$67, N$72, N$71, N$70);
  and U$82(N$70, A[1], N$73);
  and U$83(N$71, N$75, N$73);
  and U$84(N$72, A[1], N$75);
  xor U$85(SUM[1], N$74, N$73);
  xor U$86(N$74, A[1], N$75);
  not U$87(N$75, B[1]);
  or U$88(N$73, A[0], N$76);
  xor U$89(SUM[0], A[0], B[0]);
  not U$90(N$76, B[0]);
endmodule

module multiplier9514(prod, num1, num2);
input   [8:0] num1;
input   [4:0] num2;
output  [13:0] prod;
wire   [13:0] \intermediate_sums[0] ;
wire   [13:0] \intermediate_sums[1] ;
wire   [13:0] \intermediate_sums[2] ;
wire   [13:0] \shifted_pps[0] ;
wire   [13:0] \shifted_pps[1] ;
wire   [13:0] \shifted_pps[2] ;
wire   [13:0] \shifted_pps[3] ;
wire   [13:0] \shifted_pps[4] ;
wire   [8:0] \partial_prods[0] ;
wire   [8:0] \partial_prods[1] ;
wire   [8:0] \partial_prods[2] ;
wire   [8:0] \partial_prods[3] ;
wire   [8:0] \partial_prods[4] ;
wire   [4:0] num2;
wire   [8:0] num1;
wire   [13:0] prod;
  assign \shifted_pps[0] [13] = 1'b0;
  assign \shifted_pps[0] [12] = 1'b0;
  assign \shifted_pps[0] [11] = 1'b0;
  assign \shifted_pps[0] [10] = 1'b0;
  assign \shifted_pps[0] [9] = 1'b0;
  assign \shifted_pps[1] [13] = 1'b0;
  assign \shifted_pps[1] [12] = 1'b0;
  assign \shifted_pps[1] [11] = 1'b0;
  assign \shifted_pps[1] [10] = 1'b0;
  assign \shifted_pps[1] [0] = 1'b0;
  assign \shifted_pps[2] [13] = 1'b0;
  assign \shifted_pps[2] [12] = 1'b0;
  assign \shifted_pps[2] [11] = 1'b0;
  assign \shifted_pps[2] [1] = 1'b0;
  assign \shifted_pps[2] [0] = 1'b0;
  assign \shifted_pps[3] [13] = 1'b0;
  assign \shifted_pps[3] [12] = 1'b0;
  assign \shifted_pps[3] [2] = 1'b0;
  assign \shifted_pps[3] [1] = 1'b0;
  assign \shifted_pps[3] [0] = 1'b0;
  assign \shifted_pps[4] [13] = 1'b0;
  assign \shifted_pps[4] [3] = 1'b0;
  assign \shifted_pps[4] [2] = 1'b0;
  assign \shifted_pps[4] [1] = 1'b0;
  assign \shifted_pps[4] [0] = 1'b0;
  VDW_ADD_14_1_0 add_183_50(.SUM({ \intermediate_sums[0] [13:0] }), .A({ \shifted_pps[0] [13:0] }), .B({ \shifted_pps[1] [13:0] }));
  VDW_ADD_14_1_0 add_184_56(.SUM({ \intermediate_sums[1] [13:0] }), .A({ \intermediate_sums[0] [13:0] }), .B({ \shifted_pps[2] [13:0] }));
  VDW_ADD_14_1_0 add_185_56(.SUM({ \intermediate_sums[2] [13:0] }), .A({ \intermediate_sums[1] [13:0] }), .B({ \shifted_pps[3] [13:0] }));
  assign \shifted_pps[0] [8] = \partial_prods[0] [8];
  assign \shifted_pps[0] [7] = \partial_prods[0] [7];
  assign \shifted_pps[0] [6] = \partial_prods[0] [6];
  assign \shifted_pps[0] [5] = \partial_prods[0] [5];
  assign \shifted_pps[0] [4] = \partial_prods[0] [4];
  assign \shifted_pps[0] [3] = \partial_prods[0] [3];
  assign \shifted_pps[0] [2] = \partial_prods[0] [2];
  assign \shifted_pps[0] [1] = \partial_prods[0] [1];
  assign \shifted_pps[0] [0] = \partial_prods[0] [0];
  assign \shifted_pps[1] [9] = \partial_prods[1] [8];
  assign \shifted_pps[1] [8] = \partial_prods[1] [7];
  assign \shifted_pps[1] [7] = \partial_prods[1] [6];
  assign \shifted_pps[1] [6] = \partial_prods[1] [5];
  assign \shifted_pps[1] [5] = \partial_prods[1] [4];
  assign \shifted_pps[1] [4] = \partial_prods[1] [3];
  assign \shifted_pps[1] [3] = \partial_prods[1] [2];
  assign \shifted_pps[1] [2] = \partial_prods[1] [1];
  assign \shifted_pps[1] [1] = \partial_prods[1] [0];
  assign \shifted_pps[2] [10] = \partial_prods[2] [8];
  assign \shifted_pps[2] [9] = \partial_prods[2] [7];
  assign \shifted_pps[2] [8] = \partial_prods[2] [6];
  assign \shifted_pps[2] [7] = \partial_prods[2] [5];
  assign \shifted_pps[2] [6] = \partial_prods[2] [4];
  assign \shifted_pps[2] [5] = \partial_prods[2] [3];
  assign \shifted_pps[2] [4] = \partial_prods[2] [2];
  assign \shifted_pps[2] [3] = \partial_prods[2] [1];
  assign \shifted_pps[2] [2] = \partial_prods[2] [0];
  assign \shifted_pps[3] [11] = \partial_prods[3] [8];
  assign \shifted_pps[3] [10] = \partial_prods[3] [7];
  assign \shifted_pps[3] [9] = \partial_prods[3] [6];
  assign \shifted_pps[3] [8] = \partial_prods[3] [5];
  assign \shifted_pps[3] [7] = \partial_prods[3] [4];
  assign \shifted_pps[3] [6] = \partial_prods[3] [3];
  assign \shifted_pps[3] [5] = \partial_prods[3] [2];
  assign \shifted_pps[3] [4] = \partial_prods[3] [1];
  assign \shifted_pps[3] [3] = \partial_prods[3] [0];
  assign \shifted_pps[4] [12] = \partial_prods[4] [8];
  assign \shifted_pps[4] [11] = \partial_prods[4] [7];
  assign \shifted_pps[4] [10] = \partial_prods[4] [6];
  assign \shifted_pps[4] [9] = \partial_prods[4] [5];
  assign \shifted_pps[4] [8] = \partial_prods[4] [4];
  assign \shifted_pps[4] [7] = \partial_prods[4] [3];
  assign \shifted_pps[4] [6] = \partial_prods[4] [2];
  assign \shifted_pps[4] [5] = \partial_prods[4] [1];
  assign \shifted_pps[4] [4] = \partial_prods[4] [0];
  VDW_WMUX9 U$46(.Z({ \partial_prods[0] [8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ num1[8:0] }), .S(num2[0]));
  VDW_WMUX9 U$47(.Z({ \partial_prods[1] [8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ num1[8:0] }), .S(num2[1]));
  VDW_WMUX9 U$48(.Z({ \partial_prods[2] [8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ num1[8:0] }), .S(num2[2]));
  VDW_WMUX9 U$49(.Z({ \partial_prods[3] [8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ num1[8:0] }), .S(num2[3]));
  VDW_WMUX9 U$50(.Z({ \partial_prods[4] [8:0] }), .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
     .B({ num1[8:0] }), .S(num2[4]));
  VDW_SUB_14_1_0 sub_186_40(.SUM({ prod[13:0] }), .A({ \intermediate_sums[2] [13:0] }), .B({ \shifted_pps[4] [13:0] }));
endmodule

module layer2(clk, rst_n, in, out);
input  clk, rst_n;
input   [179:0] in;
output  [179:0] out;
wire  n5835, rst_n, clk;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18;
wire   [18:0] n5823_19;
wire   [18:0] n5822_30;
wire   [18:0] n5822_29;
wire   [18:0] n5822_28;
wire   [18:0] n5821_30;
wire   [18:0] n5821_29;
wire   [18:0] n5821_28;
wire   [18:0] n5820_30;
wire   [18:0] n5820_29;
wire   [18:0] n5820_28;
wire   [18:0] n5819_30;
wire   [18:0] n5819_29;
wire   [18:0] n5819_28;
wire   [18:0] n5818_30;
wire   [18:0] n5818_29;
wire   [17:0] n5818_28;
wire   [16:0] n5817_30;
wire   [15:0] n5817_29;
wire   [14:0] n5817_28;
wire   [18:0] n5823_17;
wire   [18:0] n5822_27;
wire   [18:0] n5822_26;
wire   [18:0] n5822_25;
wire   [18:0] n5821_27;
wire   [18:0] n5821_26;
wire   [18:0] n5821_25;
wire   [18:0] n5820_27;
wire   [18:0] n5820_26;
wire   [18:0] n5820_25;
wire   [18:0] n5819_27;
wire   [18:0] n5819_26;
wire   [18:0] n5819_25;
wire   [18:0] n5818_27;
wire   [18:0] n5818_26;
wire   [17:0] n5818_25;
wire   [16:0] n5817_27;
wire   [15:0] n5817_26;
wire   [14:0] n5817_25;
wire   [18:0] n5823_15;
wire   [18:0] n5822_24;
wire   [18:0] n5822_23;
wire   [18:0] n5822_22;
wire   [18:0] n5821_24;
wire   [18:0] n5821_23;
wire   [18:0] n5821_22;
wire   [18:0] n5820_24;
wire   [18:0] n5820_23;
wire   [18:0] n5820_22;
wire   [18:0] n5819_24;
wire   [18:0] n5819_23;
wire   [18:0] n5819_22;
wire   [18:0] n5818_24;
wire   [18:0] n5818_23;
wire   [17:0] n5818_22;
wire   [16:0] n5817_24;
wire   [15:0] n5817_23;
wire   [14:0] n5817_22;
wire   [18:0] n5823_13;
wire   [18:0] n5822_21;
wire   [18:0] n5822_20;
wire   [18:0] n5822_19;
wire   [18:0] n5821_21;
wire   [18:0] n5821_20;
wire   [18:0] n5821_19;
wire   [18:0] n5820_21;
wire   [18:0] n5820_20;
wire   [18:0] n5820_19;
wire   [18:0] n5819_21;
wire   [18:0] n5819_20;
wire   [18:0] n5819_19;
wire   [18:0] n5818_21;
wire   [18:0] n5818_20;
wire   [17:0] n5818_19;
wire   [16:0] n5817_21;
wire   [15:0] n5817_20;
wire   [14:0] n5817_19;
wire   [18:0] n5823_11;
wire   [18:0] n5822_18;
wire   [18:0] n5822_17;
wire   [18:0] n5822_16;
wire   [18:0] n5821_18;
wire   [18:0] n5821_17;
wire   [18:0] n5821_16;
wire   [18:0] n5820_18;
wire   [18:0] n5820_17;
wire   [18:0] n5820_16;
wire   [18:0] n5819_18;
wire   [18:0] n5819_17;
wire   [18:0] n5819_16;
wire   [18:0] n5818_18;
wire   [18:0] n5818_17;
wire   [17:0] n5818_16;
wire   [16:0] n5817_18;
wire   [15:0] n5817_17;
wire   [14:0] n5817_16;
wire   [18:0] n5823_9;
wire   [18:0] n5822_15;
wire   [18:0] n5822_14;
wire   [18:0] n5822_13;
wire   [18:0] n5821_15;
wire   [18:0] n5821_14;
wire   [18:0] n5821_13;
wire   [18:0] n5820_15;
wire   [18:0] n5820_14;
wire   [18:0] n5820_13;
wire   [18:0] n5819_15;
wire   [18:0] n5819_14;
wire   [18:0] n5819_13;
wire   [18:0] n5818_15;
wire   [18:0] n5818_14;
wire   [17:0] n5818_13;
wire   [16:0] n5817_15;
wire   [15:0] n5817_14;
wire   [14:0] n5817_13;
wire   [18:0] n5823_7;
wire   [18:0] n5822_12;
wire   [18:0] n5822_11;
wire   [18:0] n5822_10;
wire   [18:0] n5821_12;
wire   [18:0] n5821_11;
wire   [18:0] n5821_10;
wire   [18:0] n5820_12;
wire   [18:0] n5820_11;
wire   [18:0] n5820_10;
wire   [18:0] n5819_12;
wire   [18:0] n5819_11;
wire   [18:0] n5819_10;
wire   [18:0] n5818_12;
wire   [18:0] n5818_11;
wire   [17:0] n5818_10;
wire   [16:0] n5817_12;
wire   [15:0] n5817_11;
wire   [14:0] n5817_10;
wire   [18:0] n5823_5;
wire   [18:0] n5822_9;
wire   [18:0] n5822_8;
wire   [18:0] n5822_7;
wire   [18:0] n5821_9;
wire   [18:0] n5821_8;
wire   [18:0] n5821_7;
wire   [18:0] n5820_9;
wire   [18:0] n5820_8;
wire   [18:0] n5820_7;
wire   [18:0] n5819_9;
wire   [18:0] n5819_8;
wire   [18:0] n5819_7;
wire   [18:0] n5818_9;
wire   [18:0] n5818_8;
wire   [17:0] n5818_7;
wire   [16:0] n5817_9;
wire   [15:0] n5817_8;
wire   [14:0] n5817_7;
wire   [18:0] n5823_3;
wire   [18:0] n5822_6;
wire   [18:0] n5822_5;
wire   [18:0] n5822_4;
wire   [18:0] n5821_6;
wire   [18:0] n5821_5;
wire   [18:0] n5821_4;
wire   [18:0] n5820_6;
wire   [18:0] n5820_5;
wire   [18:0] n5820_4;
wire   [18:0] n5819_6;
wire   [18:0] n5819_5;
wire   [18:0] n5819_4;
wire   [18:0] n5818_6;
wire   [18:0] n5818_5;
wire   [17:0] n5818_4;
wire   [16:0] n5817_6;
wire   [15:0] n5817_5;
wire   [14:0] n5817_4;
wire   [18:0] n5823;
wire   [18:0] n5822_3;
wire   [18:0] n5822_2;
wire   [18:0] n5822;
wire   [18:0] n5821_3;
wire   [18:0] n5821_2;
wire   [18:0] n5821;
wire   [18:0] n5820_3;
wire   [18:0] n5820_2;
wire   [18:0] n5820;
wire   [18:0] n5819_3;
wire   [18:0] n5819_2;
wire   [18:0] n5819;
wire   [18:0] n5818_3;
wire   [18:0] n5818_2;
wire   [17:0] n5818;
wire   [16:0] n5817_3;
wire   [15:0] n5817_2;
wire   [14:0] n5817;
wire   [17:0] \out_reg[0] ;
wire   [17:0] \out_reg[1] ;
wire   [17:0] \out_reg[2] ;
wire   [17:0] \out_reg[3] ;
wire   [17:0] \out_reg[4] ;
wire   [17:0] \out_reg[5] ;
wire   [17:0] \out_reg[6] ;
wire   [17:0] \out_reg[7] ;
wire   [17:0] \out_reg[8] ;
wire   [17:0] \out_reg[9] ;
wire   [17:0] \row_output[0] ;
wire   [17:0] \row_output[1] ;
wire   [17:0] \row_output[2] ;
wire   [17:0] \row_output[3] ;
wire   [17:0] \row_output[4] ;
wire   [17:0] \row_output[5] ;
wire   [17:0] \row_output[6] ;
wire   [17:0] \row_output[7] ;
wire   [17:0] \row_output[8] ;
wire   [17:0] \row_output[9] ;
wire   [18:0] \row_sums[0] ;
wire   [18:0] \row_sums[1] ;
wire   [18:0] \row_sums[2] ;
wire   [18:0] \row_sums[3] ;
wire   [18:0] \row_sums[4] ;
wire   [18:0] \row_sums[5] ;
wire   [18:0] \row_sums[6] ;
wire   [18:0] \row_sums[7] ;
wire   [18:0] \row_sums[8] ;
wire   [18:0] \row_sums[9] ;
wire   [13:0] \b2_extended[0] ;
wire   [13:0] \b2_extended[1] ;
wire   [13:0] \b2_extended[2] ;
wire   [13:0] \b2_extended[3] ;
wire   [13:0] \b2_extended[4] ;
wire   [13:0] \b2_extended[5] ;
wire   [13:0] \b2_extended[6] ;
wire   [13:0] \b2_extended[7] ;
wire   [13:0] \b2_extended[8] ;
wire   [13:0] \b2_extended[9] ;
wire   [13:0] \prod_terms[0][0] ;
wire   [13:0] \prod_terms[0][1] ;
wire   [13:0] \prod_terms[0][2] ;
wire   [13:0] \prod_terms[0][3] ;
wire   [13:0] \prod_terms[0][4] ;
wire   [13:0] \prod_terms[0][5] ;
wire   [13:0] \prod_terms[0][6] ;
wire   [13:0] \prod_terms[0][7] ;
wire   [13:0] \prod_terms[0][8] ;
wire   [13:0] \prod_terms[0][9] ;
wire   [13:0] \prod_terms[0][10] ;
wire   [13:0] \prod_terms[0][11] ;
wire   [13:0] \prod_terms[0][12] ;
wire   [13:0] \prod_terms[0][13] ;
wire   [13:0] \prod_terms[0][14] ;
wire   [13:0] \prod_terms[0][15] ;
wire   [13:0] \prod_terms[0][16] ;
wire   [13:0] \prod_terms[0][17] ;
wire   [13:0] \prod_terms[0][18] ;
wire   [13:0] \prod_terms[0][19] ;
wire   [13:0] \prod_terms[1][0] ;
wire   [13:0] \prod_terms[1][1] ;
wire   [13:0] \prod_terms[1][2] ;
wire   [13:0] \prod_terms[1][3] ;
wire   [13:0] \prod_terms[1][4] ;
wire   [13:0] \prod_terms[1][5] ;
wire   [13:0] \prod_terms[1][6] ;
wire   [13:0] \prod_terms[1][7] ;
wire   [13:0] \prod_terms[1][8] ;
wire   [13:0] \prod_terms[1][9] ;
wire   [13:0] \prod_terms[1][10] ;
wire   [13:0] \prod_terms[1][11] ;
wire   [13:0] \prod_terms[1][12] ;
wire   [13:0] \prod_terms[1][13] ;
wire   [13:0] \prod_terms[1][14] ;
wire   [13:0] \prod_terms[1][15] ;
wire   [13:0] \prod_terms[1][16] ;
wire   [13:0] \prod_terms[1][17] ;
wire   [13:0] \prod_terms[1][18] ;
wire   [13:0] \prod_terms[1][19] ;
wire   [13:0] \prod_terms[2][0] ;
wire   [13:0] \prod_terms[2][1] ;
wire   [13:0] \prod_terms[2][2] ;
wire   [13:0] \prod_terms[2][3] ;
wire   [13:0] \prod_terms[2][4] ;
wire   [13:0] \prod_terms[2][5] ;
wire   [13:0] \prod_terms[2][6] ;
wire   [13:0] \prod_terms[2][7] ;
wire   [13:0] \prod_terms[2][8] ;
wire   [13:0] \prod_terms[2][9] ;
wire   [13:0] \prod_terms[2][10] ;
wire   [13:0] \prod_terms[2][11] ;
wire   [13:0] \prod_terms[2][12] ;
wire   [13:0] \prod_terms[2][13] ;
wire   [13:0] \prod_terms[2][14] ;
wire   [13:0] \prod_terms[2][15] ;
wire   [13:0] \prod_terms[2][16] ;
wire   [13:0] \prod_terms[2][17] ;
wire   [13:0] \prod_terms[2][18] ;
wire   [13:0] \prod_terms[2][19] ;
wire   [13:0] \prod_terms[3][0] ;
wire   [13:0] \prod_terms[3][1] ;
wire   [13:0] \prod_terms[3][2] ;
wire   [13:0] \prod_terms[3][3] ;
wire   [13:0] \prod_terms[3][4] ;
wire   [13:0] \prod_terms[3][5] ;
wire   [13:0] \prod_terms[3][6] ;
wire   [13:0] \prod_terms[3][7] ;
wire   [13:0] \prod_terms[3][8] ;
wire   [13:0] \prod_terms[3][9] ;
wire   [13:0] \prod_terms[3][10] ;
wire   [13:0] \prod_terms[3][11] ;
wire   [13:0] \prod_terms[3][12] ;
wire   [13:0] \prod_terms[3][13] ;
wire   [13:0] \prod_terms[3][14] ;
wire   [13:0] \prod_terms[3][15] ;
wire   [13:0] \prod_terms[3][16] ;
wire   [13:0] \prod_terms[3][17] ;
wire   [13:0] \prod_terms[3][18] ;
wire   [13:0] \prod_terms[3][19] ;
wire   [13:0] \prod_terms[4][0] ;
wire   [13:0] \prod_terms[4][1] ;
wire   [13:0] \prod_terms[4][2] ;
wire   [13:0] \prod_terms[4][3] ;
wire   [13:0] \prod_terms[4][4] ;
wire   [13:0] \prod_terms[4][5] ;
wire   [13:0] \prod_terms[4][6] ;
wire   [13:0] \prod_terms[4][7] ;
wire   [13:0] \prod_terms[4][8] ;
wire   [13:0] \prod_terms[4][9] ;
wire   [13:0] \prod_terms[4][10] ;
wire   [13:0] \prod_terms[4][11] ;
wire   [13:0] \prod_terms[4][12] ;
wire   [13:0] \prod_terms[4][13] ;
wire   [13:0] \prod_terms[4][14] ;
wire   [13:0] \prod_terms[4][15] ;
wire   [13:0] \prod_terms[4][16] ;
wire   [13:0] \prod_terms[4][17] ;
wire   [13:0] \prod_terms[4][18] ;
wire   [13:0] \prod_terms[4][19] ;
wire   [13:0] \prod_terms[5][0] ;
wire   [13:0] \prod_terms[5][1] ;
wire   [13:0] \prod_terms[5][2] ;
wire   [13:0] \prod_terms[5][3] ;
wire   [13:0] \prod_terms[5][4] ;
wire   [13:0] \prod_terms[5][5] ;
wire   [13:0] \prod_terms[5][6] ;
wire   [13:0] \prod_terms[5][7] ;
wire   [13:0] \prod_terms[5][8] ;
wire   [13:0] \prod_terms[5][9] ;
wire   [13:0] \prod_terms[5][10] ;
wire   [13:0] \prod_terms[5][11] ;
wire   [13:0] \prod_terms[5][12] ;
wire   [13:0] \prod_terms[5][13] ;
wire   [13:0] \prod_terms[5][14] ;
wire   [13:0] \prod_terms[5][15] ;
wire   [13:0] \prod_terms[5][16] ;
wire   [13:0] \prod_terms[5][17] ;
wire   [13:0] \prod_terms[5][18] ;
wire   [13:0] \prod_terms[5][19] ;
wire   [13:0] \prod_terms[6][0] ;
wire   [13:0] \prod_terms[6][1] ;
wire   [13:0] \prod_terms[6][2] ;
wire   [13:0] \prod_terms[6][3] ;
wire   [13:0] \prod_terms[6][4] ;
wire   [13:0] \prod_terms[6][5] ;
wire   [13:0] \prod_terms[6][6] ;
wire   [13:0] \prod_terms[6][7] ;
wire   [13:0] \prod_terms[6][8] ;
wire   [13:0] \prod_terms[6][9] ;
wire   [13:0] \prod_terms[6][10] ;
wire   [13:0] \prod_terms[6][11] ;
wire   [13:0] \prod_terms[6][12] ;
wire   [13:0] \prod_terms[6][13] ;
wire   [13:0] \prod_terms[6][14] ;
wire   [13:0] \prod_terms[6][15] ;
wire   [13:0] \prod_terms[6][16] ;
wire   [13:0] \prod_terms[6][17] ;
wire   [13:0] \prod_terms[6][18] ;
wire   [13:0] \prod_terms[6][19] ;
wire   [13:0] \prod_terms[7][0] ;
wire   [13:0] \prod_terms[7][1] ;
wire   [13:0] \prod_terms[7][2] ;
wire   [13:0] \prod_terms[7][3] ;
wire   [13:0] \prod_terms[7][4] ;
wire   [13:0] \prod_terms[7][5] ;
wire   [13:0] \prod_terms[7][6] ;
wire   [13:0] \prod_terms[7][7] ;
wire   [13:0] \prod_terms[7][8] ;
wire   [13:0] \prod_terms[7][9] ;
wire   [13:0] \prod_terms[7][10] ;
wire   [13:0] \prod_terms[7][11] ;
wire   [13:0] \prod_terms[7][12] ;
wire   [13:0] \prod_terms[7][13] ;
wire   [13:0] \prod_terms[7][14] ;
wire   [13:0] \prod_terms[7][15] ;
wire   [13:0] \prod_terms[7][16] ;
wire   [13:0] \prod_terms[7][17] ;
wire   [13:0] \prod_terms[7][18] ;
wire   [13:0] \prod_terms[7][19] ;
wire   [13:0] \prod_terms[8][0] ;
wire   [13:0] \prod_terms[8][1] ;
wire   [13:0] \prod_terms[8][2] ;
wire   [13:0] \prod_terms[8][3] ;
wire   [13:0] \prod_terms[8][4] ;
wire   [13:0] \prod_terms[8][5] ;
wire   [13:0] \prod_terms[8][6] ;
wire   [13:0] \prod_terms[8][7] ;
wire   [13:0] \prod_terms[8][8] ;
wire   [13:0] \prod_terms[8][9] ;
wire   [13:0] \prod_terms[8][10] ;
wire   [13:0] \prod_terms[8][11] ;
wire   [13:0] \prod_terms[8][12] ;
wire   [13:0] \prod_terms[8][13] ;
wire   [13:0] \prod_terms[8][14] ;
wire   [13:0] \prod_terms[8][15] ;
wire   [13:0] \prod_terms[8][16] ;
wire   [13:0] \prod_terms[8][17] ;
wire   [13:0] \prod_terms[8][18] ;
wire   [13:0] \prod_terms[8][19] ;
wire   [13:0] \prod_terms[9][0] ;
wire   [13:0] \prod_terms[9][1] ;
wire   [13:0] \prod_terms[9][2] ;
wire   [13:0] \prod_terms[9][3] ;
wire   [13:0] \prod_terms[9][4] ;
wire   [13:0] \prod_terms[9][5] ;
wire   [13:0] \prod_terms[9][6] ;
wire   [13:0] \prod_terms[9][7] ;
wire   [13:0] \prod_terms[9][8] ;
wire   [13:0] \prod_terms[9][9] ;
wire   [13:0] \prod_terms[9][10] ;
wire   [13:0] \prod_terms[9][11] ;
wire   [13:0] \prod_terms[9][12] ;
wire   [13:0] \prod_terms[9][13] ;
wire   [13:0] \prod_terms[9][14] ;
wire   [13:0] \prod_terms[9][15] ;
wire   [13:0] \prod_terms[9][16] ;
wire   [13:0] \prod_terms[9][17] ;
wire   [13:0] \prod_terms[9][18] ;
wire   [13:0] \prod_terms[9][19] ;
wire   [5:0] \biases_l2[0] ;
wire   [5:0] \biases_l2[1] ;
wire   [5:0] \biases_l2[2] ;
wire   [5:0] \biases_l2[3] ;
wire   [5:0] \biases_l2[4] ;
wire   [5:0] \biases_l2[5] ;
wire   [5:0] \biases_l2[6] ;
wire   [5:0] \biases_l2[7] ;
wire   [5:0] \biases_l2[8] ;
wire   [5:0] \biases_l2[9] ;
wire   [4:0] \w2[0][0] ;
wire   [4:0] \w2[0][1] ;
wire   [4:0] \w2[0][2] ;
wire   [4:0] \w2[0][3] ;
wire   [4:0] \w2[0][4] ;
wire   [4:0] \w2[0][5] ;
wire   [4:0] \w2[0][6] ;
wire   [4:0] \w2[0][7] ;
wire   [4:0] \w2[0][8] ;
wire   [4:0] \w2[0][9] ;
wire   [4:0] \w2[0][10] ;
wire   [4:0] \w2[0][11] ;
wire   [4:0] \w2[0][12] ;
wire   [4:0] \w2[0][13] ;
wire   [4:0] \w2[0][14] ;
wire   [4:0] \w2[0][15] ;
wire   [4:0] \w2[0][16] ;
wire   [4:0] \w2[0][17] ;
wire   [4:0] \w2[0][18] ;
wire   [4:0] \w2[0][19] ;
wire   [4:0] \w2[1][0] ;
wire   [4:0] \w2[1][1] ;
wire   [4:0] \w2[1][2] ;
wire   [4:0] \w2[1][3] ;
wire   [4:0] \w2[1][4] ;
wire   [4:0] \w2[1][5] ;
wire   [4:0] \w2[1][6] ;
wire   [4:0] \w2[1][7] ;
wire   [4:0] \w2[1][8] ;
wire   [4:0] \w2[1][9] ;
wire   [4:0] \w2[1][10] ;
wire   [4:0] \w2[1][11] ;
wire   [4:0] \w2[1][12] ;
wire   [4:0] \w2[1][13] ;
wire   [4:0] \w2[1][14] ;
wire   [4:0] \w2[1][15] ;
wire   [4:0] \w2[1][16] ;
wire   [4:0] \w2[1][17] ;
wire   [4:0] \w2[1][18] ;
wire   [4:0] \w2[1][19] ;
wire   [4:0] \w2[2][0] ;
wire   [4:0] \w2[2][1] ;
wire   [4:0] \w2[2][2] ;
wire   [4:0] \w2[2][3] ;
wire   [4:0] \w2[2][4] ;
wire   [4:0] \w2[2][5] ;
wire   [4:0] \w2[2][6] ;
wire   [4:0] \w2[2][7] ;
wire   [4:0] \w2[2][8] ;
wire   [4:0] \w2[2][9] ;
wire   [4:0] \w2[2][10] ;
wire   [4:0] \w2[2][11] ;
wire   [4:0] \w2[2][12] ;
wire   [4:0] \w2[2][13] ;
wire   [4:0] \w2[2][14] ;
wire   [4:0] \w2[2][15] ;
wire   [4:0] \w2[2][16] ;
wire   [4:0] \w2[2][17] ;
wire   [4:0] \w2[2][18] ;
wire   [4:0] \w2[2][19] ;
wire   [4:0] \w2[3][0] ;
wire   [4:0] \w2[3][1] ;
wire   [4:0] \w2[3][2] ;
wire   [4:0] \w2[3][3] ;
wire   [4:0] \w2[3][4] ;
wire   [4:0] \w2[3][5] ;
wire   [4:0] \w2[3][6] ;
wire   [4:0] \w2[3][7] ;
wire   [4:0] \w2[3][8] ;
wire   [4:0] \w2[3][9] ;
wire   [4:0] \w2[3][10] ;
wire   [4:0] \w2[3][11] ;
wire   [4:0] \w2[3][12] ;
wire   [4:0] \w2[3][13] ;
wire   [4:0] \w2[3][14] ;
wire   [4:0] \w2[3][15] ;
wire   [4:0] \w2[3][16] ;
wire   [4:0] \w2[3][17] ;
wire   [4:0] \w2[3][18] ;
wire   [4:0] \w2[3][19] ;
wire   [4:0] \w2[4][0] ;
wire   [4:0] \w2[4][1] ;
wire   [4:0] \w2[4][2] ;
wire   [4:0] \w2[4][3] ;
wire   [4:0] \w2[4][4] ;
wire   [4:0] \w2[4][5] ;
wire   [4:0] \w2[4][6] ;
wire   [4:0] \w2[4][7] ;
wire   [4:0] \w2[4][8] ;
wire   [4:0] \w2[4][9] ;
wire   [4:0] \w2[4][10] ;
wire   [4:0] \w2[4][11] ;
wire   [4:0] \w2[4][12] ;
wire   [4:0] \w2[4][13] ;
wire   [4:0] \w2[4][14] ;
wire   [4:0] \w2[4][15] ;
wire   [4:0] \w2[4][16] ;
wire   [4:0] \w2[4][17] ;
wire   [4:0] \w2[4][18] ;
wire   [4:0] \w2[4][19] ;
wire   [4:0] \w2[5][0] ;
wire   [4:0] \w2[5][1] ;
wire   [4:0] \w2[5][2] ;
wire   [4:0] \w2[5][3] ;
wire   [4:0] \w2[5][4] ;
wire   [4:0] \w2[5][5] ;
wire   [4:0] \w2[5][6] ;
wire   [4:0] \w2[5][7] ;
wire   [4:0] \w2[5][8] ;
wire   [4:0] \w2[5][9] ;
wire   [4:0] \w2[5][10] ;
wire   [4:0] \w2[5][11] ;
wire   [4:0] \w2[5][12] ;
wire   [4:0] \w2[5][13] ;
wire   [4:0] \w2[5][14] ;
wire   [4:0] \w2[5][15] ;
wire   [4:0] \w2[5][16] ;
wire   [4:0] \w2[5][17] ;
wire   [4:0] \w2[5][18] ;
wire   [4:0] \w2[5][19] ;
wire   [4:0] \w2[6][0] ;
wire   [4:0] \w2[6][1] ;
wire   [4:0] \w2[6][2] ;
wire   [4:0] \w2[6][3] ;
wire   [4:0] \w2[6][4] ;
wire   [4:0] \w2[6][5] ;
wire   [4:0] \w2[6][6] ;
wire   [4:0] \w2[6][7] ;
wire   [4:0] \w2[6][8] ;
wire   [4:0] \w2[6][9] ;
wire   [4:0] \w2[6][10] ;
wire   [4:0] \w2[6][11] ;
wire   [4:0] \w2[6][12] ;
wire   [4:0] \w2[6][13] ;
wire   [4:0] \w2[6][14] ;
wire   [4:0] \w2[6][15] ;
wire   [4:0] \w2[6][16] ;
wire   [4:0] \w2[6][17] ;
wire   [4:0] \w2[6][18] ;
wire   [4:0] \w2[6][19] ;
wire   [4:0] \w2[7][0] ;
wire   [4:0] \w2[7][1] ;
wire   [4:0] \w2[7][2] ;
wire   [4:0] \w2[7][3] ;
wire   [4:0] \w2[7][4] ;
wire   [4:0] \w2[7][5] ;
wire   [4:0] \w2[7][6] ;
wire   [4:0] \w2[7][7] ;
wire   [4:0] \w2[7][8] ;
wire   [4:0] \w2[7][9] ;
wire   [4:0] \w2[7][10] ;
wire   [4:0] \w2[7][11] ;
wire   [4:0] \w2[7][12] ;
wire   [4:0] \w2[7][13] ;
wire   [4:0] \w2[7][14] ;
wire   [4:0] \w2[7][15] ;
wire   [4:0] \w2[7][16] ;
wire   [4:0] \w2[7][17] ;
wire   [4:0] \w2[7][18] ;
wire   [4:0] \w2[7][19] ;
wire   [4:0] \w2[8][0] ;
wire   [4:0] \w2[8][1] ;
wire   [4:0] \w2[8][2] ;
wire   [4:0] \w2[8][3] ;
wire   [4:0] \w2[8][4] ;
wire   [4:0] \w2[8][5] ;
wire   [4:0] \w2[8][6] ;
wire   [4:0] \w2[8][7] ;
wire   [4:0] \w2[8][8] ;
wire   [4:0] \w2[8][9] ;
wire   [4:0] \w2[8][10] ;
wire   [4:0] \w2[8][11] ;
wire   [4:0] \w2[8][12] ;
wire   [4:0] \w2[8][13] ;
wire   [4:0] \w2[8][14] ;
wire   [4:0] \w2[8][15] ;
wire   [4:0] \w2[8][16] ;
wire   [4:0] \w2[8][17] ;
wire   [4:0] \w2[8][18] ;
wire   [4:0] \w2[8][19] ;
wire   [4:0] \w2[9][0] ;
wire   [4:0] \w2[9][1] ;
wire   [4:0] \w2[9][2] ;
wire   [4:0] \w2[9][3] ;
wire   [4:0] \w2[9][4] ;
wire   [4:0] \w2[9][5] ;
wire   [4:0] \w2[9][6] ;
wire   [4:0] \w2[9][7] ;
wire   [4:0] \w2[9][8] ;
wire   [4:0] \w2[9][9] ;
wire   [4:0] \w2[9][10] ;
wire   [4:0] \w2[9][11] ;
wire   [4:0] \w2[9][12] ;
wire   [4:0] \w2[9][13] ;
wire   [4:0] \w2[9][14] ;
wire   [4:0] \w2[9][15] ;
wire   [4:0] \w2[9][16] ;
wire   [4:0] \w2[9][17] ;
wire   [4:0] \w2[9][18] ;
wire   [4:0] \w2[9][19] ;
wire   [179:0] out;
wire   [179:0] in;
  assign N$1 = 1'b0;
  assign N$2 = 1'b0;
  assign N$3 = 1'b0;
  assign N$4 = 1'b0;
  assign N$5 = 1'b0;
  assign N$6 = 1'b0;
  assign N$7 = 1'b0;
  assign N$8 = 1'b0;
  assign N$9 = 1'b0;
  assign N$10 = 1'b0;
  assign N$11 = 1'b0;
  assign N$12 = 1'b0;
  assign N$13 = 1'b0;
  assign N$14 = 1'b0;
  assign N$15 = 1'b0;
  assign N$16 = 1'b0;
  assign N$17 = 1'b0;
  assign N$18 = 1'b0;
  assign \b2_extended[0] [3] = 1'b0;
  assign \b2_extended[0] [2] = 1'b0;
  assign \b2_extended[0] [1] = 1'b0;
  assign \b2_extended[0] [0] = 1'b0;
  assign \b2_extended[1] [3] = 1'b0;
  assign \b2_extended[1] [2] = 1'b0;
  assign \b2_extended[1] [1] = 1'b0;
  assign \b2_extended[1] [0] = 1'b0;
  assign \b2_extended[2] [3] = 1'b0;
  assign \b2_extended[2] [2] = 1'b0;
  assign \b2_extended[2] [1] = 1'b0;
  assign \b2_extended[2] [0] = 1'b0;
  assign \b2_extended[3] [3] = 1'b0;
  assign \b2_extended[3] [2] = 1'b0;
  assign \b2_extended[3] [1] = 1'b0;
  assign \b2_extended[3] [0] = 1'b0;
  assign \b2_extended[4] [3] = 1'b0;
  assign \b2_extended[4] [2] = 1'b0;
  assign \b2_extended[4] [1] = 1'b0;
  assign \b2_extended[4] [0] = 1'b0;
  assign \b2_extended[5] [3] = 1'b0;
  assign \b2_extended[5] [2] = 1'b0;
  assign \b2_extended[5] [1] = 1'b0;
  assign \b2_extended[5] [0] = 1'b0;
  assign \b2_extended[6] [3] = 1'b0;
  assign \b2_extended[6] [2] = 1'b0;
  assign \b2_extended[6] [1] = 1'b0;
  assign \b2_extended[6] [0] = 1'b0;
  assign \b2_extended[7] [3] = 1'b0;
  assign \b2_extended[7] [2] = 1'b0;
  assign \b2_extended[7] [1] = 1'b0;
  assign \b2_extended[7] [0] = 1'b0;
  assign \b2_extended[8] [3] = 1'b0;
  assign \b2_extended[8] [2] = 1'b0;
  assign \b2_extended[8] [1] = 1'b0;
  assign \b2_extended[8] [0] = 1'b0;
  assign \b2_extended[9] [3] = 1'b0;
  assign \b2_extended[9] [2] = 1'b0;
  assign \b2_extended[9] [1] = 1'b0;
  assign \b2_extended[9] [0] = 1'b0;
  assign \biases_l2[0] [5] = 1'b0;
  assign \biases_l2[0] [4] = 1'b0;
  assign \biases_l2[0] [2] = 1'b0;
  assign \biases_l2[0] [1] = 1'b0;
  assign \biases_l2[1] [5] = 1'b0;
  assign \biases_l2[1] [4] = 1'b0;
  assign \biases_l2[1] [1] = 1'b0;
  assign \biases_l2[2] [0] = 1'b0;
  assign \biases_l2[3] [2] = 1'b0;
  assign \biases_l2[3] [1] = 1'b0;
  assign \biases_l2[4] [3] = 1'b0;
  assign \biases_l2[4] [2] = 1'b0;
  assign \biases_l2[4] [1] = 1'b0;
  assign \biases_l2[5] [5] = 1'b0;
  assign \biases_l2[5] [4] = 1'b0;
  assign \biases_l2[5] [3] = 1'b0;
  assign \biases_l2[5] [2] = 1'b0;
  assign \biases_l2[5] [0] = 1'b0;
  assign \biases_l2[6] [4] = 1'b0;
  assign \biases_l2[6] [1] = 1'b0;
  assign \biases_l2[7] [3] = 1'b0;
  assign \biases_l2[7] [0] = 1'b0;
  assign \biases_l2[8] [3] = 1'b0;
  assign \biases_l2[8] [2] = 1'b0;
  assign \biases_l2[8] [1] = 1'b0;
  assign \biases_l2[9] [5] = 1'b0;
  assign \biases_l2[9] [4] = 1'b0;
  assign \biases_l2[9] [3] = 1'b0;
  assign \biases_l2[9] [0] = 1'b0;
  assign \w2[0][0] [0] = 1'b0;
  assign \w2[0][1] [4] = 1'b0;
  assign \w2[0][1] [3] = 1'b0;
  assign \w2[0][1] [2] = 1'b0;
  assign \w2[0][2] [1] = 1'b0;
  assign \w2[0][3] [1] = 1'b0;
  assign \w2[0][4] [2] = 1'b0;
  assign \w2[0][4] [0] = 1'b0;
  assign \w2[0][5] [1] = 1'b0;
  assign \w2[0][6] [4] = 1'b0;
  assign \w2[0][6] [3] = 1'b0;
  assign \w2[0][6] [2] = 1'b0;
  assign \w2[0][6] [1] = 1'b0;
  assign \w2[0][7] [0] = 1'b0;
  assign \w2[0][8] [4] = 1'b0;
  assign \w2[0][8] [3] = 1'b0;
  assign \w2[0][8] [2] = 1'b0;
  assign \w2[0][8] [1] = 1'b0;
  assign \w2[0][8] [0] = 1'b0;
  assign \w2[0][9] [3] = 1'b0;
  assign \w2[0][10] [0] = 1'b0;
  assign \w2[0][12] [4] = 1'b0;
  assign \w2[0][12] [3] = 1'b0;
  assign \w2[0][12] [2] = 1'b0;
  assign \w2[0][12] [1] = 1'b0;
  assign \w2[0][13] [4] = 1'b0;
  assign \w2[0][13] [3] = 1'b0;
  assign \w2[0][13] [2] = 1'b0;
  assign \w2[0][13] [1] = 1'b0;
  assign \w2[0][14] [4] = 1'b0;
  assign \w2[0][14] [3] = 1'b0;
  assign \w2[0][14] [2] = 1'b0;
  assign \w2[0][15] [4] = 1'b0;
  assign \w2[0][15] [3] = 1'b0;
  assign \w2[0][15] [2] = 1'b0;
  assign \w2[0][15] [0] = 1'b0;
  assign \w2[0][17] [1] = 1'b0;
  assign \w2[0][18] [4] = 1'b0;
  assign \w2[0][18] [3] = 1'b0;
  assign \w2[0][18] [1] = 1'b0;
  assign \w2[0][18] [0] = 1'b0;
  assign \w2[0][19] [2] = 1'b0;
  assign \w2[1][0] [4] = 1'b0;
  assign \w2[1][0] [3] = 1'b0;
  assign \w2[1][0] [1] = 1'b0;
  assign \w2[1][0] [0] = 1'b0;
  assign \w2[1][1] [1] = 1'b0;
  assign \w2[1][2] [4] = 1'b0;
  assign \w2[1][2] [2] = 1'b0;
  assign \w2[1][2] [1] = 1'b0;
  assign \w2[1][3] [4] = 1'b0;
  assign \w2[1][3] [3] = 1'b0;
  assign \w2[1][3] [1] = 1'b0;
  assign \w2[1][4] [4] = 1'b0;
  assign \w2[1][4] [3] = 1'b0;
  assign \w2[1][4] [1] = 1'b0;
  assign \w2[1][5] [4] = 1'b0;
  assign \w2[1][5] [2] = 1'b0;
  assign \w2[1][5] [0] = 1'b0;
  assign \w2[1][6] [3] = 1'b0;
  assign \w2[1][7] [0] = 1'b0;
  assign \w2[1][8] [0] = 1'b0;
  assign \w2[1][9] [0] = 1'b0;
  assign \w2[1][10] [4] = 1'b0;
  assign \w2[1][10] [3] = 1'b0;
  assign \w2[1][10] [1] = 1'b0;
  assign \w2[1][11] [3] = 1'b0;
  assign \w2[1][11] [0] = 1'b0;
  assign \w2[1][12] [4] = 1'b0;
  assign \w2[1][12] [3] = 1'b0;
  assign \w2[1][12] [1] = 1'b0;
  assign \w2[1][12] [0] = 1'b0;
  assign \w2[1][13] [2] = 1'b0;
  assign \w2[1][14] [3] = 1'b0;
  assign \w2[1][14] [2] = 1'b0;
  assign \w2[1][15] [4] = 1'b0;
  assign \w2[1][15] [3] = 1'b0;
  assign \w2[1][16] [4] = 1'b0;
  assign \w2[1][16] [3] = 1'b0;
  assign \w2[1][17] [1] = 1'b0;
  assign \w2[1][18] [4] = 1'b0;
  assign \w2[1][18] [3] = 1'b0;
  assign \w2[1][18] [2] = 1'b0;
  assign \w2[1][18] [0] = 1'b0;
  assign \w2[1][19] [1] = 1'b0;
  assign \w2[1][19] [0] = 1'b0;
  assign \w2[2][0] [2] = 1'b0;
  assign \w2[2][2] [2] = 1'b0;
  assign \w2[2][2] [1] = 1'b0;
  assign \w2[2][2] [0] = 1'b0;
  assign \w2[2][4] [4] = 1'b0;
  assign \w2[2][4] [3] = 1'b0;
  assign \w2[2][4] [2] = 1'b0;
  assign \w2[2][4] [0] = 1'b0;
  assign \w2[2][5] [0] = 1'b0;
  assign \w2[2][6] [2] = 1'b0;
  assign \w2[2][6] [0] = 1'b0;
  assign \w2[2][7] [0] = 1'b0;
  assign \w2[2][8] [4] = 1'b0;
  assign \w2[2][8] [3] = 1'b0;
  assign \w2[2][8] [1] = 1'b0;
  assign \w2[2][9] [1] = 1'b0;
  assign \w2[2][9] [0] = 1'b0;
  assign \w2[2][10] [4] = 1'b0;
  assign \w2[2][10] [3] = 1'b0;
  assign \w2[2][10] [1] = 1'b0;
  assign \w2[2][11] [3] = 1'b0;
  assign \w2[2][11] [1] = 1'b0;
  assign \w2[2][12] [4] = 1'b0;
  assign \w2[2][12] [3] = 1'b0;
  assign \w2[2][12] [2] = 1'b0;
  assign \w2[2][12] [1] = 1'b0;
  assign \w2[2][12] [0] = 1'b0;
  assign \w2[2][13] [4] = 1'b0;
  assign \w2[2][13] [3] = 1'b0;
  assign \w2[2][14] [4] = 1'b0;
  assign \w2[2][14] [3] = 1'b0;
  assign \w2[2][14] [2] = 1'b0;
  assign \w2[2][14] [1] = 1'b0;
  assign \w2[2][15] [4] = 1'b0;
  assign \w2[2][15] [3] = 1'b0;
  assign \w2[2][15] [2] = 1'b0;
  assign \w2[2][15] [1] = 1'b0;
  assign \w2[2][15] [0] = 1'b0;
  assign \w2[2][16] [4] = 1'b0;
  assign \w2[2][16] [2] = 1'b0;
  assign \w2[2][17] [4] = 1'b0;
  assign \w2[2][17] [3] = 1'b0;
  assign \w2[2][17] [1] = 1'b0;
  assign \w2[2][17] [0] = 1'b0;
  assign \w2[2][18] [4] = 1'b0;
  assign \w2[2][18] [3] = 1'b0;
  assign \w2[2][18] [2] = 1'b0;
  assign \w2[2][18] [1] = 1'b0;
  assign \w2[2][18] [0] = 1'b0;
  assign \w2[2][19] [4] = 1'b0;
  assign \w2[2][19] [3] = 1'b0;
  assign \w2[2][19] [2] = 1'b0;
  assign \w2[2][19] [1] = 1'b0;
  assign \w2[3][0] [4] = 1'b0;
  assign \w2[3][0] [3] = 1'b0;
  assign \w2[3][0] [2] = 1'b0;
  assign \w2[3][0] [1] = 1'b0;
  assign \w2[3][1] [1] = 1'b0;
  assign \w2[3][1] [0] = 1'b0;
  assign \w2[3][2] [2] = 1'b0;
  assign \w2[3][2] [1] = 1'b0;
  assign \w2[3][2] [0] = 1'b0;
  assign \w2[3][3] [2] = 1'b0;
  assign \w2[3][3] [1] = 1'b0;
  assign \w2[3][3] [0] = 1'b0;
  assign \w2[3][4] [4] = 1'b0;
  assign \w2[3][4] [3] = 1'b0;
  assign \w2[3][4] [2] = 1'b0;
  assign \w2[3][4] [0] = 1'b0;
  assign \w2[3][5] [4] = 1'b0;
  assign \w2[3][5] [3] = 1'b0;
  assign \w2[3][5] [2] = 1'b0;
  assign \w2[3][5] [0] = 1'b0;
  assign \w2[3][6] [1] = 1'b0;
  assign \w2[3][6] [0] = 1'b0;
  assign \w2[3][7] [4] = 1'b0;
  assign \w2[3][7] [3] = 1'b0;
  assign \w2[3][7] [2] = 1'b0;
  assign \w2[3][8] [3] = 1'b0;
  assign \w2[3][9] [4] = 1'b0;
  assign \w2[3][9] [3] = 1'b0;
  assign \w2[3][9] [2] = 1'b0;
  assign \w2[3][10] [4] = 1'b0;
  assign \w2[3][10] [3] = 1'b0;
  assign \w2[3][10] [2] = 1'b0;
  assign \w2[3][10] [1] = 1'b0;
  assign \w2[3][10] [0] = 1'b0;
  assign \w2[3][11] [4] = 1'b0;
  assign \w2[3][11] [3] = 1'b0;
  assign \w2[3][11] [2] = 1'b0;
  assign \w2[3][11] [0] = 1'b0;
  assign \w2[3][12] [1] = 1'b0;
  assign \w2[3][12] [0] = 1'b0;
  assign \w2[3][13] [4] = 1'b0;
  assign \w2[3][13] [3] = 1'b0;
  assign \w2[3][13] [2] = 1'b0;
  assign \w2[3][13] [1] = 1'b0;
  assign \w2[3][13] [0] = 1'b0;
  assign \w2[3][14] [4] = 1'b0;
  assign \w2[3][14] [3] = 1'b0;
  assign \w2[3][14] [1] = 1'b0;
  assign \w2[3][15] [4] = 1'b0;
  assign \w2[3][15] [3] = 1'b0;
  assign \w2[3][15] [2] = 1'b0;
  assign \w2[3][15] [1] = 1'b0;
  assign \w2[3][15] [0] = 1'b0;
  assign \w2[3][16] [4] = 1'b0;
  assign \w2[3][16] [3] = 1'b0;
  assign \w2[3][16] [2] = 1'b0;
  assign \w2[3][16] [1] = 1'b0;
  assign \w2[3][17] [4] = 1'b0;
  assign \w2[3][17] [3] = 1'b0;
  assign \w2[3][17] [1] = 1'b0;
  assign \w2[3][18] [4] = 1'b0;
  assign \w2[3][18] [3] = 1'b0;
  assign \w2[3][19] [4] = 1'b0;
  assign \w2[3][19] [3] = 1'b0;
  assign \w2[3][19] [1] = 1'b0;
  assign \w2[3][19] [0] = 1'b0;
  assign \w2[4][0] [4] = 1'b0;
  assign \w2[4][0] [3] = 1'b0;
  assign \w2[4][0] [2] = 1'b0;
  assign \w2[4][0] [1] = 1'b0;
  assign \w2[4][0] [0] = 1'b0;
  assign \w2[4][1] [4] = 1'b0;
  assign \w2[4][1] [3] = 1'b0;
  assign \w2[4][1] [2] = 1'b0;
  assign \w2[4][1] [0] = 1'b0;
  assign \w2[4][2] [4] = 1'b0;
  assign \w2[4][2] [2] = 1'b0;
  assign \w2[4][2] [0] = 1'b0;
  assign \w2[4][3] [1] = 1'b0;
  assign \w2[4][4] [4] = 1'b0;
  assign \w2[4][4] [3] = 1'b0;
  assign \w2[4][4] [1] = 1'b0;
  assign \w2[4][4] [0] = 1'b0;
  assign \w2[4][5] [4] = 1'b0;
  assign \w2[4][5] [3] = 1'b0;
  assign \w2[4][5] [2] = 1'b0;
  assign \w2[4][5] [0] = 1'b0;
  assign \w2[4][6] [4] = 1'b0;
  assign \w2[4][6] [3] = 1'b0;
  assign \w2[4][6] [1] = 1'b0;
  assign \w2[4][7] [1] = 1'b0;
  assign \w2[4][7] [0] = 1'b0;
  assign \w2[4][8] [4] = 1'b0;
  assign \w2[4][8] [3] = 1'b0;
  assign \w2[4][8] [2] = 1'b0;
  assign \w2[4][8] [1] = 1'b0;
  assign \w2[4][9] [0] = 1'b0;
  assign \w2[4][10] [4] = 1'b0;
  assign \w2[4][10] [3] = 1'b0;
  assign \w2[4][10] [2] = 1'b0;
  assign \w2[4][10] [1] = 1'b0;
  assign \w2[4][10] [0] = 1'b0;
  assign \w2[4][11] [4] = 1'b0;
  assign \w2[4][11] [3] = 1'b0;
  assign \w2[4][11] [1] = 1'b0;
  assign \w2[4][12] [2] = 1'b0;
  assign \w2[4][12] [1] = 1'b0;
  assign \w2[4][13] [4] = 1'b0;
  assign \w2[4][13] [3] = 1'b0;
  assign \w2[4][13] [2] = 1'b0;
  assign \w2[4][13] [1] = 1'b0;
  assign \w2[4][15] [4] = 1'b0;
  assign \w2[4][15] [3] = 1'b0;
  assign \w2[4][15] [2] = 1'b0;
  assign \w2[4][15] [0] = 1'b0;
  assign \w2[4][16] [0] = 1'b0;
  assign \w2[4][18] [1] = 1'b0;
  assign \w2[4][18] [0] = 1'b0;
  assign \w2[4][19] [4] = 1'b0;
  assign \w2[4][19] [3] = 1'b0;
  assign \w2[4][19] [2] = 1'b0;
  assign \w2[4][19] [0] = 1'b0;
  assign \w2[5][0] [4] = 1'b0;
  assign \w2[5][0] [2] = 1'b0;
  assign \w2[5][0] [1] = 1'b0;
  assign \w2[5][0] [0] = 1'b0;
  assign \w2[5][1] [4] = 1'b0;
  assign \w2[5][1] [3] = 1'b0;
  assign \w2[5][1] [2] = 1'b0;
  assign \w2[5][1] [0] = 1'b0;
  assign \w2[5][2] [4] = 1'b0;
  assign \w2[5][2] [3] = 1'b0;
  assign \w2[5][2] [2] = 1'b0;
  assign \w2[5][2] [1] = 1'b0;
  assign \w2[5][4] [1] = 1'b0;
  assign \w2[5][4] [0] = 1'b0;
  assign \w2[5][5] [1] = 1'b0;
  assign \w2[5][5] [0] = 1'b0;
  assign \w2[5][6] [4] = 1'b0;
  assign \w2[5][6] [3] = 1'b0;
  assign \w2[5][6] [2] = 1'b0;
  assign \w2[5][6] [0] = 1'b0;
  assign \w2[5][7] [4] = 1'b0;
  assign \w2[5][7] [3] = 1'b0;
  assign \w2[5][7] [2] = 1'b0;
  assign \w2[5][7] [1] = 1'b0;
  assign \w2[5][7] [0] = 1'b0;
  assign \w2[5][8] [0] = 1'b0;
  assign \w2[5][9] [1] = 1'b0;
  assign \w2[5][9] [0] = 1'b0;
  assign \w2[5][10] [4] = 1'b0;
  assign \w2[5][10] [3] = 1'b0;
  assign \w2[5][10] [1] = 1'b0;
  assign \w2[5][10] [0] = 1'b0;
  assign \w2[5][11] [1] = 1'b0;
  assign \w2[5][11] [0] = 1'b0;
  assign \w2[5][12] [1] = 1'b0;
  assign \w2[5][13] [1] = 1'b0;
  assign \w2[5][13] [0] = 1'b0;
  assign \w2[5][14] [4] = 1'b0;
  assign \w2[5][14] [3] = 1'b0;
  assign \w2[5][14] [2] = 1'b0;
  assign \w2[5][15] [4] = 1'b0;
  assign \w2[5][15] [3] = 1'b0;
  assign \w2[5][16] [0] = 1'b0;
  assign \w2[5][17] [3] = 1'b0;
  assign \w2[5][17] [0] = 1'b0;
  assign \w2[5][18] [1] = 1'b0;
  assign \w2[5][18] [0] = 1'b0;
  assign \w2[5][19] [4] = 1'b0;
  assign \w2[5][19] [3] = 1'b0;
  assign \w2[6][0] [4] = 1'b0;
  assign \w2[6][0] [3] = 1'b0;
  assign \w2[6][0] [2] = 1'b0;
  assign \w2[6][0] [0] = 1'b0;
  assign \w2[6][1] [4] = 1'b0;
  assign \w2[6][1] [2] = 1'b0;
  assign \w2[6][1] [1] = 1'b0;
  assign \w2[6][2] [3] = 1'b0;
  assign \w2[6][2] [0] = 1'b0;
  assign \w2[6][3] [4] = 1'b0;
  assign \w2[6][3] [3] = 1'b0;
  assign \w2[6][3] [2] = 1'b0;
  assign \w2[6][3] [1] = 1'b0;
  assign \w2[6][4] [4] = 1'b0;
  assign \w2[6][4] [3] = 1'b0;
  assign \w2[6][4] [2] = 1'b0;
  assign \w2[6][4] [1] = 1'b0;
  assign \w2[6][5] [3] = 1'b0;
  assign \w2[6][5] [0] = 1'b0;
  assign \w2[6][6] [4] = 1'b0;
  assign \w2[6][6] [3] = 1'b0;
  assign \w2[6][6] [2] = 1'b0;
  assign \w2[6][6] [1] = 1'b0;
  assign \w2[6][6] [0] = 1'b0;
  assign \w2[6][7] [4] = 1'b0;
  assign \w2[6][7] [3] = 1'b0;
  assign \w2[6][7] [2] = 1'b0;
  assign \w2[6][8] [4] = 1'b0;
  assign \w2[6][8] [3] = 1'b0;
  assign \w2[6][8] [2] = 1'b0;
  assign \w2[6][9] [1] = 1'b0;
  assign \w2[6][9] [0] = 1'b0;
  assign \w2[6][10] [3] = 1'b0;
  assign \w2[6][11] [4] = 1'b0;
  assign \w2[6][11] [3] = 1'b0;
  assign \w2[6][11] [0] = 1'b0;
  assign \w2[6][12] [2] = 1'b0;
  assign \w2[6][12] [1] = 1'b0;
  assign \w2[6][13] [4] = 1'b0;
  assign \w2[6][13] [3] = 1'b0;
  assign \w2[6][13] [2] = 1'b0;
  assign \w2[6][14] [1] = 1'b0;
  assign \w2[6][14] [0] = 1'b0;
  assign \w2[6][15] [3] = 1'b0;
  assign \w2[6][15] [2] = 1'b0;
  assign \w2[6][17] [0] = 1'b0;
  assign \w2[6][18] [4] = 1'b0;
  assign \w2[6][18] [3] = 1'b0;
  assign \w2[6][18] [2] = 1'b0;
  assign \w2[6][18] [1] = 1'b0;
  assign \w2[6][19] [4] = 1'b0;
  assign \w2[6][19] [3] = 1'b0;
  assign \w2[6][19] [2] = 1'b0;
  assign \w2[6][19] [1] = 1'b0;
  assign \w2[7][0] [4] = 1'b0;
  assign \w2[7][0] [3] = 1'b0;
  assign \w2[7][0] [2] = 1'b0;
  assign \w2[7][0] [1] = 1'b0;
  assign \w2[7][0] [0] = 1'b0;
  assign \w2[7][1] [4] = 1'b0;
  assign \w2[7][1] [2] = 1'b0;
  assign \w2[7][1] [1] = 1'b0;
  assign \w2[7][3] [3] = 1'b0;
  assign \w2[7][4] [2] = 1'b0;
  assign \w2[7][4] [1] = 1'b0;
  assign \w2[7][5] [2] = 1'b0;
  assign \w2[7][5] [1] = 1'b0;
  assign \w2[7][6] [2] = 1'b0;
  assign \w2[7][6] [0] = 1'b0;
  assign \w2[7][8] [4] = 1'b0;
  assign \w2[7][8] [3] = 1'b0;
  assign \w2[7][8] [1] = 1'b0;
  assign \w2[7][9] [4] = 1'b0;
  assign \w2[7][9] [2] = 1'b0;
  assign \w2[7][9] [1] = 1'b0;
  assign \w2[7][10] [4] = 1'b0;
  assign \w2[7][10] [3] = 1'b0;
  assign \w2[7][10] [2] = 1'b0;
  assign \w2[7][10] [1] = 1'b0;
  assign \w2[7][10] [0] = 1'b0;
  assign \w2[7][11] [0] = 1'b0;
  assign \w2[7][12] [4] = 1'b0;
  assign \w2[7][12] [3] = 1'b0;
  assign \w2[7][12] [0] = 1'b0;
  assign \w2[7][13] [4] = 1'b0;
  assign \w2[7][13] [3] = 1'b0;
  assign \w2[7][13] [2] = 1'b0;
  assign \w2[7][13] [1] = 1'b0;
  assign \w2[7][13] [0] = 1'b0;
  assign \w2[7][14] [4] = 1'b0;
  assign \w2[7][14] [3] = 1'b0;
  assign \w2[7][14] [2] = 1'b0;
  assign \w2[7][14] [1] = 1'b0;
  assign \w2[7][15] [3] = 1'b0;
  assign \w2[7][16] [4] = 1'b0;
  assign \w2[7][16] [3] = 1'b0;
  assign \w2[7][16] [1] = 1'b0;
  assign \w2[7][16] [0] = 1'b0;
  assign \w2[7][17] [3] = 1'b0;
  assign \w2[7][18] [4] = 1'b0;
  assign \w2[7][18] [3] = 1'b0;
  assign \w2[7][18] [2] = 1'b0;
  assign \w2[7][19] [4] = 1'b0;
  assign \w2[7][19] [3] = 1'b0;
  assign \w2[7][19] [2] = 1'b0;
  assign \w2[7][19] [1] = 1'b0;
  assign \w2[7][19] [0] = 1'b0;
  assign \w2[8][0] [2] = 1'b0;
  assign \w2[8][0] [1] = 1'b0;
  assign \w2[8][1] [4] = 1'b0;
  assign \w2[8][1] [3] = 1'b0;
  assign \w2[8][1] [1] = 1'b0;
  assign \w2[8][1] [0] = 1'b0;
  assign \w2[8][2] [1] = 1'b0;
  assign \w2[8][2] [0] = 1'b0;
  assign \w2[8][3] [4] = 1'b0;
  assign \w2[8][3] [3] = 1'b0;
  assign \w2[8][3] [2] = 1'b0;
  assign \w2[8][3] [0] = 1'b0;
  assign \w2[8][4] [4] = 1'b0;
  assign \w2[8][4] [3] = 1'b0;
  assign \w2[8][4] [2] = 1'b0;
  assign \w2[8][4] [1] = 1'b0;
  assign \w2[8][4] [0] = 1'b0;
  assign \w2[8][5] [4] = 1'b0;
  assign \w2[8][5] [3] = 1'b0;
  assign \w2[8][5] [2] = 1'b0;
  assign \w2[8][5] [1] = 1'b0;
  assign \w2[8][6] [4] = 1'b0;
  assign \w2[8][6] [3] = 1'b0;
  assign \w2[8][6] [2] = 1'b0;
  assign \w2[8][6] [0] = 1'b0;
  assign \w2[8][7] [4] = 1'b0;
  assign \w2[8][7] [2] = 1'b0;
  assign \w2[8][7] [0] = 1'b0;
  assign \w2[8][8] [4] = 1'b0;
  assign \w2[8][8] [3] = 1'b0;
  assign \w2[8][8] [2] = 1'b0;
  assign \w2[8][9] [4] = 1'b0;
  assign \w2[8][9] [3] = 1'b0;
  assign \w2[8][9] [2] = 1'b0;
  assign \w2[8][9] [1] = 1'b0;
  assign \w2[8][10] [4] = 1'b0;
  assign \w2[8][10] [3] = 1'b0;
  assign \w2[8][10] [2] = 1'b0;
  assign \w2[8][10] [1] = 1'b0;
  assign \w2[8][10] [0] = 1'b0;
  assign \w2[8][11] [3] = 1'b0;
  assign \w2[8][11] [1] = 1'b0;
  assign \w2[8][11] [0] = 1'b0;
  assign \w2[8][12] [4] = 1'b0;
  assign \w2[8][12] [3] = 1'b0;
  assign \w2[8][12] [2] = 1'b0;
  assign \w2[8][12] [1] = 1'b0;
  assign \w2[8][12] [0] = 1'b0;
  assign \w2[8][13] [4] = 1'b0;
  assign \w2[8][13] [3] = 1'b0;
  assign \w2[8][13] [2] = 1'b0;
  assign \w2[8][13] [0] = 1'b0;
  assign \w2[8][14] [1] = 1'b0;
  assign \w2[8][15] [4] = 1'b0;
  assign \w2[8][15] [3] = 1'b0;
  assign \w2[8][15] [0] = 1'b0;
  assign \w2[8][18] [2] = 1'b0;
  assign \w2[8][18] [0] = 1'b0;
  assign \w2[8][19] [3] = 1'b0;
  assign \w2[8][19] [2] = 1'b0;
  assign \w2[9][0] [2] = 1'b0;
  assign \w2[9][0] [1] = 1'b0;
  assign \w2[9][0] [0] = 1'b0;
  assign \w2[9][1] [4] = 1'b0;
  assign \w2[9][1] [3] = 1'b0;
  assign \w2[9][1] [0] = 1'b0;
  assign \w2[9][2] [3] = 1'b0;
  assign \w2[9][3] [4] = 1'b0;
  assign \w2[9][3] [2] = 1'b0;
  assign \w2[9][3] [1] = 1'b0;
  assign \w2[9][4] [3] = 1'b0;
  assign \w2[9][6] [4] = 1'b0;
  assign \w2[9][6] [3] = 1'b0;
  assign \w2[9][6] [1] = 1'b0;
  assign \w2[9][6] [0] = 1'b0;
  assign \w2[9][7] [1] = 1'b0;
  assign \w2[9][7] [0] = 1'b0;
  assign \w2[9][8] [2] = 1'b0;
  assign \w2[9][9] [4] = 1'b0;
  assign \w2[9][9] [3] = 1'b0;
  assign \w2[9][9] [2] = 1'b0;
  assign \w2[9][9] [1] = 1'b0;
  assign \w2[9][10] [4] = 1'b0;
  assign \w2[9][10] [3] = 1'b0;
  assign \w2[9][10] [2] = 1'b0;
  assign \w2[9][10] [0] = 1'b0;
  assign \w2[9][11] [4] = 1'b0;
  assign \w2[9][11] [3] = 1'b0;
  assign \w2[9][11] [2] = 1'b0;
  assign \w2[9][11] [1] = 1'b0;
  assign \w2[9][11] [0] = 1'b0;
  assign \w2[9][12] [3] = 1'b0;
  assign \w2[9][13] [0] = 1'b0;
  assign \w2[9][14] [4] = 1'b0;
  assign \w2[9][14] [3] = 1'b0;
  assign \w2[9][14] [1] = 1'b0;
  assign \w2[9][15] [4] = 1'b0;
  assign \w2[9][15] [2] = 1'b0;
  assign \w2[9][15] [1] = 1'b0;
  assign \w2[9][16] [4] = 1'b0;
  assign \w2[9][16] [2] = 1'b0;
  assign \w2[9][16] [0] = 1'b0;
  assign \w2[9][17] [4] = 1'b0;
  assign \w2[9][17] [3] = 1'b0;
  assign \w2[9][17] [2] = 1'b0;
  assign \w2[9][18] [3] = 1'b0;
  assign \w2[9][19] [2] = 1'b0;
  assign \biases_l2[0] [3] = 1'b1;
  assign \biases_l2[0] [0] = 1'b1;
  assign \biases_l2[1] [3] = 1'b1;
  assign \biases_l2[1] [2] = 1'b1;
  assign \biases_l2[1] [0] = 1'b1;
  assign \biases_l2[2] [5] = 1'b1;
  assign \biases_l2[2] [4] = 1'b1;
  assign \biases_l2[2] [3] = 1'b1;
  assign \biases_l2[2] [2] = 1'b1;
  assign \biases_l2[2] [1] = 1'b1;
  assign \biases_l2[3] [5] = 1'b1;
  assign \biases_l2[3] [4] = 1'b1;
  assign \biases_l2[3] [3] = 1'b1;
  assign \biases_l2[3] [0] = 1'b1;
  assign \biases_l2[4] [5] = 1'b1;
  assign \biases_l2[4] [4] = 1'b1;
  assign \biases_l2[4] [0] = 1'b1;
  assign \biases_l2[5] [1] = 1'b1;
  assign \biases_l2[6] [5] = 1'b1;
  assign \biases_l2[6] [3] = 1'b1;
  assign \biases_l2[6] [2] = 1'b1;
  assign \biases_l2[6] [0] = 1'b1;
  assign \biases_l2[7] [5] = 1'b1;
  assign \biases_l2[7] [4] = 1'b1;
  assign \biases_l2[7] [2] = 1'b1;
  assign \biases_l2[7] [1] = 1'b1;
  assign \biases_l2[8] [5] = 1'b1;
  assign \biases_l2[8] [4] = 1'b1;
  assign \biases_l2[8] [0] = 1'b1;
  assign \biases_l2[9] [2] = 1'b1;
  assign \biases_l2[9] [1] = 1'b1;
  assign \w2[0][0] [4] = 1'b1;
  assign \w2[0][0] [3] = 1'b1;
  assign \w2[0][0] [2] = 1'b1;
  assign \w2[0][0] [1] = 1'b1;
  assign \w2[0][1] [1] = 1'b1;
  assign \w2[0][1] [0] = 1'b1;
  assign \w2[0][2] [4] = 1'b1;
  assign \w2[0][2] [3] = 1'b1;
  assign \w2[0][2] [2] = 1'b1;
  assign \w2[0][2] [0] = 1'b1;
  assign \w2[0][3] [4] = 1'b1;
  assign \w2[0][3] [3] = 1'b1;
  assign \w2[0][3] [2] = 1'b1;
  assign \w2[0][3] [0] = 1'b1;
  assign \w2[0][4] [4] = 1'b1;
  assign \w2[0][4] [3] = 1'b1;
  assign \w2[0][4] [1] = 1'b1;
  assign \w2[0][5] [4] = 1'b1;
  assign \w2[0][5] [3] = 1'b1;
  assign \w2[0][5] [2] = 1'b1;
  assign \w2[0][5] [0] = 1'b1;
  assign \w2[0][6] [0] = 1'b1;
  assign \w2[0][7] [4] = 1'b1;
  assign \w2[0][7] [3] = 1'b1;
  assign \w2[0][7] [2] = 1'b1;
  assign \w2[0][7] [1] = 1'b1;
  assign \w2[0][9] [4] = 1'b1;
  assign \w2[0][9] [2] = 1'b1;
  assign \w2[0][9] [1] = 1'b1;
  assign \w2[0][9] [0] = 1'b1;
  assign \w2[0][10] [4] = 1'b1;
  assign \w2[0][10] [3] = 1'b1;
  assign \w2[0][10] [2] = 1'b1;
  assign \w2[0][10] [1] = 1'b1;
  assign \w2[0][11] [4] = 1'b1;
  assign \w2[0][11] [3] = 1'b1;
  assign \w2[0][11] [2] = 1'b1;
  assign \w2[0][11] [1] = 1'b1;
  assign \w2[0][11] [0] = 1'b1;
  assign \w2[0][12] [0] = 1'b1;
  assign \w2[0][13] [0] = 1'b1;
  assign \w2[0][14] [1] = 1'b1;
  assign \w2[0][14] [0] = 1'b1;
  assign \w2[0][15] [1] = 1'b1;
  assign \w2[0][16] [4] = 1'b1;
  assign \w2[0][16] [3] = 1'b1;
  assign \w2[0][16] [2] = 1'b1;
  assign \w2[0][16] [1] = 1'b1;
  assign \w2[0][16] [0] = 1'b1;
  assign \w2[0][17] [4] = 1'b1;
  assign \w2[0][17] [3] = 1'b1;
  assign \w2[0][17] [2] = 1'b1;
  assign \w2[0][17] [0] = 1'b1;
  assign \w2[0][18] [2] = 1'b1;
  assign \w2[0][19] [4] = 1'b1;
  assign \w2[0][19] [3] = 1'b1;
  assign \w2[0][19] [1] = 1'b1;
  assign \w2[0][19] [0] = 1'b1;
  assign \w2[1][0] [2] = 1'b1;
  assign \w2[1][1] [4] = 1'b1;
  assign \w2[1][1] [3] = 1'b1;
  assign \w2[1][1] [2] = 1'b1;
  assign \w2[1][1] [0] = 1'b1;
  assign \w2[1][2] [3] = 1'b1;
  assign \w2[1][2] [0] = 1'b1;
  assign \w2[1][3] [2] = 1'b1;
  assign \w2[1][3] [0] = 1'b1;
  assign \w2[1][4] [2] = 1'b1;
  assign \w2[1][4] [0] = 1'b1;
  assign \w2[1][5] [3] = 1'b1;
  assign \w2[1][5] [1] = 1'b1;
  assign \w2[1][6] [4] = 1'b1;
  assign \w2[1][6] [2] = 1'b1;
  assign \w2[1][6] [1] = 1'b1;
  assign \w2[1][6] [0] = 1'b1;
  assign \w2[1][7] [4] = 1'b1;
  assign \w2[1][7] [3] = 1'b1;
  assign \w2[1][7] [2] = 1'b1;
  assign \w2[1][7] [1] = 1'b1;
  assign \w2[1][8] [4] = 1'b1;
  assign \w2[1][8] [3] = 1'b1;
  assign \w2[1][8] [2] = 1'b1;
  assign \w2[1][8] [1] = 1'b1;
  assign \w2[1][9] [4] = 1'b1;
  assign \w2[1][9] [3] = 1'b1;
  assign \w2[1][9] [2] = 1'b1;
  assign \w2[1][9] [1] = 1'b1;
  assign \w2[1][10] [2] = 1'b1;
  assign \w2[1][10] [0] = 1'b1;
  assign \w2[1][11] [4] = 1'b1;
  assign \w2[1][11] [2] = 1'b1;
  assign \w2[1][11] [1] = 1'b1;
  assign \w2[1][12] [2] = 1'b1;
  assign \w2[1][13] [4] = 1'b1;
  assign \w2[1][13] [3] = 1'b1;
  assign \w2[1][13] [1] = 1'b1;
  assign \w2[1][13] [0] = 1'b1;
  assign \w2[1][14] [4] = 1'b1;
  assign \w2[1][14] [1] = 1'b1;
  assign \w2[1][14] [0] = 1'b1;
  assign \w2[1][15] [2] = 1'b1;
  assign \w2[1][15] [1] = 1'b1;
  assign \w2[1][15] [0] = 1'b1;
  assign \w2[1][16] [2] = 1'b1;
  assign \w2[1][16] [1] = 1'b1;
  assign \w2[1][16] [0] = 1'b1;
  assign \w2[1][17] [4] = 1'b1;
  assign \w2[1][17] [3] = 1'b1;
  assign \w2[1][17] [2] = 1'b1;
  assign \w2[1][17] [0] = 1'b1;
  assign \w2[1][18] [1] = 1'b1;
  assign \w2[1][19] [4] = 1'b1;
  assign \w2[1][19] [3] = 1'b1;
  assign \w2[1][19] [2] = 1'b1;
  assign \w2[2][0] [4] = 1'b1;
  assign \w2[2][0] [3] = 1'b1;
  assign \w2[2][0] [1] = 1'b1;
  assign \w2[2][0] [0] = 1'b1;
  assign \w2[2][1] [4] = 1'b1;
  assign \w2[2][1] [3] = 1'b1;
  assign \w2[2][1] [2] = 1'b1;
  assign \w2[2][1] [1] = 1'b1;
  assign \w2[2][1] [0] = 1'b1;
  assign \w2[2][2] [4] = 1'b1;
  assign \w2[2][2] [3] = 1'b1;
  assign \w2[2][3] [4] = 1'b1;
  assign \w2[2][3] [3] = 1'b1;
  assign \w2[2][3] [2] = 1'b1;
  assign \w2[2][3] [1] = 1'b1;
  assign \w2[2][3] [0] = 1'b1;
  assign \w2[2][4] [1] = 1'b1;
  assign \w2[2][5] [4] = 1'b1;
  assign \w2[2][5] [3] = 1'b1;
  assign \w2[2][5] [2] = 1'b1;
  assign \w2[2][5] [1] = 1'b1;
  assign \w2[2][6] [4] = 1'b1;
  assign \w2[2][6] [3] = 1'b1;
  assign \w2[2][6] [1] = 1'b1;
  assign \w2[2][7] [4] = 1'b1;
  assign \w2[2][7] [3] = 1'b1;
  assign \w2[2][7] [2] = 1'b1;
  assign \w2[2][7] [1] = 1'b1;
  assign \w2[2][8] [2] = 1'b1;
  assign \w2[2][8] [0] = 1'b1;
  assign \w2[2][9] [4] = 1'b1;
  assign \w2[2][9] [3] = 1'b1;
  assign \w2[2][9] [2] = 1'b1;
  assign \w2[2][10] [2] = 1'b1;
  assign \w2[2][10] [0] = 1'b1;
  assign \w2[2][11] [4] = 1'b1;
  assign \w2[2][11] [2] = 1'b1;
  assign \w2[2][11] [0] = 1'b1;
  assign \w2[2][13] [2] = 1'b1;
  assign \w2[2][13] [1] = 1'b1;
  assign \w2[2][13] [0] = 1'b1;
  assign \w2[2][14] [0] = 1'b1;
  assign \w2[2][16] [3] = 1'b1;
  assign \w2[2][16] [1] = 1'b1;
  assign \w2[2][16] [0] = 1'b1;
  assign \w2[2][17] [2] = 1'b1;
  assign \w2[2][19] [0] = 1'b1;
  assign \w2[3][0] [0] = 1'b1;
  assign \w2[3][1] [4] = 1'b1;
  assign \w2[3][1] [3] = 1'b1;
  assign \w2[3][1] [2] = 1'b1;
  assign \w2[3][2] [4] = 1'b1;
  assign \w2[3][2] [3] = 1'b1;
  assign \w2[3][3] [4] = 1'b1;
  assign \w2[3][3] [3] = 1'b1;
  assign \w2[3][4] [1] = 1'b1;
  assign \w2[3][5] [1] = 1'b1;
  assign \w2[3][6] [4] = 1'b1;
  assign \w2[3][6] [3] = 1'b1;
  assign \w2[3][6] [2] = 1'b1;
  assign \w2[3][7] [1] = 1'b1;
  assign \w2[3][7] [0] = 1'b1;
  assign \w2[3][8] [4] = 1'b1;
  assign \w2[3][8] [2] = 1'b1;
  assign \w2[3][8] [1] = 1'b1;
  assign \w2[3][8] [0] = 1'b1;
  assign \w2[3][9] [1] = 1'b1;
  assign \w2[3][9] [0] = 1'b1;
  assign \w2[3][11] [1] = 1'b1;
  assign \w2[3][12] [4] = 1'b1;
  assign \w2[3][12] [3] = 1'b1;
  assign \w2[3][12] [2] = 1'b1;
  assign \w2[3][14] [2] = 1'b1;
  assign \w2[3][14] [0] = 1'b1;
  assign \w2[3][16] [0] = 1'b1;
  assign \w2[3][17] [2] = 1'b1;
  assign \w2[3][17] [0] = 1'b1;
  assign \w2[3][18] [2] = 1'b1;
  assign \w2[3][18] [1] = 1'b1;
  assign \w2[3][18] [0] = 1'b1;
  assign \w2[3][19] [2] = 1'b1;
  assign \w2[4][1] [1] = 1'b1;
  assign \w2[4][2] [3] = 1'b1;
  assign \w2[4][2] [1] = 1'b1;
  assign \w2[4][3] [4] = 1'b1;
  assign \w2[4][3] [3] = 1'b1;
  assign \w2[4][3] [2] = 1'b1;
  assign \w2[4][3] [0] = 1'b1;
  assign \w2[4][4] [2] = 1'b1;
  assign \w2[4][5] [1] = 1'b1;
  assign \w2[4][6] [2] = 1'b1;
  assign \w2[4][6] [0] = 1'b1;
  assign \w2[4][7] [4] = 1'b1;
  assign \w2[4][7] [3] = 1'b1;
  assign \w2[4][7] [2] = 1'b1;
  assign \w2[4][8] [0] = 1'b1;
  assign \w2[4][9] [4] = 1'b1;
  assign \w2[4][9] [3] = 1'b1;
  assign \w2[4][9] [2] = 1'b1;
  assign \w2[4][9] [1] = 1'b1;
  assign \w2[4][11] [2] = 1'b1;
  assign \w2[4][11] [0] = 1'b1;
  assign \w2[4][12] [4] = 1'b1;
  assign \w2[4][12] [3] = 1'b1;
  assign \w2[4][12] [0] = 1'b1;
  assign \w2[4][13] [0] = 1'b1;
  assign \w2[4][14] [4] = 1'b1;
  assign \w2[4][14] [3] = 1'b1;
  assign \w2[4][14] [2] = 1'b1;
  assign \w2[4][14] [1] = 1'b1;
  assign \w2[4][14] [0] = 1'b1;
  assign \w2[4][15] [1] = 1'b1;
  assign \w2[4][16] [4] = 1'b1;
  assign \w2[4][16] [3] = 1'b1;
  assign \w2[4][16] [2] = 1'b1;
  assign \w2[4][16] [1] = 1'b1;
  assign \w2[4][17] [4] = 1'b1;
  assign \w2[4][17] [3] = 1'b1;
  assign \w2[4][17] [2] = 1'b1;
  assign \w2[4][17] [1] = 1'b1;
  assign \w2[4][17] [0] = 1'b1;
  assign \w2[4][18] [4] = 1'b1;
  assign \w2[4][18] [3] = 1'b1;
  assign \w2[4][18] [2] = 1'b1;
  assign \w2[4][19] [1] = 1'b1;
  assign \w2[5][0] [3] = 1'b1;
  assign \w2[5][1] [1] = 1'b1;
  assign \w2[5][2] [0] = 1'b1;
  assign \w2[5][3] [4] = 1'b1;
  assign \w2[5][3] [3] = 1'b1;
  assign \w2[5][3] [2] = 1'b1;
  assign \w2[5][3] [1] = 1'b1;
  assign \w2[5][3] [0] = 1'b1;
  assign \w2[5][4] [4] = 1'b1;
  assign \w2[5][4] [3] = 1'b1;
  assign \w2[5][4] [2] = 1'b1;
  assign \w2[5][5] [4] = 1'b1;
  assign \w2[5][5] [3] = 1'b1;
  assign \w2[5][5] [2] = 1'b1;
  assign \w2[5][6] [1] = 1'b1;
  assign \w2[5][8] [4] = 1'b1;
  assign \w2[5][8] [3] = 1'b1;
  assign \w2[5][8] [2] = 1'b1;
  assign \w2[5][8] [1] = 1'b1;
  assign \w2[5][9] [4] = 1'b1;
  assign \w2[5][9] [3] = 1'b1;
  assign \w2[5][9] [2] = 1'b1;
  assign \w2[5][10] [2] = 1'b1;
  assign \w2[5][11] [4] = 1'b1;
  assign \w2[5][11] [3] = 1'b1;
  assign \w2[5][11] [2] = 1'b1;
  assign \w2[5][12] [4] = 1'b1;
  assign \w2[5][12] [3] = 1'b1;
  assign \w2[5][12] [2] = 1'b1;
  assign \w2[5][12] [0] = 1'b1;
  assign \w2[5][13] [4] = 1'b1;
  assign \w2[5][13] [3] = 1'b1;
  assign \w2[5][13] [2] = 1'b1;
  assign \w2[5][14] [1] = 1'b1;
  assign \w2[5][14] [0] = 1'b1;
  assign \w2[5][15] [2] = 1'b1;
  assign \w2[5][15] [1] = 1'b1;
  assign \w2[5][15] [0] = 1'b1;
  assign \w2[5][16] [4] = 1'b1;
  assign \w2[5][16] [3] = 1'b1;
  assign \w2[5][16] [2] = 1'b1;
  assign \w2[5][16] [1] = 1'b1;
  assign \w2[5][17] [4] = 1'b1;
  assign \w2[5][17] [2] = 1'b1;
  assign \w2[5][17] [1] = 1'b1;
  assign \w2[5][18] [4] = 1'b1;
  assign \w2[5][18] [3] = 1'b1;
  assign \w2[5][18] [2] = 1'b1;
  assign \w2[5][19] [2] = 1'b1;
  assign \w2[5][19] [1] = 1'b1;
  assign \w2[5][19] [0] = 1'b1;
  assign \w2[6][0] [1] = 1'b1;
  assign \w2[6][1] [3] = 1'b1;
  assign \w2[6][1] [0] = 1'b1;
  assign \w2[6][2] [4] = 1'b1;
  assign \w2[6][2] [2] = 1'b1;
  assign \w2[6][2] [1] = 1'b1;
  assign \w2[6][3] [0] = 1'b1;
  assign \w2[6][4] [0] = 1'b1;
  assign \w2[6][5] [4] = 1'b1;
  assign \w2[6][5] [2] = 1'b1;
  assign \w2[6][5] [1] = 1'b1;
  assign \w2[6][7] [1] = 1'b1;
  assign \w2[6][7] [0] = 1'b1;
  assign \w2[6][8] [1] = 1'b1;
  assign \w2[6][8] [0] = 1'b1;
  assign \w2[6][9] [4] = 1'b1;
  assign \w2[6][9] [3] = 1'b1;
  assign \w2[6][9] [2] = 1'b1;
  assign \w2[6][10] [4] = 1'b1;
  assign \w2[6][10] [2] = 1'b1;
  assign \w2[6][10] [1] = 1'b1;
  assign \w2[6][10] [0] = 1'b1;
  assign \w2[6][11] [2] = 1'b1;
  assign \w2[6][11] [1] = 1'b1;
  assign \w2[6][12] [4] = 1'b1;
  assign \w2[6][12] [3] = 1'b1;
  assign \w2[6][12] [0] = 1'b1;
  assign \w2[6][13] [1] = 1'b1;
  assign \w2[6][13] [0] = 1'b1;
  assign \w2[6][14] [4] = 1'b1;
  assign \w2[6][14] [3] = 1'b1;
  assign \w2[6][14] [2] = 1'b1;
  assign \w2[6][15] [4] = 1'b1;
  assign \w2[6][15] [1] = 1'b1;
  assign \w2[6][15] [0] = 1'b1;
  assign \w2[6][16] [4] = 1'b1;
  assign \w2[6][16] [3] = 1'b1;
  assign \w2[6][16] [2] = 1'b1;
  assign \w2[6][16] [1] = 1'b1;
  assign \w2[6][16] [0] = 1'b1;
  assign \w2[6][17] [4] = 1'b1;
  assign \w2[6][17] [3] = 1'b1;
  assign \w2[6][17] [2] = 1'b1;
  assign \w2[6][17] [1] = 1'b1;
  assign \w2[6][18] [0] = 1'b1;
  assign \w2[6][19] [0] = 1'b1;
  assign \w2[7][1] [3] = 1'b1;
  assign \w2[7][1] [0] = 1'b1;
  assign \w2[7][2] [4] = 1'b1;
  assign \w2[7][2] [3] = 1'b1;
  assign \w2[7][2] [2] = 1'b1;
  assign \w2[7][2] [1] = 1'b1;
  assign \w2[7][2] [0] = 1'b1;
  assign \w2[7][3] [4] = 1'b1;
  assign \w2[7][3] [2] = 1'b1;
  assign \w2[7][3] [1] = 1'b1;
  assign \w2[7][3] [0] = 1'b1;
  assign \w2[7][4] [4] = 1'b1;
  assign \w2[7][4] [3] = 1'b1;
  assign \w2[7][4] [0] = 1'b1;
  assign \w2[7][5] [4] = 1'b1;
  assign \w2[7][5] [3] = 1'b1;
  assign \w2[7][5] [0] = 1'b1;
  assign \w2[7][6] [4] = 1'b1;
  assign \w2[7][6] [3] = 1'b1;
  assign \w2[7][6] [1] = 1'b1;
  assign \w2[7][7] [4] = 1'b1;
  assign \w2[7][7] [3] = 1'b1;
  assign \w2[7][7] [2] = 1'b1;
  assign \w2[7][7] [1] = 1'b1;
  assign \w2[7][7] [0] = 1'b1;
  assign \w2[7][8] [2] = 1'b1;
  assign \w2[7][8] [0] = 1'b1;
  assign \w2[7][9] [3] = 1'b1;
  assign \w2[7][9] [0] = 1'b1;
  assign \w2[7][11] [4] = 1'b1;
  assign \w2[7][11] [3] = 1'b1;
  assign \w2[7][11] [2] = 1'b1;
  assign \w2[7][11] [1] = 1'b1;
  assign \w2[7][12] [2] = 1'b1;
  assign \w2[7][12] [1] = 1'b1;
  assign \w2[7][14] [0] = 1'b1;
  assign \w2[7][15] [4] = 1'b1;
  assign \w2[7][15] [2] = 1'b1;
  assign \w2[7][15] [1] = 1'b1;
  assign \w2[7][15] [0] = 1'b1;
  assign \w2[7][16] [2] = 1'b1;
  assign \w2[7][17] [4] = 1'b1;
  assign \w2[7][17] [2] = 1'b1;
  assign \w2[7][17] [1] = 1'b1;
  assign \w2[7][17] [0] = 1'b1;
  assign \w2[7][18] [1] = 1'b1;
  assign \w2[7][18] [0] = 1'b1;
  assign \w2[8][0] [4] = 1'b1;
  assign \w2[8][0] [3] = 1'b1;
  assign \w2[8][0] [0] = 1'b1;
  assign \w2[8][1] [2] = 1'b1;
  assign \w2[8][2] [4] = 1'b1;
  assign \w2[8][2] [3] = 1'b1;
  assign \w2[8][2] [2] = 1'b1;
  assign \w2[8][3] [1] = 1'b1;
  assign \w2[8][5] [0] = 1'b1;
  assign \w2[8][6] [1] = 1'b1;
  assign \w2[8][7] [3] = 1'b1;
  assign \w2[8][7] [1] = 1'b1;
  assign \w2[8][8] [1] = 1'b1;
  assign \w2[8][8] [0] = 1'b1;
  assign \w2[8][9] [0] = 1'b1;
  assign \w2[8][11] [4] = 1'b1;
  assign \w2[8][11] [2] = 1'b1;
  assign \w2[8][13] [1] = 1'b1;
  assign \w2[8][14] [4] = 1'b1;
  assign \w2[8][14] [3] = 1'b1;
  assign \w2[8][14] [2] = 1'b1;
  assign \w2[8][14] [0] = 1'b1;
  assign \w2[8][15] [2] = 1'b1;
  assign \w2[8][15] [1] = 1'b1;
  assign \w2[8][16] [4] = 1'b1;
  assign \w2[8][16] [3] = 1'b1;
  assign \w2[8][16] [2] = 1'b1;
  assign \w2[8][16] [1] = 1'b1;
  assign \w2[8][16] [0] = 1'b1;
  assign \w2[8][17] [4] = 1'b1;
  assign \w2[8][17] [3] = 1'b1;
  assign \w2[8][17] [2] = 1'b1;
  assign \w2[8][17] [1] = 1'b1;
  assign \w2[8][17] [0] = 1'b1;
  assign \w2[8][18] [4] = 1'b1;
  assign \w2[8][18] [3] = 1'b1;
  assign \w2[8][18] [1] = 1'b1;
  assign \w2[8][19] [4] = 1'b1;
  assign \w2[8][19] [1] = 1'b1;
  assign \w2[8][19] [0] = 1'b1;
  assign \w2[9][0] [4] = 1'b1;
  assign \w2[9][0] [3] = 1'b1;
  assign \w2[9][1] [2] = 1'b1;
  assign \w2[9][1] [1] = 1'b1;
  assign \w2[9][2] [4] = 1'b1;
  assign \w2[9][2] [2] = 1'b1;
  assign \w2[9][2] [1] = 1'b1;
  assign \w2[9][2] [0] = 1'b1;
  assign \w2[9][3] [3] = 1'b1;
  assign \w2[9][3] [0] = 1'b1;
  assign \w2[9][4] [4] = 1'b1;
  assign \w2[9][4] [2] = 1'b1;
  assign \w2[9][4] [1] = 1'b1;
  assign \w2[9][4] [0] = 1'b1;
  assign \w2[9][5] [4] = 1'b1;
  assign \w2[9][5] [3] = 1'b1;
  assign \w2[9][5] [2] = 1'b1;
  assign \w2[9][5] [1] = 1'b1;
  assign \w2[9][5] [0] = 1'b1;
  assign \w2[9][6] [2] = 1'b1;
  assign \w2[9][7] [4] = 1'b1;
  assign \w2[9][7] [3] = 1'b1;
  assign \w2[9][7] [2] = 1'b1;
  assign \w2[9][8] [4] = 1'b1;
  assign \w2[9][8] [3] = 1'b1;
  assign \w2[9][8] [1] = 1'b1;
  assign \w2[9][8] [0] = 1'b1;
  assign \w2[9][9] [0] = 1'b1;
  assign \w2[9][10] [1] = 1'b1;
  assign \w2[9][12] [4] = 1'b1;
  assign \w2[9][12] [2] = 1'b1;
  assign \w2[9][12] [1] = 1'b1;
  assign \w2[9][12] [0] = 1'b1;
  assign \w2[9][13] [4] = 1'b1;
  assign \w2[9][13] [3] = 1'b1;
  assign \w2[9][13] [2] = 1'b1;
  assign \w2[9][13] [1] = 1'b1;
  assign \w2[9][14] [2] = 1'b1;
  assign \w2[9][14] [0] = 1'b1;
  assign \w2[9][15] [3] = 1'b1;
  assign \w2[9][15] [0] = 1'b1;
  assign \w2[9][16] [3] = 1'b1;
  assign \w2[9][16] [1] = 1'b1;
  assign \w2[9][17] [1] = 1'b1;
  assign \w2[9][17] [0] = 1'b1;
  assign \w2[9][18] [4] = 1'b1;
  assign \w2[9][18] [2] = 1'b1;
  assign \w2[9][18] [1] = 1'b1;
  assign \w2[9][18] [0] = 1'b1;
  assign \w2[9][19] [4] = 1'b1;
  assign \w2[9][19] [3] = 1'b1;
  assign \w2[9][19] [1] = 1'b1;
  assign \w2[9][19] [0] = 1'b1;
  _HDFF_verplex \out_reg_reg[0][17] (.Q(\out_reg[0] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[0] [17]));
  _HDFF_verplex \out_reg_reg[0][16] (.Q(\out_reg[0] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[0] [16]));
  _HDFF_verplex \out_reg_reg[0][15] (.Q(\out_reg[0] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[0] [15]));
  _HDFF_verplex \out_reg_reg[0][14] (.Q(\out_reg[0] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[0] [14]));
  _HDFF_verplex \out_reg_reg[0][13] (.Q(\out_reg[0] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[0] [13]));
  _HDFF_verplex \out_reg_reg[0][12] (.Q(\out_reg[0] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[0] [12]));
  _HDFF_verplex \out_reg_reg[0][11] (.Q(\out_reg[0] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[0] [11]));
  _HDFF_verplex \out_reg_reg[0][10] (.Q(\out_reg[0] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[0] [10]));
  _HDFF_verplex \out_reg_reg[0][9] (.Q(\out_reg[0] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[0] [9]));
  _HDFF_verplex \out_reg_reg[0][8] (.Q(\out_reg[0] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[0] [8]));
  _HDFF_verplex \out_reg_reg[0][7] (.Q(\out_reg[0] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[0] [7]));
  _HDFF_verplex \out_reg_reg[0][6] (.Q(\out_reg[0] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[0] [6]));
  _HDFF_verplex \out_reg_reg[0][5] (.Q(\out_reg[0] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[0] [5]));
  _HDFF_verplex \out_reg_reg[0][4] (.Q(\out_reg[0] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[0] [4]));
  _HDFF_verplex \out_reg_reg[0][3] (.Q(\out_reg[0] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[0] [3]));
  _HDFF_verplex \out_reg_reg[0][2] (.Q(\out_reg[0] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[0] [2]));
  _HDFF_verplex \out_reg_reg[0][1] (.Q(\out_reg[0] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[0] [1]));
  _HDFF_verplex \out_reg_reg[0][0] (.Q(\out_reg[0] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[0] [0]));
  _HDFF_verplex \out_reg_reg[1][17] (.Q(\out_reg[1] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[1] [17]));
  _HDFF_verplex \out_reg_reg[1][16] (.Q(\out_reg[1] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[1] [16]));
  _HDFF_verplex \out_reg_reg[1][15] (.Q(\out_reg[1] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[1] [15]));
  _HDFF_verplex \out_reg_reg[1][14] (.Q(\out_reg[1] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[1] [14]));
  _HDFF_verplex \out_reg_reg[1][13] (.Q(\out_reg[1] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[1] [13]));
  _HDFF_verplex \out_reg_reg[1][12] (.Q(\out_reg[1] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[1] [12]));
  _HDFF_verplex \out_reg_reg[1][11] (.Q(\out_reg[1] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[1] [11]));
  _HDFF_verplex \out_reg_reg[1][10] (.Q(\out_reg[1] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[1] [10]));
  _HDFF_verplex \out_reg_reg[1][9] (.Q(\out_reg[1] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[1] [9]));
  _HDFF_verplex \out_reg_reg[1][8] (.Q(\out_reg[1] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[1] [8]));
  _HDFF_verplex \out_reg_reg[1][7] (.Q(\out_reg[1] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[1] [7]));
  _HDFF_verplex \out_reg_reg[1][6] (.Q(\out_reg[1] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[1] [6]));
  _HDFF_verplex \out_reg_reg[1][5] (.Q(\out_reg[1] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[1] [5]));
  _HDFF_verplex \out_reg_reg[1][4] (.Q(\out_reg[1] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[1] [4]));
  _HDFF_verplex \out_reg_reg[1][3] (.Q(\out_reg[1] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[1] [3]));
  _HDFF_verplex \out_reg_reg[1][2] (.Q(\out_reg[1] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[1] [2]));
  _HDFF_verplex \out_reg_reg[1][1] (.Q(\out_reg[1] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[1] [1]));
  _HDFF_verplex \out_reg_reg[1][0] (.Q(\out_reg[1] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[1] [0]));
  _HDFF_verplex \out_reg_reg[2][17] (.Q(\out_reg[2] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[2] [17]));
  _HDFF_verplex \out_reg_reg[2][16] (.Q(\out_reg[2] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[2] [16]));
  _HDFF_verplex \out_reg_reg[2][15] (.Q(\out_reg[2] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[2] [15]));
  _HDFF_verplex \out_reg_reg[2][14] (.Q(\out_reg[2] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[2] [14]));
  _HDFF_verplex \out_reg_reg[2][13] (.Q(\out_reg[2] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[2] [13]));
  _HDFF_verplex \out_reg_reg[2][12] (.Q(\out_reg[2] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[2] [12]));
  _HDFF_verplex \out_reg_reg[2][11] (.Q(\out_reg[2] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[2] [11]));
  _HDFF_verplex \out_reg_reg[2][10] (.Q(\out_reg[2] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[2] [10]));
  _HDFF_verplex \out_reg_reg[2][9] (.Q(\out_reg[2] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[2] [9]));
  _HDFF_verplex \out_reg_reg[2][8] (.Q(\out_reg[2] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[2] [8]));
  _HDFF_verplex \out_reg_reg[2][7] (.Q(\out_reg[2] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[2] [7]));
  _HDFF_verplex \out_reg_reg[2][6] (.Q(\out_reg[2] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[2] [6]));
  _HDFF_verplex \out_reg_reg[2][5] (.Q(\out_reg[2] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[2] [5]));
  _HDFF_verplex \out_reg_reg[2][4] (.Q(\out_reg[2] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[2] [4]));
  _HDFF_verplex \out_reg_reg[2][3] (.Q(\out_reg[2] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[2] [3]));
  _HDFF_verplex \out_reg_reg[2][2] (.Q(\out_reg[2] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[2] [2]));
  _HDFF_verplex \out_reg_reg[2][1] (.Q(\out_reg[2] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[2] [1]));
  _HDFF_verplex \out_reg_reg[2][0] (.Q(\out_reg[2] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[2] [0]));
  _HDFF_verplex \out_reg_reg[3][17] (.Q(\out_reg[3] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[3] [17]));
  _HDFF_verplex \out_reg_reg[3][16] (.Q(\out_reg[3] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[3] [16]));
  _HDFF_verplex \out_reg_reg[3][15] (.Q(\out_reg[3] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[3] [15]));
  _HDFF_verplex \out_reg_reg[3][14] (.Q(\out_reg[3] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[3] [14]));
  _HDFF_verplex \out_reg_reg[3][13] (.Q(\out_reg[3] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[3] [13]));
  _HDFF_verplex \out_reg_reg[3][12] (.Q(\out_reg[3] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[3] [12]));
  _HDFF_verplex \out_reg_reg[3][11] (.Q(\out_reg[3] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[3] [11]));
  _HDFF_verplex \out_reg_reg[3][10] (.Q(\out_reg[3] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[3] [10]));
  _HDFF_verplex \out_reg_reg[3][9] (.Q(\out_reg[3] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[3] [9]));
  _HDFF_verplex \out_reg_reg[3][8] (.Q(\out_reg[3] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[3] [8]));
  _HDFF_verplex \out_reg_reg[3][7] (.Q(\out_reg[3] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[3] [7]));
  _HDFF_verplex \out_reg_reg[3][6] (.Q(\out_reg[3] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[3] [6]));
  _HDFF_verplex \out_reg_reg[3][5] (.Q(\out_reg[3] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[3] [5]));
  _HDFF_verplex \out_reg_reg[3][4] (.Q(\out_reg[3] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[3] [4]));
  _HDFF_verplex \out_reg_reg[3][3] (.Q(\out_reg[3] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[3] [3]));
  _HDFF_verplex \out_reg_reg[3][2] (.Q(\out_reg[3] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[3] [2]));
  _HDFF_verplex \out_reg_reg[3][1] (.Q(\out_reg[3] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[3] [1]));
  _HDFF_verplex \out_reg_reg[3][0] (.Q(\out_reg[3] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[3] [0]));
  _HDFF_verplex \out_reg_reg[4][17] (.Q(\out_reg[4] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[4] [17]));
  _HDFF_verplex \out_reg_reg[4][16] (.Q(\out_reg[4] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[4] [16]));
  _HDFF_verplex \out_reg_reg[4][15] (.Q(\out_reg[4] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[4] [15]));
  _HDFF_verplex \out_reg_reg[4][14] (.Q(\out_reg[4] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[4] [14]));
  _HDFF_verplex \out_reg_reg[4][13] (.Q(\out_reg[4] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[4] [13]));
  _HDFF_verplex \out_reg_reg[4][12] (.Q(\out_reg[4] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[4] [12]));
  _HDFF_verplex \out_reg_reg[4][11] (.Q(\out_reg[4] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[4] [11]));
  _HDFF_verplex \out_reg_reg[4][10] (.Q(\out_reg[4] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[4] [10]));
  _HDFF_verplex \out_reg_reg[4][9] (.Q(\out_reg[4] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[4] [9]));
  _HDFF_verplex \out_reg_reg[4][8] (.Q(\out_reg[4] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[4] [8]));
  _HDFF_verplex \out_reg_reg[4][7] (.Q(\out_reg[4] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[4] [7]));
  _HDFF_verplex \out_reg_reg[4][6] (.Q(\out_reg[4] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[4] [6]));
  _HDFF_verplex \out_reg_reg[4][5] (.Q(\out_reg[4] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[4] [5]));
  _HDFF_verplex \out_reg_reg[4][4] (.Q(\out_reg[4] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[4] [4]));
  _HDFF_verplex \out_reg_reg[4][3] (.Q(\out_reg[4] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[4] [3]));
  _HDFF_verplex \out_reg_reg[4][2] (.Q(\out_reg[4] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[4] [2]));
  _HDFF_verplex \out_reg_reg[4][1] (.Q(\out_reg[4] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[4] [1]));
  _HDFF_verplex \out_reg_reg[4][0] (.Q(\out_reg[4] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[4] [0]));
  _HDFF_verplex \out_reg_reg[5][17] (.Q(\out_reg[5] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[5] [17]));
  _HDFF_verplex \out_reg_reg[5][16] (.Q(\out_reg[5] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[5] [16]));
  _HDFF_verplex \out_reg_reg[5][15] (.Q(\out_reg[5] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[5] [15]));
  _HDFF_verplex \out_reg_reg[5][14] (.Q(\out_reg[5] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[5] [14]));
  _HDFF_verplex \out_reg_reg[5][13] (.Q(\out_reg[5] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[5] [13]));
  _HDFF_verplex \out_reg_reg[5][12] (.Q(\out_reg[5] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[5] [12]));
  _HDFF_verplex \out_reg_reg[5][11] (.Q(\out_reg[5] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[5] [11]));
  _HDFF_verplex \out_reg_reg[5][10] (.Q(\out_reg[5] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[5] [10]));
  _HDFF_verplex \out_reg_reg[5][9] (.Q(\out_reg[5] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[5] [9]));
  _HDFF_verplex \out_reg_reg[5][8] (.Q(\out_reg[5] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[5] [8]));
  _HDFF_verplex \out_reg_reg[5][7] (.Q(\out_reg[5] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[5] [7]));
  _HDFF_verplex \out_reg_reg[5][6] (.Q(\out_reg[5] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[5] [6]));
  _HDFF_verplex \out_reg_reg[5][5] (.Q(\out_reg[5] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[5] [5]));
  _HDFF_verplex \out_reg_reg[5][4] (.Q(\out_reg[5] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[5] [4]));
  _HDFF_verplex \out_reg_reg[5][3] (.Q(\out_reg[5] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[5] [3]));
  _HDFF_verplex \out_reg_reg[5][2] (.Q(\out_reg[5] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[5] [2]));
  _HDFF_verplex \out_reg_reg[5][1] (.Q(\out_reg[5] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[5] [1]));
  _HDFF_verplex \out_reg_reg[5][0] (.Q(\out_reg[5] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[5] [0]));
  _HDFF_verplex \out_reg_reg[6][17] (.Q(\out_reg[6] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[6] [17]));
  _HDFF_verplex \out_reg_reg[6][16] (.Q(\out_reg[6] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[6] [16]));
  _HDFF_verplex \out_reg_reg[6][15] (.Q(\out_reg[6] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[6] [15]));
  _HDFF_verplex \out_reg_reg[6][14] (.Q(\out_reg[6] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[6] [14]));
  _HDFF_verplex \out_reg_reg[6][13] (.Q(\out_reg[6] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[6] [13]));
  _HDFF_verplex \out_reg_reg[6][12] (.Q(\out_reg[6] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[6] [12]));
  _HDFF_verplex \out_reg_reg[6][11] (.Q(\out_reg[6] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[6] [11]));
  _HDFF_verplex \out_reg_reg[6][10] (.Q(\out_reg[6] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[6] [10]));
  _HDFF_verplex \out_reg_reg[6][9] (.Q(\out_reg[6] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[6] [9]));
  _HDFF_verplex \out_reg_reg[6][8] (.Q(\out_reg[6] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[6] [8]));
  _HDFF_verplex \out_reg_reg[6][7] (.Q(\out_reg[6] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[6] [7]));
  _HDFF_verplex \out_reg_reg[6][6] (.Q(\out_reg[6] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[6] [6]));
  _HDFF_verplex \out_reg_reg[6][5] (.Q(\out_reg[6] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[6] [5]));
  _HDFF_verplex \out_reg_reg[6][4] (.Q(\out_reg[6] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[6] [4]));
  _HDFF_verplex \out_reg_reg[6][3] (.Q(\out_reg[6] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[6] [3]));
  _HDFF_verplex \out_reg_reg[6][2] (.Q(\out_reg[6] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[6] [2]));
  _HDFF_verplex \out_reg_reg[6][1] (.Q(\out_reg[6] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[6] [1]));
  _HDFF_verplex \out_reg_reg[6][0] (.Q(\out_reg[6] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[6] [0]));
  _HDFF_verplex \out_reg_reg[7][17] (.Q(\out_reg[7] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[7] [17]));
  _HDFF_verplex \out_reg_reg[7][16] (.Q(\out_reg[7] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[7] [16]));
  _HDFF_verplex \out_reg_reg[7][15] (.Q(\out_reg[7] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[7] [15]));
  _HDFF_verplex \out_reg_reg[7][14] (.Q(\out_reg[7] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[7] [14]));
  _HDFF_verplex \out_reg_reg[7][13] (.Q(\out_reg[7] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[7] [13]));
  _HDFF_verplex \out_reg_reg[7][12] (.Q(\out_reg[7] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[7] [12]));
  _HDFF_verplex \out_reg_reg[7][11] (.Q(\out_reg[7] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[7] [11]));
  _HDFF_verplex \out_reg_reg[7][10] (.Q(\out_reg[7] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[7] [10]));
  _HDFF_verplex \out_reg_reg[7][9] (.Q(\out_reg[7] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[7] [9]));
  _HDFF_verplex \out_reg_reg[7][8] (.Q(\out_reg[7] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[7] [8]));
  _HDFF_verplex \out_reg_reg[7][7] (.Q(\out_reg[7] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[7] [7]));
  _HDFF_verplex \out_reg_reg[7][6] (.Q(\out_reg[7] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[7] [6]));
  _HDFF_verplex \out_reg_reg[7][5] (.Q(\out_reg[7] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[7] [5]));
  _HDFF_verplex \out_reg_reg[7][4] (.Q(\out_reg[7] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[7] [4]));
  _HDFF_verplex \out_reg_reg[7][3] (.Q(\out_reg[7] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[7] [3]));
  _HDFF_verplex \out_reg_reg[7][2] (.Q(\out_reg[7] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[7] [2]));
  _HDFF_verplex \out_reg_reg[7][1] (.Q(\out_reg[7] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[7] [1]));
  _HDFF_verplex \out_reg_reg[7][0] (.Q(\out_reg[7] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[7] [0]));
  _HDFF_verplex \out_reg_reg[8][17] (.Q(\out_reg[8] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[8] [17]));
  _HDFF_verplex \out_reg_reg[8][16] (.Q(\out_reg[8] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[8] [16]));
  _HDFF_verplex \out_reg_reg[8][15] (.Q(\out_reg[8] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[8] [15]));
  _HDFF_verplex \out_reg_reg[8][14] (.Q(\out_reg[8] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[8] [14]));
  _HDFF_verplex \out_reg_reg[8][13] (.Q(\out_reg[8] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[8] [13]));
  _HDFF_verplex \out_reg_reg[8][12] (.Q(\out_reg[8] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[8] [12]));
  _HDFF_verplex \out_reg_reg[8][11] (.Q(\out_reg[8] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[8] [11]));
  _HDFF_verplex \out_reg_reg[8][10] (.Q(\out_reg[8] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[8] [10]));
  _HDFF_verplex \out_reg_reg[8][9] (.Q(\out_reg[8] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[8] [9]));
  _HDFF_verplex \out_reg_reg[8][8] (.Q(\out_reg[8] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[8] [8]));
  _HDFF_verplex \out_reg_reg[8][7] (.Q(\out_reg[8] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[8] [7]));
  _HDFF_verplex \out_reg_reg[8][6] (.Q(\out_reg[8] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[8] [6]));
  _HDFF_verplex \out_reg_reg[8][5] (.Q(\out_reg[8] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[8] [5]));
  _HDFF_verplex \out_reg_reg[8][4] (.Q(\out_reg[8] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[8] [4]));
  _HDFF_verplex \out_reg_reg[8][3] (.Q(\out_reg[8] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[8] [3]));
  _HDFF_verplex \out_reg_reg[8][2] (.Q(\out_reg[8] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[8] [2]));
  _HDFF_verplex \out_reg_reg[8][1] (.Q(\out_reg[8] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[8] [1]));
  _HDFF_verplex \out_reg_reg[8][0] (.Q(\out_reg[8] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[8] [0]));
  _HDFF_verplex \out_reg_reg[9][17] (.Q(\out_reg[9] [17]), .QN( ), .S(N$18), .R(
    n5835), .CK(clk), .D(\row_output[9] [17]));
  _HDFF_verplex \out_reg_reg[9][16] (.Q(\out_reg[9] [16]), .QN( ), .S(N$17), .R(
    n5835), .CK(clk), .D(\row_output[9] [16]));
  _HDFF_verplex \out_reg_reg[9][15] (.Q(\out_reg[9] [15]), .QN( ), .S(N$16), .R(
    n5835), .CK(clk), .D(\row_output[9] [15]));
  _HDFF_verplex \out_reg_reg[9][14] (.Q(\out_reg[9] [14]), .QN( ), .S(N$15), .R(
    n5835), .CK(clk), .D(\row_output[9] [14]));
  _HDFF_verplex \out_reg_reg[9][13] (.Q(\out_reg[9] [13]), .QN( ), .S(N$14), .R(
    n5835), .CK(clk), .D(\row_output[9] [13]));
  _HDFF_verplex \out_reg_reg[9][12] (.Q(\out_reg[9] [12]), .QN( ), .S(N$13), .R(
    n5835), .CK(clk), .D(\row_output[9] [12]));
  _HDFF_verplex \out_reg_reg[9][11] (.Q(\out_reg[9] [11]), .QN( ), .S(N$12), .R(
    n5835), .CK(clk), .D(\row_output[9] [11]));
  _HDFF_verplex \out_reg_reg[9][10] (.Q(\out_reg[9] [10]), .QN( ), .S(N$11), .R(
    n5835), .CK(clk), .D(\row_output[9] [10]));
  _HDFF_verplex \out_reg_reg[9][9] (.Q(\out_reg[9] [9]), .QN( ), .S(N$10), .R(
    n5835), .CK(clk), .D(\row_output[9] [9]));
  _HDFF_verplex \out_reg_reg[9][8] (.Q(\out_reg[9] [8]), .QN( ), .S(N$9), .R(
    n5835), .CK(clk), .D(\row_output[9] [8]));
  _HDFF_verplex \out_reg_reg[9][7] (.Q(\out_reg[9] [7]), .QN( ), .S(N$8), .R(
    n5835), .CK(clk), .D(\row_output[9] [7]));
  _HDFF_verplex \out_reg_reg[9][6] (.Q(\out_reg[9] [6]), .QN( ), .S(N$7), .R(
    n5835), .CK(clk), .D(\row_output[9] [6]));
  _HDFF_verplex \out_reg_reg[9][5] (.Q(\out_reg[9] [5]), .QN( ), .S(N$6), .R(
    n5835), .CK(clk), .D(\row_output[9] [5]));
  _HDFF_verplex \out_reg_reg[9][4] (.Q(\out_reg[9] [4]), .QN( ), .S(N$5), .R(
    n5835), .CK(clk), .D(\row_output[9] [4]));
  _HDFF_verplex \out_reg_reg[9][3] (.Q(\out_reg[9] [3]), .QN( ), .S(N$4), .R(
    n5835), .CK(clk), .D(\row_output[9] [3]));
  _HDFF_verplex \out_reg_reg[9][2] (.Q(\out_reg[9] [2]), .QN( ), .S(N$3), .R(
    n5835), .CK(clk), .D(\row_output[9] [2]));
  _HDFF_verplex \out_reg_reg[9][1] (.Q(\out_reg[9] [1]), .QN( ), .S(N$2), .R(
    n5835), .CK(clk), .D(\row_output[9] [1]));
  _HDFF_verplex \out_reg_reg[9][0] (.Q(\out_reg[9] [0]), .QN( ), .S(N$1), .R(
    n5835), .CK(clk), .D(\row_output[9] [0]));
  not U$1(n5835, rst_n);
  VDW_ADD_19_1_0 add_5823_68_I1(.SUM({ \row_sums[0] [18:0] }), .A({ n5823_19[18:0] }), .B({\b2_extended[0] [13], 
    \b2_extended[0] [13], \b2_extended[0] [13], \b2_extended[0] [13], 
    \b2_extended[0] [13],  \b2_extended[0] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I1(.SUM({ n5823_19[18:0] }), .A({ n5822_30[18:0] }), .B({\prod_terms[0][19] [13], 
    \prod_terms[0][19] [13], \prod_terms[0][19] [13], \prod_terms[0][19] [13], 
    \prod_terms[0][19] [13],  \prod_terms[0][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I1(.SUM({ n5822_30[18:0] }), .A({ n5822_29[18:0] }), .B({\prod_terms[0][18] [13], 
    \prod_terms[0][18] [13], \prod_terms[0][18] [13], \prod_terms[0][18] [13], 
    \prod_terms[0][18] [13],  \prod_terms[0][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I1(.SUM({ n5822_29[18:0] }), .A({ n5822_28[18:0] }), .B({\prod_terms[0][17] [13], 
    \prod_terms[0][17] [13], \prod_terms[0][17] [13], \prod_terms[0][17] [13], 
    \prod_terms[0][17] [13],  \prod_terms[0][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I1(.SUM({ n5822_28[18:0] }), .A({ n5821_30[18:0] }), .B({\prod_terms[0][16] [13], 
    \prod_terms[0][16] [13], \prod_terms[0][16] [13], \prod_terms[0][16] [13], 
    \prod_terms[0][16] [13],  \prod_terms[0][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I1(.SUM({ n5821_30[18:0] }), .A({ n5821_29[18:0] }), .B({\prod_terms[0][15] [13], 
    \prod_terms[0][15] [13], \prod_terms[0][15] [13], \prod_terms[0][15] [13], 
    \prod_terms[0][15] [13],  \prod_terms[0][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I1(.SUM({ n5821_29[18:0] }), .A({ n5821_28[18:0] }), .B({\prod_terms[0][14] [13], 
    \prod_terms[0][14] [13], \prod_terms[0][14] [13], \prod_terms[0][14] [13], 
    \prod_terms[0][14] [13],  \prod_terms[0][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I1(.SUM({ n5821_28[18:0] }), .A({ n5820_30[18:0] }), .B({\prod_terms[0][13] [13], 
    \prod_terms[0][13] [13], \prod_terms[0][13] [13], \prod_terms[0][13] [13], 
    \prod_terms[0][13] [13],  \prod_terms[0][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I1(.SUM({ n5820_30[18:0] }), .A({ n5820_29[18:0] }), .B({\prod_terms[0][12] [13], 
    \prod_terms[0][12] [13], \prod_terms[0][12] [13], \prod_terms[0][12] [13], 
    \prod_terms[0][12] [13],  \prod_terms[0][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I1(.SUM({ n5820_29[18:0] }), .A({ n5820_28[18:0] }), .B({\prod_terms[0][11] [13], 
    \prod_terms[0][11] [13], \prod_terms[0][11] [13], \prod_terms[0][11] [13], 
    \prod_terms[0][11] [13],  \prod_terms[0][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I1(.SUM({ n5820_28[18:0] }), .A({ n5819_30[18:0] }), .B({\prod_terms[0][10] [13], 
    \prod_terms[0][10] [13], \prod_terms[0][10] [13], \prod_terms[0][10] [13], 
    \prod_terms[0][10] [13],  \prod_terms[0][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I1(.SUM({ n5819_30[18:0] }), .A({ n5819_29[18:0] }), .B({\prod_terms[0][9] [13], 
    \prod_terms[0][9] [13], \prod_terms[0][9] [13], \prod_terms[0][9] [13], 
    \prod_terms[0][9] [13],  \prod_terms[0][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I1(.SUM({ n5819_29[18:0] }), .A({ n5819_28[18:0] }), .B({\prod_terms[0][8] [13], 
    \prod_terms[0][8] [13], \prod_terms[0][8] [13], \prod_terms[0][8] [13], 
    \prod_terms[0][8] [13],  \prod_terms[0][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I1(.SUM({ n5819_28[18:0] }), .A({ n5818_30[18:0] }), .B({\prod_terms[0][7] [13], 
    \prod_terms[0][7] [13], \prod_terms[0][7] [13], \prod_terms[0][7] [13], 
    \prod_terms[0][7] [13],  \prod_terms[0][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I1(.SUM({ n5818_30[18:0] }), .A({ n5818_29[18:0] }), .B({\prod_terms[0][6] [13], 
    \prod_terms[0][6] [13], \prod_terms[0][6] [13], \prod_terms[0][6] [13], 
    \prod_terms[0][6] [13],  \prod_terms[0][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I1(.SUM({ n5818_29[18:0] }), .A({n5818_28[17],  n5818_28[17:0] }), .B({
    \prod_terms[0][5] [13], \prod_terms[0][5] [13], \prod_terms[0][5] [13], 
    \prod_terms[0][5] [13], \prod_terms[0][5] [13],  \prod_terms[0][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I1(.SUM({ n5818_28[17:0] }), .A({n5817_30[16],  n5817_30[16:0] }), .B({
    \prod_terms[0][4] [13], \prod_terms[0][4] [13], \prod_terms[0][4] [13], 
    \prod_terms[0][4] [13],  \prod_terms[0][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I1(.SUM({ n5817_30[16:0] }), .A({n5817_29[15],  n5817_29[15:0] }), .B({
    \prod_terms[0][3] [13], \prod_terms[0][3] [13], \prod_terms[0][3] [13],  \prod_terms[0][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I1(.SUM({ n5817_29[15:0] }), .A({n5817_28[14],  n5817_28[14:0] }), .B({
    \prod_terms[0][2] [13], \prod_terms[0][2] [13],  \prod_terms[0][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I1(.SUM({ n5817_28[14:0] }), .A({\prod_terms[0][0] [13],  \prod_terms[0][0] [13:0] }), .B({
    \prod_terms[0][1] [13],  \prod_terms[0][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I2(.SUM({ \row_sums[1] [18:0] }), .A({ n5823_17[18:0] }), .B({\b2_extended[1] [13], 
    \b2_extended[1] [13], \b2_extended[1] [13], \b2_extended[1] [13], 
    \b2_extended[1] [13],  \b2_extended[1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I2(.SUM({ n5823_17[18:0] }), .A({ n5822_27[18:0] }), .B({\prod_terms[1][19] [13], 
    \prod_terms[1][19] [13], \prod_terms[1][19] [13], \prod_terms[1][19] [13], 
    \prod_terms[1][19] [13],  \prod_terms[1][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I2(.SUM({ n5822_27[18:0] }), .A({ n5822_26[18:0] }), .B({\prod_terms[1][18] [13], 
    \prod_terms[1][18] [13], \prod_terms[1][18] [13], \prod_terms[1][18] [13], 
    \prod_terms[1][18] [13],  \prod_terms[1][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I2(.SUM({ n5822_26[18:0] }), .A({ n5822_25[18:0] }), .B({\prod_terms[1][17] [13], 
    \prod_terms[1][17] [13], \prod_terms[1][17] [13], \prod_terms[1][17] [13], 
    \prod_terms[1][17] [13],  \prod_terms[1][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I2(.SUM({ n5822_25[18:0] }), .A({ n5821_27[18:0] }), .B({\prod_terms[1][16] [13], 
    \prod_terms[1][16] [13], \prod_terms[1][16] [13], \prod_terms[1][16] [13], 
    \prod_terms[1][16] [13],  \prod_terms[1][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I2(.SUM({ n5821_27[18:0] }), .A({ n5821_26[18:0] }), .B({\prod_terms[1][15] [13], 
    \prod_terms[1][15] [13], \prod_terms[1][15] [13], \prod_terms[1][15] [13], 
    \prod_terms[1][15] [13],  \prod_terms[1][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I2(.SUM({ n5821_26[18:0] }), .A({ n5821_25[18:0] }), .B({\prod_terms[1][14] [13], 
    \prod_terms[1][14] [13], \prod_terms[1][14] [13], \prod_terms[1][14] [13], 
    \prod_terms[1][14] [13],  \prod_terms[1][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I2(.SUM({ n5821_25[18:0] }), .A({ n5820_27[18:0] }), .B({\prod_terms[1][13] [13], 
    \prod_terms[1][13] [13], \prod_terms[1][13] [13], \prod_terms[1][13] [13], 
    \prod_terms[1][13] [13],  \prod_terms[1][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I2(.SUM({ n5820_27[18:0] }), .A({ n5820_26[18:0] }), .B({\prod_terms[1][12] [13], 
    \prod_terms[1][12] [13], \prod_terms[1][12] [13], \prod_terms[1][12] [13], 
    \prod_terms[1][12] [13],  \prod_terms[1][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I2(.SUM({ n5820_26[18:0] }), .A({ n5820_25[18:0] }), .B({\prod_terms[1][11] [13], 
    \prod_terms[1][11] [13], \prod_terms[1][11] [13], \prod_terms[1][11] [13], 
    \prod_terms[1][11] [13],  \prod_terms[1][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I2(.SUM({ n5820_25[18:0] }), .A({ n5819_27[18:0] }), .B({\prod_terms[1][10] [13], 
    \prod_terms[1][10] [13], \prod_terms[1][10] [13], \prod_terms[1][10] [13], 
    \prod_terms[1][10] [13],  \prod_terms[1][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I2(.SUM({ n5819_27[18:0] }), .A({ n5819_26[18:0] }), .B({\prod_terms[1][9] [13], 
    \prod_terms[1][9] [13], \prod_terms[1][9] [13], \prod_terms[1][9] [13], 
    \prod_terms[1][9] [13],  \prod_terms[1][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I2(.SUM({ n5819_26[18:0] }), .A({ n5819_25[18:0] }), .B({\prod_terms[1][8] [13], 
    \prod_terms[1][8] [13], \prod_terms[1][8] [13], \prod_terms[1][8] [13], 
    \prod_terms[1][8] [13],  \prod_terms[1][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I2(.SUM({ n5819_25[18:0] }), .A({ n5818_27[18:0] }), .B({\prod_terms[1][7] [13], 
    \prod_terms[1][7] [13], \prod_terms[1][7] [13], \prod_terms[1][7] [13], 
    \prod_terms[1][7] [13],  \prod_terms[1][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I2(.SUM({ n5818_27[18:0] }), .A({ n5818_26[18:0] }), .B({\prod_terms[1][6] [13], 
    \prod_terms[1][6] [13], \prod_terms[1][6] [13], \prod_terms[1][6] [13], 
    \prod_terms[1][6] [13],  \prod_terms[1][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I2(.SUM({ n5818_26[18:0] }), .A({n5818_25[17],  n5818_25[17:0] }), .B({
    \prod_terms[1][5] [13], \prod_terms[1][5] [13], \prod_terms[1][5] [13], 
    \prod_terms[1][5] [13], \prod_terms[1][5] [13],  \prod_terms[1][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I2(.SUM({ n5818_25[17:0] }), .A({n5817_27[16],  n5817_27[16:0] }), .B({
    \prod_terms[1][4] [13], \prod_terms[1][4] [13], \prod_terms[1][4] [13], 
    \prod_terms[1][4] [13],  \prod_terms[1][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I2(.SUM({ n5817_27[16:0] }), .A({n5817_26[15],  n5817_26[15:0] }), .B({
    \prod_terms[1][3] [13], \prod_terms[1][3] [13], \prod_terms[1][3] [13],  \prod_terms[1][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I2(.SUM({ n5817_26[15:0] }), .A({n5817_25[14],  n5817_25[14:0] }), .B({
    \prod_terms[1][2] [13], \prod_terms[1][2] [13],  \prod_terms[1][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I2(.SUM({ n5817_25[14:0] }), .A({\prod_terms[1][0] [13],  \prod_terms[1][0] [13:0] }), .B({
    \prod_terms[1][1] [13],  \prod_terms[1][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I3(.SUM({ \row_sums[2] [18:0] }), .A({ n5823_15[18:0] }), .B({\b2_extended[2] [13], 
    \b2_extended[2] [13], \b2_extended[2] [13], \b2_extended[2] [13], 
    \b2_extended[2] [13],  \b2_extended[2] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I3(.SUM({ n5823_15[18:0] }), .A({ n5822_24[18:0] }), .B({\prod_terms[2][19] [13], 
    \prod_terms[2][19] [13], \prod_terms[2][19] [13], \prod_terms[2][19] [13], 
    \prod_terms[2][19] [13],  \prod_terms[2][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I3(.SUM({ n5822_24[18:0] }), .A({ n5822_23[18:0] }), .B({\prod_terms[2][18] [13], 
    \prod_terms[2][18] [13], \prod_terms[2][18] [13], \prod_terms[2][18] [13], 
    \prod_terms[2][18] [13],  \prod_terms[2][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I3(.SUM({ n5822_23[18:0] }), .A({ n5822_22[18:0] }), .B({\prod_terms[2][17] [13], 
    \prod_terms[2][17] [13], \prod_terms[2][17] [13], \prod_terms[2][17] [13], 
    \prod_terms[2][17] [13],  \prod_terms[2][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I3(.SUM({ n5822_22[18:0] }), .A({ n5821_24[18:0] }), .B({\prod_terms[2][16] [13], 
    \prod_terms[2][16] [13], \prod_terms[2][16] [13], \prod_terms[2][16] [13], 
    \prod_terms[2][16] [13],  \prod_terms[2][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I3(.SUM({ n5821_24[18:0] }), .A({ n5821_23[18:0] }), .B({\prod_terms[2][15] [13], 
    \prod_terms[2][15] [13], \prod_terms[2][15] [13], \prod_terms[2][15] [13], 
    \prod_terms[2][15] [13],  \prod_terms[2][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I3(.SUM({ n5821_23[18:0] }), .A({ n5821_22[18:0] }), .B({\prod_terms[2][14] [13], 
    \prod_terms[2][14] [13], \prod_terms[2][14] [13], \prod_terms[2][14] [13], 
    \prod_terms[2][14] [13],  \prod_terms[2][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I3(.SUM({ n5821_22[18:0] }), .A({ n5820_24[18:0] }), .B({\prod_terms[2][13] [13], 
    \prod_terms[2][13] [13], \prod_terms[2][13] [13], \prod_terms[2][13] [13], 
    \prod_terms[2][13] [13],  \prod_terms[2][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I3(.SUM({ n5820_24[18:0] }), .A({ n5820_23[18:0] }), .B({\prod_terms[2][12] [13], 
    \prod_terms[2][12] [13], \prod_terms[2][12] [13], \prod_terms[2][12] [13], 
    \prod_terms[2][12] [13],  \prod_terms[2][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I3(.SUM({ n5820_23[18:0] }), .A({ n5820_22[18:0] }), .B({\prod_terms[2][11] [13], 
    \prod_terms[2][11] [13], \prod_terms[2][11] [13], \prod_terms[2][11] [13], 
    \prod_terms[2][11] [13],  \prod_terms[2][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I3(.SUM({ n5820_22[18:0] }), .A({ n5819_24[18:0] }), .B({\prod_terms[2][10] [13], 
    \prod_terms[2][10] [13], \prod_terms[2][10] [13], \prod_terms[2][10] [13], 
    \prod_terms[2][10] [13],  \prod_terms[2][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I3(.SUM({ n5819_24[18:0] }), .A({ n5819_23[18:0] }), .B({\prod_terms[2][9] [13], 
    \prod_terms[2][9] [13], \prod_terms[2][9] [13], \prod_terms[2][9] [13], 
    \prod_terms[2][9] [13],  \prod_terms[2][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I3(.SUM({ n5819_23[18:0] }), .A({ n5819_22[18:0] }), .B({\prod_terms[2][8] [13], 
    \prod_terms[2][8] [13], \prod_terms[2][8] [13], \prod_terms[2][8] [13], 
    \prod_terms[2][8] [13],  \prod_terms[2][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I3(.SUM({ n5819_22[18:0] }), .A({ n5818_24[18:0] }), .B({\prod_terms[2][7] [13], 
    \prod_terms[2][7] [13], \prod_terms[2][7] [13], \prod_terms[2][7] [13], 
    \prod_terms[2][7] [13],  \prod_terms[2][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I3(.SUM({ n5818_24[18:0] }), .A({ n5818_23[18:0] }), .B({\prod_terms[2][6] [13], 
    \prod_terms[2][6] [13], \prod_terms[2][6] [13], \prod_terms[2][6] [13], 
    \prod_terms[2][6] [13],  \prod_terms[2][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I3(.SUM({ n5818_23[18:0] }), .A({n5818_22[17],  n5818_22[17:0] }), .B({
    \prod_terms[2][5] [13], \prod_terms[2][5] [13], \prod_terms[2][5] [13], 
    \prod_terms[2][5] [13], \prod_terms[2][5] [13],  \prod_terms[2][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I3(.SUM({ n5818_22[17:0] }), .A({n5817_24[16],  n5817_24[16:0] }), .B({
    \prod_terms[2][4] [13], \prod_terms[2][4] [13], \prod_terms[2][4] [13], 
    \prod_terms[2][4] [13],  \prod_terms[2][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I3(.SUM({ n5817_24[16:0] }), .A({n5817_23[15],  n5817_23[15:0] }), .B({
    \prod_terms[2][3] [13], \prod_terms[2][3] [13], \prod_terms[2][3] [13],  \prod_terms[2][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I3(.SUM({ n5817_23[15:0] }), .A({n5817_22[14],  n5817_22[14:0] }), .B({
    \prod_terms[2][2] [13], \prod_terms[2][2] [13],  \prod_terms[2][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I3(.SUM({ n5817_22[14:0] }), .A({\prod_terms[2][0] [13],  \prod_terms[2][0] [13:0] }), .B({
    \prod_terms[2][1] [13],  \prod_terms[2][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I4(.SUM({ \row_sums[3] [18:0] }), .A({ n5823_13[18:0] }), .B({\b2_extended[3] [13], 
    \b2_extended[3] [13], \b2_extended[3] [13], \b2_extended[3] [13], 
    \b2_extended[3] [13],  \b2_extended[3] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I4(.SUM({ n5823_13[18:0] }), .A({ n5822_21[18:0] }), .B({\prod_terms[3][19] [13], 
    \prod_terms[3][19] [13], \prod_terms[3][19] [13], \prod_terms[3][19] [13], 
    \prod_terms[3][19] [13],  \prod_terms[3][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I4(.SUM({ n5822_21[18:0] }), .A({ n5822_20[18:0] }), .B({\prod_terms[3][18] [13], 
    \prod_terms[3][18] [13], \prod_terms[3][18] [13], \prod_terms[3][18] [13], 
    \prod_terms[3][18] [13],  \prod_terms[3][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I4(.SUM({ n5822_20[18:0] }), .A({ n5822_19[18:0] }), .B({\prod_terms[3][17] [13], 
    \prod_terms[3][17] [13], \prod_terms[3][17] [13], \prod_terms[3][17] [13], 
    \prod_terms[3][17] [13],  \prod_terms[3][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I4(.SUM({ n5822_19[18:0] }), .A({ n5821_21[18:0] }), .B({\prod_terms[3][16] [13], 
    \prod_terms[3][16] [13], \prod_terms[3][16] [13], \prod_terms[3][16] [13], 
    \prod_terms[3][16] [13],  \prod_terms[3][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I4(.SUM({ n5821_21[18:0] }), .A({ n5821_20[18:0] }), .B({\prod_terms[3][15] [13], 
    \prod_terms[3][15] [13], \prod_terms[3][15] [13], \prod_terms[3][15] [13], 
    \prod_terms[3][15] [13],  \prod_terms[3][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I4(.SUM({ n5821_20[18:0] }), .A({ n5821_19[18:0] }), .B({\prod_terms[3][14] [13], 
    \prod_terms[3][14] [13], \prod_terms[3][14] [13], \prod_terms[3][14] [13], 
    \prod_terms[3][14] [13],  \prod_terms[3][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I4(.SUM({ n5821_19[18:0] }), .A({ n5820_21[18:0] }), .B({\prod_terms[3][13] [13], 
    \prod_terms[3][13] [13], \prod_terms[3][13] [13], \prod_terms[3][13] [13], 
    \prod_terms[3][13] [13],  \prod_terms[3][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I4(.SUM({ n5820_21[18:0] }), .A({ n5820_20[18:0] }), .B({\prod_terms[3][12] [13], 
    \prod_terms[3][12] [13], \prod_terms[3][12] [13], \prod_terms[3][12] [13], 
    \prod_terms[3][12] [13],  \prod_terms[3][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I4(.SUM({ n5820_20[18:0] }), .A({ n5820_19[18:0] }), .B({\prod_terms[3][11] [13], 
    \prod_terms[3][11] [13], \prod_terms[3][11] [13], \prod_terms[3][11] [13], 
    \prod_terms[3][11] [13],  \prod_terms[3][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I4(.SUM({ n5820_19[18:0] }), .A({ n5819_21[18:0] }), .B({\prod_terms[3][10] [13], 
    \prod_terms[3][10] [13], \prod_terms[3][10] [13], \prod_terms[3][10] [13], 
    \prod_terms[3][10] [13],  \prod_terms[3][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I4(.SUM({ n5819_21[18:0] }), .A({ n5819_20[18:0] }), .B({\prod_terms[3][9] [13], 
    \prod_terms[3][9] [13], \prod_terms[3][9] [13], \prod_terms[3][9] [13], 
    \prod_terms[3][9] [13],  \prod_terms[3][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I4(.SUM({ n5819_20[18:0] }), .A({ n5819_19[18:0] }), .B({\prod_terms[3][8] [13], 
    \prod_terms[3][8] [13], \prod_terms[3][8] [13], \prod_terms[3][8] [13], 
    \prod_terms[3][8] [13],  \prod_terms[3][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I4(.SUM({ n5819_19[18:0] }), .A({ n5818_21[18:0] }), .B({\prod_terms[3][7] [13], 
    \prod_terms[3][7] [13], \prod_terms[3][7] [13], \prod_terms[3][7] [13], 
    \prod_terms[3][7] [13],  \prod_terms[3][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I4(.SUM({ n5818_21[18:0] }), .A({ n5818_20[18:0] }), .B({\prod_terms[3][6] [13], 
    \prod_terms[3][6] [13], \prod_terms[3][6] [13], \prod_terms[3][6] [13], 
    \prod_terms[3][6] [13],  \prod_terms[3][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I4(.SUM({ n5818_20[18:0] }), .A({n5818_19[17],  n5818_19[17:0] }), .B({
    \prod_terms[3][5] [13], \prod_terms[3][5] [13], \prod_terms[3][5] [13], 
    \prod_terms[3][5] [13], \prod_terms[3][5] [13],  \prod_terms[3][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I4(.SUM({ n5818_19[17:0] }), .A({n5817_21[16],  n5817_21[16:0] }), .B({
    \prod_terms[3][4] [13], \prod_terms[3][4] [13], \prod_terms[3][4] [13], 
    \prod_terms[3][4] [13],  \prod_terms[3][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I4(.SUM({ n5817_21[16:0] }), .A({n5817_20[15],  n5817_20[15:0] }), .B({
    \prod_terms[3][3] [13], \prod_terms[3][3] [13], \prod_terms[3][3] [13],  \prod_terms[3][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I4(.SUM({ n5817_20[15:0] }), .A({n5817_19[14],  n5817_19[14:0] }), .B({
    \prod_terms[3][2] [13], \prod_terms[3][2] [13],  \prod_terms[3][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I4(.SUM({ n5817_19[14:0] }), .A({\prod_terms[3][0] [13],  \prod_terms[3][0] [13:0] }), .B({
    \prod_terms[3][1] [13],  \prod_terms[3][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I5(.SUM({ \row_sums[4] [18:0] }), .A({ n5823_11[18:0] }), .B({\b2_extended[4] [13], 
    \b2_extended[4] [13], \b2_extended[4] [13], \b2_extended[4] [13], 
    \b2_extended[4] [13],  \b2_extended[4] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I5(.SUM({ n5823_11[18:0] }), .A({ n5822_18[18:0] }), .B({\prod_terms[4][19] [13], 
    \prod_terms[4][19] [13], \prod_terms[4][19] [13], \prod_terms[4][19] [13], 
    \prod_terms[4][19] [13],  \prod_terms[4][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I5(.SUM({ n5822_18[18:0] }), .A({ n5822_17[18:0] }), .B({\prod_terms[4][18] [13], 
    \prod_terms[4][18] [13], \prod_terms[4][18] [13], \prod_terms[4][18] [13], 
    \prod_terms[4][18] [13],  \prod_terms[4][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I5(.SUM({ n5822_17[18:0] }), .A({ n5822_16[18:0] }), .B({\prod_terms[4][17] [13], 
    \prod_terms[4][17] [13], \prod_terms[4][17] [13], \prod_terms[4][17] [13], 
    \prod_terms[4][17] [13],  \prod_terms[4][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I5(.SUM({ n5822_16[18:0] }), .A({ n5821_18[18:0] }), .B({\prod_terms[4][16] [13], 
    \prod_terms[4][16] [13], \prod_terms[4][16] [13], \prod_terms[4][16] [13], 
    \prod_terms[4][16] [13],  \prod_terms[4][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I5(.SUM({ n5821_18[18:0] }), .A({ n5821_17[18:0] }), .B({\prod_terms[4][15] [13], 
    \prod_terms[4][15] [13], \prod_terms[4][15] [13], \prod_terms[4][15] [13], 
    \prod_terms[4][15] [13],  \prod_terms[4][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I5(.SUM({ n5821_17[18:0] }), .A({ n5821_16[18:0] }), .B({\prod_terms[4][14] [13], 
    \prod_terms[4][14] [13], \prod_terms[4][14] [13], \prod_terms[4][14] [13], 
    \prod_terms[4][14] [13],  \prod_terms[4][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I5(.SUM({ n5821_16[18:0] }), .A({ n5820_18[18:0] }), .B({\prod_terms[4][13] [13], 
    \prod_terms[4][13] [13], \prod_terms[4][13] [13], \prod_terms[4][13] [13], 
    \prod_terms[4][13] [13],  \prod_terms[4][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I5(.SUM({ n5820_18[18:0] }), .A({ n5820_17[18:0] }), .B({\prod_terms[4][12] [13], 
    \prod_terms[4][12] [13], \prod_terms[4][12] [13], \prod_terms[4][12] [13], 
    \prod_terms[4][12] [13],  \prod_terms[4][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I5(.SUM({ n5820_17[18:0] }), .A({ n5820_16[18:0] }), .B({\prod_terms[4][11] [13], 
    \prod_terms[4][11] [13], \prod_terms[4][11] [13], \prod_terms[4][11] [13], 
    \prod_terms[4][11] [13],  \prod_terms[4][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I5(.SUM({ n5820_16[18:0] }), .A({ n5819_18[18:0] }), .B({\prod_terms[4][10] [13], 
    \prod_terms[4][10] [13], \prod_terms[4][10] [13], \prod_terms[4][10] [13], 
    \prod_terms[4][10] [13],  \prod_terms[4][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I5(.SUM({ n5819_18[18:0] }), .A({ n5819_17[18:0] }), .B({\prod_terms[4][9] [13], 
    \prod_terms[4][9] [13], \prod_terms[4][9] [13], \prod_terms[4][9] [13], 
    \prod_terms[4][9] [13],  \prod_terms[4][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I5(.SUM({ n5819_17[18:0] }), .A({ n5819_16[18:0] }), .B({\prod_terms[4][8] [13], 
    \prod_terms[4][8] [13], \prod_terms[4][8] [13], \prod_terms[4][8] [13], 
    \prod_terms[4][8] [13],  \prod_terms[4][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I5(.SUM({ n5819_16[18:0] }), .A({ n5818_18[18:0] }), .B({\prod_terms[4][7] [13], 
    \prod_terms[4][7] [13], \prod_terms[4][7] [13], \prod_terms[4][7] [13], 
    \prod_terms[4][7] [13],  \prod_terms[4][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I5(.SUM({ n5818_18[18:0] }), .A({ n5818_17[18:0] }), .B({\prod_terms[4][6] [13], 
    \prod_terms[4][6] [13], \prod_terms[4][6] [13], \prod_terms[4][6] [13], 
    \prod_terms[4][6] [13],  \prod_terms[4][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I5(.SUM({ n5818_17[18:0] }), .A({n5818_16[17],  n5818_16[17:0] }), .B({
    \prod_terms[4][5] [13], \prod_terms[4][5] [13], \prod_terms[4][5] [13], 
    \prod_terms[4][5] [13], \prod_terms[4][5] [13],  \prod_terms[4][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I5(.SUM({ n5818_16[17:0] }), .A({n5817_18[16],  n5817_18[16:0] }), .B({
    \prod_terms[4][4] [13], \prod_terms[4][4] [13], \prod_terms[4][4] [13], 
    \prod_terms[4][4] [13],  \prod_terms[4][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I5(.SUM({ n5817_18[16:0] }), .A({n5817_17[15],  n5817_17[15:0] }), .B({
    \prod_terms[4][3] [13], \prod_terms[4][3] [13], \prod_terms[4][3] [13],  \prod_terms[4][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I5(.SUM({ n5817_17[15:0] }), .A({n5817_16[14],  n5817_16[14:0] }), .B({
    \prod_terms[4][2] [13], \prod_terms[4][2] [13],  \prod_terms[4][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I5(.SUM({ n5817_16[14:0] }), .A({\prod_terms[4][0] [13],  \prod_terms[4][0] [13:0] }), .B({
    \prod_terms[4][1] [13],  \prod_terms[4][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I6(.SUM({ \row_sums[5] [18:0] }), .A({ n5823_9[18:0] }), .B({\b2_extended[5] [13], 
    \b2_extended[5] [13], \b2_extended[5] [13], \b2_extended[5] [13], 
    \b2_extended[5] [13],  \b2_extended[5] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I6(.SUM({ n5823_9[18:0] }), .A({ n5822_15[18:0] }), .B({\prod_terms[5][19] [13], 
    \prod_terms[5][19] [13], \prod_terms[5][19] [13], \prod_terms[5][19] [13], 
    \prod_terms[5][19] [13],  \prod_terms[5][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I6(.SUM({ n5822_15[18:0] }), .A({ n5822_14[18:0] }), .B({\prod_terms[5][18] [13], 
    \prod_terms[5][18] [13], \prod_terms[5][18] [13], \prod_terms[5][18] [13], 
    \prod_terms[5][18] [13],  \prod_terms[5][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I6(.SUM({ n5822_14[18:0] }), .A({ n5822_13[18:0] }), .B({\prod_terms[5][17] [13], 
    \prod_terms[5][17] [13], \prod_terms[5][17] [13], \prod_terms[5][17] [13], 
    \prod_terms[5][17] [13],  \prod_terms[5][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I6(.SUM({ n5822_13[18:0] }), .A({ n5821_15[18:0] }), .B({\prod_terms[5][16] [13], 
    \prod_terms[5][16] [13], \prod_terms[5][16] [13], \prod_terms[5][16] [13], 
    \prod_terms[5][16] [13],  \prod_terms[5][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I6(.SUM({ n5821_15[18:0] }), .A({ n5821_14[18:0] }), .B({\prod_terms[5][15] [13], 
    \prod_terms[5][15] [13], \prod_terms[5][15] [13], \prod_terms[5][15] [13], 
    \prod_terms[5][15] [13],  \prod_terms[5][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I6(.SUM({ n5821_14[18:0] }), .A({ n5821_13[18:0] }), .B({\prod_terms[5][14] [13], 
    \prod_terms[5][14] [13], \prod_terms[5][14] [13], \prod_terms[5][14] [13], 
    \prod_terms[5][14] [13],  \prod_terms[5][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I6(.SUM({ n5821_13[18:0] }), .A({ n5820_15[18:0] }), .B({\prod_terms[5][13] [13], 
    \prod_terms[5][13] [13], \prod_terms[5][13] [13], \prod_terms[5][13] [13], 
    \prod_terms[5][13] [13],  \prod_terms[5][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I6(.SUM({ n5820_15[18:0] }), .A({ n5820_14[18:0] }), .B({\prod_terms[5][12] [13], 
    \prod_terms[5][12] [13], \prod_terms[5][12] [13], \prod_terms[5][12] [13], 
    \prod_terms[5][12] [13],  \prod_terms[5][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I6(.SUM({ n5820_14[18:0] }), .A({ n5820_13[18:0] }), .B({\prod_terms[5][11] [13], 
    \prod_terms[5][11] [13], \prod_terms[5][11] [13], \prod_terms[5][11] [13], 
    \prod_terms[5][11] [13],  \prod_terms[5][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I6(.SUM({ n5820_13[18:0] }), .A({ n5819_15[18:0] }), .B({\prod_terms[5][10] [13], 
    \prod_terms[5][10] [13], \prod_terms[5][10] [13], \prod_terms[5][10] [13], 
    \prod_terms[5][10] [13],  \prod_terms[5][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I6(.SUM({ n5819_15[18:0] }), .A({ n5819_14[18:0] }), .B({\prod_terms[5][9] [13], 
    \prod_terms[5][9] [13], \prod_terms[5][9] [13], \prod_terms[5][9] [13], 
    \prod_terms[5][9] [13],  \prod_terms[5][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I6(.SUM({ n5819_14[18:0] }), .A({ n5819_13[18:0] }), .B({\prod_terms[5][8] [13], 
    \prod_terms[5][8] [13], \prod_terms[5][8] [13], \prod_terms[5][8] [13], 
    \prod_terms[5][8] [13],  \prod_terms[5][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I6(.SUM({ n5819_13[18:0] }), .A({ n5818_15[18:0] }), .B({\prod_terms[5][7] [13], 
    \prod_terms[5][7] [13], \prod_terms[5][7] [13], \prod_terms[5][7] [13], 
    \prod_terms[5][7] [13],  \prod_terms[5][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I6(.SUM({ n5818_15[18:0] }), .A({ n5818_14[18:0] }), .B({\prod_terms[5][6] [13], 
    \prod_terms[5][6] [13], \prod_terms[5][6] [13], \prod_terms[5][6] [13], 
    \prod_terms[5][6] [13],  \prod_terms[5][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I6(.SUM({ n5818_14[18:0] }), .A({n5818_13[17],  n5818_13[17:0] }), .B({
    \prod_terms[5][5] [13], \prod_terms[5][5] [13], \prod_terms[5][5] [13], 
    \prod_terms[5][5] [13], \prod_terms[5][5] [13],  \prod_terms[5][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I6(.SUM({ n5818_13[17:0] }), .A({n5817_15[16],  n5817_15[16:0] }), .B({
    \prod_terms[5][4] [13], \prod_terms[5][4] [13], \prod_terms[5][4] [13], 
    \prod_terms[5][4] [13],  \prod_terms[5][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I6(.SUM({ n5817_15[16:0] }), .A({n5817_14[15],  n5817_14[15:0] }), .B({
    \prod_terms[5][3] [13], \prod_terms[5][3] [13], \prod_terms[5][3] [13],  \prod_terms[5][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I6(.SUM({ n5817_14[15:0] }), .A({n5817_13[14],  n5817_13[14:0] }), .B({
    \prod_terms[5][2] [13], \prod_terms[5][2] [13],  \prod_terms[5][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I6(.SUM({ n5817_13[14:0] }), .A({\prod_terms[5][0] [13],  \prod_terms[5][0] [13:0] }), .B({
    \prod_terms[5][1] [13],  \prod_terms[5][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I7(.SUM({ \row_sums[6] [18:0] }), .A({ n5823_7[18:0] }), .B({\b2_extended[6] [13], 
    \b2_extended[6] [13], \b2_extended[6] [13], \b2_extended[6] [13], 
    \b2_extended[6] [13],  \b2_extended[6] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I7(.SUM({ n5823_7[18:0] }), .A({ n5822_12[18:0] }), .B({\prod_terms[6][19] [13], 
    \prod_terms[6][19] [13], \prod_terms[6][19] [13], \prod_terms[6][19] [13], 
    \prod_terms[6][19] [13],  \prod_terms[6][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I7(.SUM({ n5822_12[18:0] }), .A({ n5822_11[18:0] }), .B({\prod_terms[6][18] [13], 
    \prod_terms[6][18] [13], \prod_terms[6][18] [13], \prod_terms[6][18] [13], 
    \prod_terms[6][18] [13],  \prod_terms[6][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I7(.SUM({ n5822_11[18:0] }), .A({ n5822_10[18:0] }), .B({\prod_terms[6][17] [13], 
    \prod_terms[6][17] [13], \prod_terms[6][17] [13], \prod_terms[6][17] [13], 
    \prod_terms[6][17] [13],  \prod_terms[6][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I7(.SUM({ n5822_10[18:0] }), .A({ n5821_12[18:0] }), .B({\prod_terms[6][16] [13], 
    \prod_terms[6][16] [13], \prod_terms[6][16] [13], \prod_terms[6][16] [13], 
    \prod_terms[6][16] [13],  \prod_terms[6][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I7(.SUM({ n5821_12[18:0] }), .A({ n5821_11[18:0] }), .B({\prod_terms[6][15] [13], 
    \prod_terms[6][15] [13], \prod_terms[6][15] [13], \prod_terms[6][15] [13], 
    \prod_terms[6][15] [13],  \prod_terms[6][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I7(.SUM({ n5821_11[18:0] }), .A({ n5821_10[18:0] }), .B({\prod_terms[6][14] [13], 
    \prod_terms[6][14] [13], \prod_terms[6][14] [13], \prod_terms[6][14] [13], 
    \prod_terms[6][14] [13],  \prod_terms[6][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I7(.SUM({ n5821_10[18:0] }), .A({ n5820_12[18:0] }), .B({\prod_terms[6][13] [13], 
    \prod_terms[6][13] [13], \prod_terms[6][13] [13], \prod_terms[6][13] [13], 
    \prod_terms[6][13] [13],  \prod_terms[6][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I7(.SUM({ n5820_12[18:0] }), .A({ n5820_11[18:0] }), .B({\prod_terms[6][12] [13], 
    \prod_terms[6][12] [13], \prod_terms[6][12] [13], \prod_terms[6][12] [13], 
    \prod_terms[6][12] [13],  \prod_terms[6][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I7(.SUM({ n5820_11[18:0] }), .A({ n5820_10[18:0] }), .B({\prod_terms[6][11] [13], 
    \prod_terms[6][11] [13], \prod_terms[6][11] [13], \prod_terms[6][11] [13], 
    \prod_terms[6][11] [13],  \prod_terms[6][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I7(.SUM({ n5820_10[18:0] }), .A({ n5819_12[18:0] }), .B({\prod_terms[6][10] [13], 
    \prod_terms[6][10] [13], \prod_terms[6][10] [13], \prod_terms[6][10] [13], 
    \prod_terms[6][10] [13],  \prod_terms[6][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I7(.SUM({ n5819_12[18:0] }), .A({ n5819_11[18:0] }), .B({\prod_terms[6][9] [13], 
    \prod_terms[6][9] [13], \prod_terms[6][9] [13], \prod_terms[6][9] [13], 
    \prod_terms[6][9] [13],  \prod_terms[6][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I7(.SUM({ n5819_11[18:0] }), .A({ n5819_10[18:0] }), .B({\prod_terms[6][8] [13], 
    \prod_terms[6][8] [13], \prod_terms[6][8] [13], \prod_terms[6][8] [13], 
    \prod_terms[6][8] [13],  \prod_terms[6][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I7(.SUM({ n5819_10[18:0] }), .A({ n5818_12[18:0] }), .B({\prod_terms[6][7] [13], 
    \prod_terms[6][7] [13], \prod_terms[6][7] [13], \prod_terms[6][7] [13], 
    \prod_terms[6][7] [13],  \prod_terms[6][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I7(.SUM({ n5818_12[18:0] }), .A({ n5818_11[18:0] }), .B({\prod_terms[6][6] [13], 
    \prod_terms[6][6] [13], \prod_terms[6][6] [13], \prod_terms[6][6] [13], 
    \prod_terms[6][6] [13],  \prod_terms[6][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I7(.SUM({ n5818_11[18:0] }), .A({n5818_10[17],  n5818_10[17:0] }), .B({
    \prod_terms[6][5] [13], \prod_terms[6][5] [13], \prod_terms[6][5] [13], 
    \prod_terms[6][5] [13], \prod_terms[6][5] [13],  \prod_terms[6][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I7(.SUM({ n5818_10[17:0] }), .A({n5817_12[16],  n5817_12[16:0] }), .B({
    \prod_terms[6][4] [13], \prod_terms[6][4] [13], \prod_terms[6][4] [13], 
    \prod_terms[6][4] [13],  \prod_terms[6][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I7(.SUM({ n5817_12[16:0] }), .A({n5817_11[15],  n5817_11[15:0] }), .B({
    \prod_terms[6][3] [13], \prod_terms[6][3] [13], \prod_terms[6][3] [13],  \prod_terms[6][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I7(.SUM({ n5817_11[15:0] }), .A({n5817_10[14],  n5817_10[14:0] }), .B({
    \prod_terms[6][2] [13], \prod_terms[6][2] [13],  \prod_terms[6][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I7(.SUM({ n5817_10[14:0] }), .A({\prod_terms[6][0] [13],  \prod_terms[6][0] [13:0] }), .B({
    \prod_terms[6][1] [13],  \prod_terms[6][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I8(.SUM({ \row_sums[7] [18:0] }), .A({ n5823_5[18:0] }), .B({\b2_extended[7] [13], 
    \b2_extended[7] [13], \b2_extended[7] [13], \b2_extended[7] [13], 
    \b2_extended[7] [13],  \b2_extended[7] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I8(.SUM({ n5823_5[18:0] }), .A({ n5822_9[18:0] }), .B({\prod_terms[7][19] [13], 
    \prod_terms[7][19] [13], \prod_terms[7][19] [13], \prod_terms[7][19] [13], 
    \prod_terms[7][19] [13],  \prod_terms[7][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I8(.SUM({ n5822_9[18:0] }), .A({ n5822_8[18:0] }), .B({\prod_terms[7][18] [13], 
    \prod_terms[7][18] [13], \prod_terms[7][18] [13], \prod_terms[7][18] [13], 
    \prod_terms[7][18] [13],  \prod_terms[7][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I8(.SUM({ n5822_8[18:0] }), .A({ n5822_7[18:0] }), .B({\prod_terms[7][17] [13], 
    \prod_terms[7][17] [13], \prod_terms[7][17] [13], \prod_terms[7][17] [13], 
    \prod_terms[7][17] [13],  \prod_terms[7][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I8(.SUM({ n5822_7[18:0] }), .A({ n5821_9[18:0] }), .B({\prod_terms[7][16] [13], 
    \prod_terms[7][16] [13], \prod_terms[7][16] [13], \prod_terms[7][16] [13], 
    \prod_terms[7][16] [13],  \prod_terms[7][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I8(.SUM({ n5821_9[18:0] }), .A({ n5821_8[18:0] }), .B({\prod_terms[7][15] [13], 
    \prod_terms[7][15] [13], \prod_terms[7][15] [13], \prod_terms[7][15] [13], 
    \prod_terms[7][15] [13],  \prod_terms[7][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I8(.SUM({ n5821_8[18:0] }), .A({ n5821_7[18:0] }), .B({\prod_terms[7][14] [13], 
    \prod_terms[7][14] [13], \prod_terms[7][14] [13], \prod_terms[7][14] [13], 
    \prod_terms[7][14] [13],  \prod_terms[7][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I8(.SUM({ n5821_7[18:0] }), .A({ n5820_9[18:0] }), .B({\prod_terms[7][13] [13], 
    \prod_terms[7][13] [13], \prod_terms[7][13] [13], \prod_terms[7][13] [13], 
    \prod_terms[7][13] [13],  \prod_terms[7][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I8(.SUM({ n5820_9[18:0] }), .A({ n5820_8[18:0] }), .B({\prod_terms[7][12] [13], 
    \prod_terms[7][12] [13], \prod_terms[7][12] [13], \prod_terms[7][12] [13], 
    \prod_terms[7][12] [13],  \prod_terms[7][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I8(.SUM({ n5820_8[18:0] }), .A({ n5820_7[18:0] }), .B({\prod_terms[7][11] [13], 
    \prod_terms[7][11] [13], \prod_terms[7][11] [13], \prod_terms[7][11] [13], 
    \prod_terms[7][11] [13],  \prod_terms[7][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I8(.SUM({ n5820_7[18:0] }), .A({ n5819_9[18:0] }), .B({\prod_terms[7][10] [13], 
    \prod_terms[7][10] [13], \prod_terms[7][10] [13], \prod_terms[7][10] [13], 
    \prod_terms[7][10] [13],  \prod_terms[7][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I8(.SUM({ n5819_9[18:0] }), .A({ n5819_8[18:0] }), .B({\prod_terms[7][9] [13], 
    \prod_terms[7][9] [13], \prod_terms[7][9] [13], \prod_terms[7][9] [13], 
    \prod_terms[7][9] [13],  \prod_terms[7][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I8(.SUM({ n5819_8[18:0] }), .A({ n5819_7[18:0] }), .B({\prod_terms[7][8] [13], 
    \prod_terms[7][8] [13], \prod_terms[7][8] [13], \prod_terms[7][8] [13], 
    \prod_terms[7][8] [13],  \prod_terms[7][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I8(.SUM({ n5819_7[18:0] }), .A({ n5818_9[18:0] }), .B({\prod_terms[7][7] [13], 
    \prod_terms[7][7] [13], \prod_terms[7][7] [13], \prod_terms[7][7] [13], 
    \prod_terms[7][7] [13],  \prod_terms[7][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I8(.SUM({ n5818_9[18:0] }), .A({ n5818_8[18:0] }), .B({\prod_terms[7][6] [13], 
    \prod_terms[7][6] [13], \prod_terms[7][6] [13], \prod_terms[7][6] [13], 
    \prod_terms[7][6] [13],  \prod_terms[7][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I8(.SUM({ n5818_8[18:0] }), .A({n5818_7[17],  n5818_7[17:0] }), .B({
    \prod_terms[7][5] [13], \prod_terms[7][5] [13], \prod_terms[7][5] [13], 
    \prod_terms[7][5] [13], \prod_terms[7][5] [13],  \prod_terms[7][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I8(.SUM({ n5818_7[17:0] }), .A({n5817_9[16],  n5817_9[16:0] }), .B({
    \prod_terms[7][4] [13], \prod_terms[7][4] [13], \prod_terms[7][4] [13], 
    \prod_terms[7][4] [13],  \prod_terms[7][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I8(.SUM({ n5817_9[16:0] }), .A({n5817_8[15],  n5817_8[15:0] }), .B({
    \prod_terms[7][3] [13], \prod_terms[7][3] [13], \prod_terms[7][3] [13],  \prod_terms[7][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I8(.SUM({ n5817_8[15:0] }), .A({n5817_7[14],  n5817_7[14:0] }), .B({
    \prod_terms[7][2] [13], \prod_terms[7][2] [13],  \prod_terms[7][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I8(.SUM({ n5817_7[14:0] }), .A({\prod_terms[7][0] [13],  \prod_terms[7][0] [13:0] }), .B({
    \prod_terms[7][1] [13],  \prod_terms[7][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I9(.SUM({ \row_sums[8] [18:0] }), .A({ n5823_3[18:0] }), .B({\b2_extended[8] [13], 
    \b2_extended[8] [13], \b2_extended[8] [13], \b2_extended[8] [13], 
    \b2_extended[8] [13],  \b2_extended[8] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I9(.SUM({ n5823_3[18:0] }), .A({ n5822_6[18:0] }), .B({\prod_terms[8][19] [13], 
    \prod_terms[8][19] [13], \prod_terms[8][19] [13], \prod_terms[8][19] [13], 
    \prod_terms[8][19] [13],  \prod_terms[8][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I9(.SUM({ n5822_6[18:0] }), .A({ n5822_5[18:0] }), .B({\prod_terms[8][18] [13], 
    \prod_terms[8][18] [13], \prod_terms[8][18] [13], \prod_terms[8][18] [13], 
    \prod_terms[8][18] [13],  \prod_terms[8][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I9(.SUM({ n5822_5[18:0] }), .A({ n5822_4[18:0] }), .B({\prod_terms[8][17] [13], 
    \prod_terms[8][17] [13], \prod_terms[8][17] [13], \prod_terms[8][17] [13], 
    \prod_terms[8][17] [13],  \prod_terms[8][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I9(.SUM({ n5822_4[18:0] }), .A({ n5821_6[18:0] }), .B({\prod_terms[8][16] [13], 
    \prod_terms[8][16] [13], \prod_terms[8][16] [13], \prod_terms[8][16] [13], 
    \prod_terms[8][16] [13],  \prod_terms[8][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I9(.SUM({ n5821_6[18:0] }), .A({ n5821_5[18:0] }), .B({\prod_terms[8][15] [13], 
    \prod_terms[8][15] [13], \prod_terms[8][15] [13], \prod_terms[8][15] [13], 
    \prod_terms[8][15] [13],  \prod_terms[8][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I9(.SUM({ n5821_5[18:0] }), .A({ n5821_4[18:0] }), .B({\prod_terms[8][14] [13], 
    \prod_terms[8][14] [13], \prod_terms[8][14] [13], \prod_terms[8][14] [13], 
    \prod_terms[8][14] [13],  \prod_terms[8][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I9(.SUM({ n5821_4[18:0] }), .A({ n5820_6[18:0] }), .B({\prod_terms[8][13] [13], 
    \prod_terms[8][13] [13], \prod_terms[8][13] [13], \prod_terms[8][13] [13], 
    \prod_terms[8][13] [13],  \prod_terms[8][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I9(.SUM({ n5820_6[18:0] }), .A({ n5820_5[18:0] }), .B({\prod_terms[8][12] [13], 
    \prod_terms[8][12] [13], \prod_terms[8][12] [13], \prod_terms[8][12] [13], 
    \prod_terms[8][12] [13],  \prod_terms[8][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I9(.SUM({ n5820_5[18:0] }), .A({ n5820_4[18:0] }), .B({\prod_terms[8][11] [13], 
    \prod_terms[8][11] [13], \prod_terms[8][11] [13], \prod_terms[8][11] [13], 
    \prod_terms[8][11] [13],  \prod_terms[8][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I9(.SUM({ n5820_4[18:0] }), .A({ n5819_6[18:0] }), .B({\prod_terms[8][10] [13], 
    \prod_terms[8][10] [13], \prod_terms[8][10] [13], \prod_terms[8][10] [13], 
    \prod_terms[8][10] [13],  \prod_terms[8][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I9(.SUM({ n5819_6[18:0] }), .A({ n5819_5[18:0] }), .B({\prod_terms[8][9] [13], 
    \prod_terms[8][9] [13], \prod_terms[8][9] [13], \prod_terms[8][9] [13], 
    \prod_terms[8][9] [13],  \prod_terms[8][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I9(.SUM({ n5819_5[18:0] }), .A({ n5819_4[18:0] }), .B({\prod_terms[8][8] [13], 
    \prod_terms[8][8] [13], \prod_terms[8][8] [13], \prod_terms[8][8] [13], 
    \prod_terms[8][8] [13],  \prod_terms[8][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I9(.SUM({ n5819_4[18:0] }), .A({ n5818_6[18:0] }), .B({\prod_terms[8][7] [13], 
    \prod_terms[8][7] [13], \prod_terms[8][7] [13], \prod_terms[8][7] [13], 
    \prod_terms[8][7] [13],  \prod_terms[8][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I9(.SUM({ n5818_6[18:0] }), .A({ n5818_5[18:0] }), .B({\prod_terms[8][6] [13], 
    \prod_terms[8][6] [13], \prod_terms[8][6] [13], \prod_terms[8][6] [13], 
    \prod_terms[8][6] [13],  \prod_terms[8][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I9(.SUM({ n5818_5[18:0] }), .A({n5818_4[17],  n5818_4[17:0] }), .B({
    \prod_terms[8][5] [13], \prod_terms[8][5] [13], \prod_terms[8][5] [13], 
    \prod_terms[8][5] [13], \prod_terms[8][5] [13],  \prod_terms[8][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I9(.SUM({ n5818_4[17:0] }), .A({n5817_6[16],  n5817_6[16:0] }), .B({
    \prod_terms[8][4] [13], \prod_terms[8][4] [13], \prod_terms[8][4] [13], 
    \prod_terms[8][4] [13],  \prod_terms[8][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I9(.SUM({ n5817_6[16:0] }), .A({n5817_5[15],  n5817_5[15:0] }), .B({
    \prod_terms[8][3] [13], \prod_terms[8][3] [13], \prod_terms[8][3] [13],  \prod_terms[8][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I9(.SUM({ n5817_5[15:0] }), .A({n5817_4[14],  n5817_4[14:0] }), .B({
    \prod_terms[8][2] [13], \prod_terms[8][2] [13],  \prod_terms[8][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I9(.SUM({ n5817_4[14:0] }), .A({\prod_terms[8][0] [13],  \prod_terms[8][0] [13:0] }), .B({
    \prod_terms[8][1] [13],  \prod_terms[8][1] [13:0] }));
  VDW_ADD_19_1_0 add_5823_68_I10(.SUM({ \row_sums[9] [18:0] }), .A({ n5823[18:0] }), .B({\b2_extended[9] [13], 
    \b2_extended[9] [13], \b2_extended[9] [13], \b2_extended[9] [13], 
    \b2_extended[9] [13],  \b2_extended[9] [13:0] }));
  VDW_ADD_19_1_0 add_5823_48_I10(.SUM({ n5823[18:0] }), .A({ n5822_3[18:0] }), .B({\prod_terms[9][19] [13], 
    \prod_terms[9][19] [13], \prod_terms[9][19] [13], \prod_terms[9][19] [13], 
    \prod_terms[9][19] [13],  \prod_terms[9][19] [13:0] }));
  VDW_ADD_19_1_0 add_5822_88_I10(.SUM({ n5822_3[18:0] }), .A({ n5822_2[18:0] }), .B({\prod_terms[9][18] [13], 
    \prod_terms[9][18] [13], \prod_terms[9][18] [13], \prod_terms[9][18] [13], 
    \prod_terms[9][18] [13],  \prod_terms[9][18] [13:0] }));
  VDW_ADD_19_1_0 add_5822_68_I10(.SUM({ n5822_2[18:0] }), .A({ n5822[18:0] }), .B({\prod_terms[9][17] [13], 
    \prod_terms[9][17] [13], \prod_terms[9][17] [13], \prod_terms[9][17] [13], 
    \prod_terms[9][17] [13],  \prod_terms[9][17] [13:0] }));
  VDW_ADD_19_1_0 add_5822_48_I10(.SUM({ n5822[18:0] }), .A({ n5821_3[18:0] }), .B({\prod_terms[9][16] [13], 
    \prod_terms[9][16] [13], \prod_terms[9][16] [13], \prod_terms[9][16] [13], 
    \prod_terms[9][16] [13],  \prod_terms[9][16] [13:0] }));
  VDW_ADD_19_1_0 add_5821_88_I10(.SUM({ n5821_3[18:0] }), .A({ n5821_2[18:0] }), .B({\prod_terms[9][15] [13], 
    \prod_terms[9][15] [13], \prod_terms[9][15] [13], \prod_terms[9][15] [13], 
    \prod_terms[9][15] [13],  \prod_terms[9][15] [13:0] }));
  VDW_ADD_19_1_0 add_5821_68_I10(.SUM({ n5821_2[18:0] }), .A({ n5821[18:0] }), .B({\prod_terms[9][14] [13], 
    \prod_terms[9][14] [13], \prod_terms[9][14] [13], \prod_terms[9][14] [13], 
    \prod_terms[9][14] [13],  \prod_terms[9][14] [13:0] }));
  VDW_ADD_19_1_0 add_5821_48_I10(.SUM({ n5821[18:0] }), .A({ n5820_3[18:0] }), .B({\prod_terms[9][13] [13], 
    \prod_terms[9][13] [13], \prod_terms[9][13] [13], \prod_terms[9][13] [13], 
    \prod_terms[9][13] [13],  \prod_terms[9][13] [13:0] }));
  VDW_ADD_19_1_0 add_5820_88_I10(.SUM({ n5820_3[18:0] }), .A({ n5820_2[18:0] }), .B({\prod_terms[9][12] [13], 
    \prod_terms[9][12] [13], \prod_terms[9][12] [13], \prod_terms[9][12] [13], 
    \prod_terms[9][12] [13],  \prod_terms[9][12] [13:0] }));
  VDW_ADD_19_1_0 add_5820_68_I10(.SUM({ n5820_2[18:0] }), .A({ n5820[18:0] }), .B({\prod_terms[9][11] [13], 
    \prod_terms[9][11] [13], \prod_terms[9][11] [13], \prod_terms[9][11] [13], 
    \prod_terms[9][11] [13],  \prod_terms[9][11] [13:0] }));
  VDW_ADD_19_1_0 add_5820_48_I10(.SUM({ n5820[18:0] }), .A({ n5819_3[18:0] }), .B({\prod_terms[9][10] [13], 
    \prod_terms[9][10] [13], \prod_terms[9][10] [13], \prod_terms[9][10] [13], 
    \prod_terms[9][10] [13],  \prod_terms[9][10] [13:0] }));
  VDW_ADD_19_1_0 add_5819_88_I10(.SUM({ n5819_3[18:0] }), .A({ n5819_2[18:0] }), .B({\prod_terms[9][9] [13], 
    \prod_terms[9][9] [13], \prod_terms[9][9] [13], \prod_terms[9][9] [13], 
    \prod_terms[9][9] [13],  \prod_terms[9][9] [13:0] }));
  VDW_ADD_19_1_0 add_5819_68_I10(.SUM({ n5819_2[18:0] }), .A({ n5819[18:0] }), .B({\prod_terms[9][8] [13], 
    \prod_terms[9][8] [13], \prod_terms[9][8] [13], \prod_terms[9][8] [13], 
    \prod_terms[9][8] [13],  \prod_terms[9][8] [13:0] }));
  VDW_ADD_19_1_0 add_5819_48_I10(.SUM({ n5819[18:0] }), .A({ n5818_3[18:0] }), .B({\prod_terms[9][7] [13], 
    \prod_terms[9][7] [13], \prod_terms[9][7] [13], \prod_terms[9][7] [13], 
    \prod_terms[9][7] [13],  \prod_terms[9][7] [13:0] }));
  VDW_ADD_19_1_0 add_5818_88_I10(.SUM({ n5818_3[18:0] }), .A({ n5818_2[18:0] }), .B({\prod_terms[9][6] [13], 
    \prod_terms[9][6] [13], \prod_terms[9][6] [13], \prod_terms[9][6] [13], 
    \prod_terms[9][6] [13],  \prod_terms[9][6] [13:0] }));
  VDW_ADD_19_1_0 add_5818_68_I10(.SUM({ n5818_2[18:0] }), .A({n5818[17],  n5818[17:0] }), .B({
    \prod_terms[9][5] [13], \prod_terms[9][5] [13], \prod_terms[9][5] [13], 
    \prod_terms[9][5] [13], \prod_terms[9][5] [13],  \prod_terms[9][5] [13:0] }));
  VDW_ADD_18_1_0 add_5818_48_I10(.SUM({ n5818[17:0] }), .A({n5817_3[16],  n5817_3[16:0] }), .B({
    \prod_terms[9][4] [13], \prod_terms[9][4] [13], \prod_terms[9][4] [13], 
    \prod_terms[9][4] [13],  \prod_terms[9][4] [13:0] }));
  VDW_ADD_17_1_0 add_5817_91_I10(.SUM({ n5817_3[16:0] }), .A({n5817_2[15],  n5817_2[15:0] }), .B({
    \prod_terms[9][3] [13], \prod_terms[9][3] [13], \prod_terms[9][3] [13],  \prod_terms[9][3] [13:0] }));
  VDW_ADD_16_1_0 add_5817_71_I10(.SUM({ n5817_2[15:0] }), .A({n5817[14],  n5817[14:0] }), .B({
    \prod_terms[9][2] [13], \prod_terms[9][2] [13],  \prod_terms[9][2] [13:0] }));
  VDW_ADD_15_1_0 add_5817_52_I10(.SUM({ n5817[14:0] }), .A({\prod_terms[9][0] [13],  \prod_terms[9][0] [13:0] }), .B({
    \prod_terms[9][1] [13],  \prod_terms[9][1] [13:0] }));
  assign \b2_extended[0] [13] = \biases_l2[0] [5];
  assign \b2_extended[0] [12] = \biases_l2[0] [5];
  assign \b2_extended[0] [11] = \biases_l2[0] [5];
  assign \b2_extended[0] [10] = \biases_l2[0] [5];
  assign \b2_extended[0] [9] = \biases_l2[0] [5];
  assign \b2_extended[0] [8] = \biases_l2[0] [4];
  assign \b2_extended[0] [7] = \biases_l2[0] [3];
  assign \b2_extended[0] [6] = \biases_l2[0] [2];
  assign \b2_extended[0] [5] = \biases_l2[0] [1];
  assign \b2_extended[0] [4] = \biases_l2[0] [0];
  assign \b2_extended[1] [13] = \biases_l2[1] [5];
  assign \b2_extended[1] [12] = \biases_l2[1] [5];
  assign \b2_extended[1] [11] = \biases_l2[1] [5];
  assign \b2_extended[1] [10] = \biases_l2[1] [5];
  assign \b2_extended[1] [9] = \biases_l2[1] [5];
  assign \b2_extended[1] [8] = \biases_l2[1] [4];
  assign \b2_extended[1] [7] = \biases_l2[1] [3];
  assign \b2_extended[1] [6] = \biases_l2[1] [2];
  assign \b2_extended[1] [5] = \biases_l2[1] [1];
  assign \b2_extended[1] [4] = \biases_l2[1] [0];
  assign \b2_extended[2] [13] = \biases_l2[2] [5];
  assign \b2_extended[2] [12] = \biases_l2[2] [5];
  assign \b2_extended[2] [11] = \biases_l2[2] [5];
  assign \b2_extended[2] [10] = \biases_l2[2] [5];
  assign \b2_extended[2] [9] = \biases_l2[2] [5];
  assign \b2_extended[2] [8] = \biases_l2[2] [4];
  assign \b2_extended[2] [7] = \biases_l2[2] [3];
  assign \b2_extended[2] [6] = \biases_l2[2] [2];
  assign \b2_extended[2] [5] = \biases_l2[2] [1];
  assign \b2_extended[2] [4] = \biases_l2[2] [0];
  assign \b2_extended[3] [13] = \biases_l2[3] [5];
  assign \b2_extended[3] [12] = \biases_l2[3] [5];
  assign \b2_extended[3] [11] = \biases_l2[3] [5];
  assign \b2_extended[3] [10] = \biases_l2[3] [5];
  assign \b2_extended[3] [9] = \biases_l2[3] [5];
  assign \b2_extended[3] [8] = \biases_l2[3] [4];
  assign \b2_extended[3] [7] = \biases_l2[3] [3];
  assign \b2_extended[3] [6] = \biases_l2[3] [2];
  assign \b2_extended[3] [5] = \biases_l2[3] [1];
  assign \b2_extended[3] [4] = \biases_l2[3] [0];
  assign \b2_extended[4] [13] = \biases_l2[4] [5];
  assign \b2_extended[4] [12] = \biases_l2[4] [5];
  assign \b2_extended[4] [11] = \biases_l2[4] [5];
  assign \b2_extended[4] [10] = \biases_l2[4] [5];
  assign \b2_extended[4] [9] = \biases_l2[4] [5];
  assign \b2_extended[4] [8] = \biases_l2[4] [4];
  assign \b2_extended[4] [7] = \biases_l2[4] [3];
  assign \b2_extended[4] [6] = \biases_l2[4] [2];
  assign \b2_extended[4] [5] = \biases_l2[4] [1];
  assign \b2_extended[4] [4] = \biases_l2[4] [0];
  assign \b2_extended[5] [13] = \biases_l2[5] [5];
  assign \b2_extended[5] [12] = \biases_l2[5] [5];
  assign \b2_extended[5] [11] = \biases_l2[5] [5];
  assign \b2_extended[5] [10] = \biases_l2[5] [5];
  assign \b2_extended[5] [9] = \biases_l2[5] [5];
  assign \b2_extended[5] [8] = \biases_l2[5] [4];
  assign \b2_extended[5] [7] = \biases_l2[5] [3];
  assign \b2_extended[5] [6] = \biases_l2[5] [2];
  assign \b2_extended[5] [5] = \biases_l2[5] [1];
  assign \b2_extended[5] [4] = \biases_l2[5] [0];
  assign \b2_extended[6] [13] = \biases_l2[6] [5];
  assign \b2_extended[6] [12] = \biases_l2[6] [5];
  assign \b2_extended[6] [11] = \biases_l2[6] [5];
  assign \b2_extended[6] [10] = \biases_l2[6] [5];
  assign \b2_extended[6] [9] = \biases_l2[6] [5];
  assign \b2_extended[6] [8] = \biases_l2[6] [4];
  assign \b2_extended[6] [7] = \biases_l2[6] [3];
  assign \b2_extended[6] [6] = \biases_l2[6] [2];
  assign \b2_extended[6] [5] = \biases_l2[6] [1];
  assign \b2_extended[6] [4] = \biases_l2[6] [0];
  assign \b2_extended[7] [13] = \biases_l2[7] [5];
  assign \b2_extended[7] [12] = \biases_l2[7] [5];
  assign \b2_extended[7] [11] = \biases_l2[7] [5];
  assign \b2_extended[7] [10] = \biases_l2[7] [5];
  assign \b2_extended[7] [9] = \biases_l2[7] [5];
  assign \b2_extended[7] [8] = \biases_l2[7] [4];
  assign \b2_extended[7] [7] = \biases_l2[7] [3];
  assign \b2_extended[7] [6] = \biases_l2[7] [2];
  assign \b2_extended[7] [5] = \biases_l2[7] [1];
  assign \b2_extended[7] [4] = \biases_l2[7] [0];
  assign \b2_extended[8] [13] = \biases_l2[8] [5];
  assign \b2_extended[8] [12] = \biases_l2[8] [5];
  assign \b2_extended[8] [11] = \biases_l2[8] [5];
  assign \b2_extended[8] [10] = \biases_l2[8] [5];
  assign \b2_extended[8] [9] = \biases_l2[8] [5];
  assign \b2_extended[8] [8] = \biases_l2[8] [4];
  assign \b2_extended[8] [7] = \biases_l2[8] [3];
  assign \b2_extended[8] [6] = \biases_l2[8] [2];
  assign \b2_extended[8] [5] = \biases_l2[8] [1];
  assign \b2_extended[8] [4] = \biases_l2[8] [0];
  assign \b2_extended[9] [13] = \biases_l2[9] [5];
  assign \b2_extended[9] [12] = \biases_l2[9] [5];
  assign \b2_extended[9] [11] = \biases_l2[9] [5];
  assign \b2_extended[9] [10] = \biases_l2[9] [5];
  assign \b2_extended[9] [9] = \biases_l2[9] [5];
  assign \b2_extended[9] [8] = \biases_l2[9] [4];
  assign \b2_extended[9] [7] = \biases_l2[9] [3];
  assign \b2_extended[9] [6] = \biases_l2[9] [2];
  assign \b2_extended[9] [5] = \biases_l2[9] [1];
  assign \b2_extended[9] [4] = \biases_l2[9] [0];
  assign out[179] = \out_reg[9] [17];
  assign out[178] = \out_reg[9] [16];
  assign out[177] = \out_reg[9] [15];
  assign out[176] = \out_reg[9] [14];
  assign out[175] = \out_reg[9] [13];
  assign out[174] = \out_reg[9] [12];
  assign out[173] = \out_reg[9] [11];
  assign out[172] = \out_reg[9] [10];
  assign out[171] = \out_reg[9] [9];
  assign out[170] = \out_reg[9] [8];
  assign out[169] = \out_reg[9] [7];
  assign out[168] = \out_reg[9] [6];
  assign out[167] = \out_reg[9] [5];
  assign out[166] = \out_reg[9] [4];
  assign out[165] = \out_reg[9] [3];
  assign out[164] = \out_reg[9] [2];
  assign out[163] = \out_reg[9] [1];
  assign out[162] = \out_reg[9] [0];
  assign out[161] = \out_reg[8] [17];
  assign out[160] = \out_reg[8] [16];
  assign out[159] = \out_reg[8] [15];
  assign out[158] = \out_reg[8] [14];
  assign out[157] = \out_reg[8] [13];
  assign out[156] = \out_reg[8] [12];
  assign out[155] = \out_reg[8] [11];
  assign out[154] = \out_reg[8] [10];
  assign out[153] = \out_reg[8] [9];
  assign out[152] = \out_reg[8] [8];
  assign out[151] = \out_reg[8] [7];
  assign out[150] = \out_reg[8] [6];
  assign out[149] = \out_reg[8] [5];
  assign out[148] = \out_reg[8] [4];
  assign out[147] = \out_reg[8] [3];
  assign out[146] = \out_reg[8] [2];
  assign out[145] = \out_reg[8] [1];
  assign out[144] = \out_reg[8] [0];
  assign out[143] = \out_reg[7] [17];
  assign out[142] = \out_reg[7] [16];
  assign out[141] = \out_reg[7] [15];
  assign out[140] = \out_reg[7] [14];
  assign out[139] = \out_reg[7] [13];
  assign out[138] = \out_reg[7] [12];
  assign out[137] = \out_reg[7] [11];
  assign out[136] = \out_reg[7] [10];
  assign out[135] = \out_reg[7] [9];
  assign out[134] = \out_reg[7] [8];
  assign out[133] = \out_reg[7] [7];
  assign out[132] = \out_reg[7] [6];
  assign out[131] = \out_reg[7] [5];
  assign out[130] = \out_reg[7] [4];
  assign out[129] = \out_reg[7] [3];
  assign out[128] = \out_reg[7] [2];
  assign out[127] = \out_reg[7] [1];
  assign out[126] = \out_reg[7] [0];
  assign out[125] = \out_reg[6] [17];
  assign out[124] = \out_reg[6] [16];
  assign out[123] = \out_reg[6] [15];
  assign out[122] = \out_reg[6] [14];
  assign out[121] = \out_reg[6] [13];
  assign out[120] = \out_reg[6] [12];
  assign out[119] = \out_reg[6] [11];
  assign out[118] = \out_reg[6] [10];
  assign out[117] = \out_reg[6] [9];
  assign out[116] = \out_reg[6] [8];
  assign out[115] = \out_reg[6] [7];
  assign out[114] = \out_reg[6] [6];
  assign out[113] = \out_reg[6] [5];
  assign out[112] = \out_reg[6] [4];
  assign out[111] = \out_reg[6] [3];
  assign out[110] = \out_reg[6] [2];
  assign out[109] = \out_reg[6] [1];
  assign out[108] = \out_reg[6] [0];
  assign out[107] = \out_reg[5] [17];
  assign out[106] = \out_reg[5] [16];
  assign out[105] = \out_reg[5] [15];
  assign out[104] = \out_reg[5] [14];
  assign out[103] = \out_reg[5] [13];
  assign out[102] = \out_reg[5] [12];
  assign out[101] = \out_reg[5] [11];
  assign out[100] = \out_reg[5] [10];
  assign out[99] = \out_reg[5] [9];
  assign out[98] = \out_reg[5] [8];
  assign out[97] = \out_reg[5] [7];
  assign out[96] = \out_reg[5] [6];
  assign out[95] = \out_reg[5] [5];
  assign out[94] = \out_reg[5] [4];
  assign out[93] = \out_reg[5] [3];
  assign out[92] = \out_reg[5] [2];
  assign out[91] = \out_reg[5] [1];
  assign out[90] = \out_reg[5] [0];
  assign out[89] = \out_reg[4] [17];
  assign out[88] = \out_reg[4] [16];
  assign out[87] = \out_reg[4] [15];
  assign out[86] = \out_reg[4] [14];
  assign out[85] = \out_reg[4] [13];
  assign out[84] = \out_reg[4] [12];
  assign out[83] = \out_reg[4] [11];
  assign out[82] = \out_reg[4] [10];
  assign out[81] = \out_reg[4] [9];
  assign out[80] = \out_reg[4] [8];
  assign out[79] = \out_reg[4] [7];
  assign out[78] = \out_reg[4] [6];
  assign out[77] = \out_reg[4] [5];
  assign out[76] = \out_reg[4] [4];
  assign out[75] = \out_reg[4] [3];
  assign out[74] = \out_reg[4] [2];
  assign out[73] = \out_reg[4] [1];
  assign out[72] = \out_reg[4] [0];
  assign out[71] = \out_reg[3] [17];
  assign out[70] = \out_reg[3] [16];
  assign out[69] = \out_reg[3] [15];
  assign out[68] = \out_reg[3] [14];
  assign out[67] = \out_reg[3] [13];
  assign out[66] = \out_reg[3] [12];
  assign out[65] = \out_reg[3] [11];
  assign out[64] = \out_reg[3] [10];
  assign out[63] = \out_reg[3] [9];
  assign out[62] = \out_reg[3] [8];
  assign out[61] = \out_reg[3] [7];
  assign out[60] = \out_reg[3] [6];
  assign out[59] = \out_reg[3] [5];
  assign out[58] = \out_reg[3] [4];
  assign out[57] = \out_reg[3] [3];
  assign out[56] = \out_reg[3] [2];
  assign out[55] = \out_reg[3] [1];
  assign out[54] = \out_reg[3] [0];
  assign out[53] = \out_reg[2] [17];
  assign out[52] = \out_reg[2] [16];
  assign out[51] = \out_reg[2] [15];
  assign out[50] = \out_reg[2] [14];
  assign out[49] = \out_reg[2] [13];
  assign out[48] = \out_reg[2] [12];
  assign out[47] = \out_reg[2] [11];
  assign out[46] = \out_reg[2] [10];
  assign out[45] = \out_reg[2] [9];
  assign out[44] = \out_reg[2] [8];
  assign out[43] = \out_reg[2] [7];
  assign out[42] = \out_reg[2] [6];
  assign out[41] = \out_reg[2] [5];
  assign out[40] = \out_reg[2] [4];
  assign out[39] = \out_reg[2] [3];
  assign out[38] = \out_reg[2] [2];
  assign out[37] = \out_reg[2] [1];
  assign out[36] = \out_reg[2] [0];
  assign out[35] = \out_reg[1] [17];
  assign out[34] = \out_reg[1] [16];
  assign out[33] = \out_reg[1] [15];
  assign out[32] = \out_reg[1] [14];
  assign out[31] = \out_reg[1] [13];
  assign out[30] = \out_reg[1] [12];
  assign out[29] = \out_reg[1] [11];
  assign out[28] = \out_reg[1] [10];
  assign out[27] = \out_reg[1] [9];
  assign out[26] = \out_reg[1] [8];
  assign out[25] = \out_reg[1] [7];
  assign out[24] = \out_reg[1] [6];
  assign out[23] = \out_reg[1] [5];
  assign out[22] = \out_reg[1] [4];
  assign out[21] = \out_reg[1] [3];
  assign out[20] = \out_reg[1] [2];
  assign out[19] = \out_reg[1] [1];
  assign out[18] = \out_reg[1] [0];
  assign out[17] = \out_reg[0] [17];
  assign out[16] = \out_reg[0] [16];
  assign out[15] = \out_reg[0] [15];
  assign out[14] = \out_reg[0] [14];
  assign out[13] = \out_reg[0] [13];
  assign out[12] = \out_reg[0] [12];
  assign out[11] = \out_reg[0] [11];
  assign out[10] = \out_reg[0] [10];
  assign out[9] = \out_reg[0] [9];
  assign out[8] = \out_reg[0] [8];
  assign out[7] = \out_reg[0] [7];
  assign out[6] = \out_reg[0] [6];
  assign out[5] = \out_reg[0] [5];
  assign out[4] = \out_reg[0] [4];
  assign out[3] = \out_reg[0] [3];
  assign out[2] = \out_reg[0] [2];
  assign out[1] = \out_reg[0] [1];
  assign out[0] = \out_reg[0] [0];
  ReLU_19bit \row_iteration[0].relu_inst (.in_data({ \row_sums[0] [18:0] }), .out_data({ \row_output[0] [17:0] }));
  multiplier9514 \row_iteration[0].prod_calc[0].mult_inst (.prod({ \prod_terms[0][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[0][0] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[1].mult_inst (.prod({ \prod_terms[0][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[0][1] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[2].mult_inst (.prod({ \prod_terms[0][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[0][2] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[3].mult_inst (.prod({ \prod_terms[0][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[0][3] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[4].mult_inst (.prod({ \prod_terms[0][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[0][4] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[5].mult_inst (.prod({ \prod_terms[0][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[0][5] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[6].mult_inst (.prod({ \prod_terms[0][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[0][6] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[7].mult_inst (.prod({ \prod_terms[0][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[0][7] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[8].mult_inst (.prod({ \prod_terms[0][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[0][8] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[9].mult_inst (.prod({ \prod_terms[0][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[0][9] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[10].mult_inst (.prod({ \prod_terms[0][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[0][10] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[11].mult_inst (.prod({ \prod_terms[0][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[0][11] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[12].mult_inst (.prod({ \prod_terms[0][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[0][12] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[13].mult_inst (.prod({ \prod_terms[0][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[0][13] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[14].mult_inst (.prod({ \prod_terms[0][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[0][14] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[15].mult_inst (.prod({ \prod_terms[0][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[0][15] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[16].mult_inst (.prod({ \prod_terms[0][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[0][16] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[17].mult_inst (.prod({ \prod_terms[0][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[0][17] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[18].mult_inst (.prod({ \prod_terms[0][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[0][18] [4:0] }));
  multiplier9514 \row_iteration[0].prod_calc[19].mult_inst (.prod({ \prod_terms[0][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[0][19] [4:0] }));
  ReLU_19bit \row_iteration[1].relu_inst (.in_data({ \row_sums[1] [18:0] }), .out_data({ \row_output[1] [17:0] }));
  multiplier9514 \row_iteration[1].prod_calc[0].mult_inst (.prod({ \prod_terms[1][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[1][0] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[1].mult_inst (.prod({ \prod_terms[1][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[1][1] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[2].mult_inst (.prod({ \prod_terms[1][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[1][2] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[3].mult_inst (.prod({ \prod_terms[1][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[1][3] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[4].mult_inst (.prod({ \prod_terms[1][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[1][4] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[5].mult_inst (.prod({ \prod_terms[1][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[1][5] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[6].mult_inst (.prod({ \prod_terms[1][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[1][6] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[7].mult_inst (.prod({ \prod_terms[1][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[1][7] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[8].mult_inst (.prod({ \prod_terms[1][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[1][8] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[9].mult_inst (.prod({ \prod_terms[1][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[1][9] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[10].mult_inst (.prod({ \prod_terms[1][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[1][10] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[11].mult_inst (.prod({ \prod_terms[1][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[1][11] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[12].mult_inst (.prod({ \prod_terms[1][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[1][12] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[13].mult_inst (.prod({ \prod_terms[1][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[1][13] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[14].mult_inst (.prod({ \prod_terms[1][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[1][14] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[15].mult_inst (.prod({ \prod_terms[1][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[1][15] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[16].mult_inst (.prod({ \prod_terms[1][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[1][16] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[17].mult_inst (.prod({ \prod_terms[1][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[1][17] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[18].mult_inst (.prod({ \prod_terms[1][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[1][18] [4:0] }));
  multiplier9514 \row_iteration[1].prod_calc[19].mult_inst (.prod({ \prod_terms[1][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[1][19] [4:0] }));
  ReLU_19bit \row_iteration[2].relu_inst (.in_data({ \row_sums[2] [18:0] }), .out_data({ \row_output[2] [17:0] }));
  multiplier9514 \row_iteration[2].prod_calc[0].mult_inst (.prod({ \prod_terms[2][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[2][0] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[1].mult_inst (.prod({ \prod_terms[2][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[2][1] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[2].mult_inst (.prod({ \prod_terms[2][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[2][2] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[3].mult_inst (.prod({ \prod_terms[2][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[2][3] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[4].mult_inst (.prod({ \prod_terms[2][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[2][4] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[5].mult_inst (.prod({ \prod_terms[2][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[2][5] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[6].mult_inst (.prod({ \prod_terms[2][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[2][6] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[7].mult_inst (.prod({ \prod_terms[2][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[2][7] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[8].mult_inst (.prod({ \prod_terms[2][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[2][8] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[9].mult_inst (.prod({ \prod_terms[2][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[2][9] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[10].mult_inst (.prod({ \prod_terms[2][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[2][10] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[11].mult_inst (.prod({ \prod_terms[2][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[2][11] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[12].mult_inst (.prod({ \prod_terms[2][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[2][12] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[13].mult_inst (.prod({ \prod_terms[2][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[2][13] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[14].mult_inst (.prod({ \prod_terms[2][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[2][14] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[15].mult_inst (.prod({ \prod_terms[2][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[2][15] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[16].mult_inst (.prod({ \prod_terms[2][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[2][16] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[17].mult_inst (.prod({ \prod_terms[2][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[2][17] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[18].mult_inst (.prod({ \prod_terms[2][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[2][18] [4:0] }));
  multiplier9514 \row_iteration[2].prod_calc[19].mult_inst (.prod({ \prod_terms[2][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[2][19] [4:0] }));
  ReLU_19bit \row_iteration[3].relu_inst (.in_data({ \row_sums[3] [18:0] }), .out_data({ \row_output[3] [17:0] }));
  multiplier9514 \row_iteration[3].prod_calc[0].mult_inst (.prod({ \prod_terms[3][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[3][0] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[1].mult_inst (.prod({ \prod_terms[3][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[3][1] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[2].mult_inst (.prod({ \prod_terms[3][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[3][2] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[3].mult_inst (.prod({ \prod_terms[3][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[3][3] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[4].mult_inst (.prod({ \prod_terms[3][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[3][4] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[5].mult_inst (.prod({ \prod_terms[3][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[3][5] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[6].mult_inst (.prod({ \prod_terms[3][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[3][6] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[7].mult_inst (.prod({ \prod_terms[3][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[3][7] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[8].mult_inst (.prod({ \prod_terms[3][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[3][8] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[9].mult_inst (.prod({ \prod_terms[3][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[3][9] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[10].mult_inst (.prod({ \prod_terms[3][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[3][10] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[11].mult_inst (.prod({ \prod_terms[3][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[3][11] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[12].mult_inst (.prod({ \prod_terms[3][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[3][12] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[13].mult_inst (.prod({ \prod_terms[3][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[3][13] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[14].mult_inst (.prod({ \prod_terms[3][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[3][14] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[15].mult_inst (.prod({ \prod_terms[3][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[3][15] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[16].mult_inst (.prod({ \prod_terms[3][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[3][16] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[17].mult_inst (.prod({ \prod_terms[3][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[3][17] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[18].mult_inst (.prod({ \prod_terms[3][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[3][18] [4:0] }));
  multiplier9514 \row_iteration[3].prod_calc[19].mult_inst (.prod({ \prod_terms[3][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[3][19] [4:0] }));
  ReLU_19bit \row_iteration[4].relu_inst (.in_data({ \row_sums[4] [18:0] }), .out_data({ \row_output[4] [17:0] }));
  multiplier9514 \row_iteration[4].prod_calc[0].mult_inst (.prod({ \prod_terms[4][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[4][0] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[1].mult_inst (.prod({ \prod_terms[4][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[4][1] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[2].mult_inst (.prod({ \prod_terms[4][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[4][2] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[3].mult_inst (.prod({ \prod_terms[4][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[4][3] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[4].mult_inst (.prod({ \prod_terms[4][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[4][4] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[5].mult_inst (.prod({ \prod_terms[4][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[4][5] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[6].mult_inst (.prod({ \prod_terms[4][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[4][6] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[7].mult_inst (.prod({ \prod_terms[4][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[4][7] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[8].mult_inst (.prod({ \prod_terms[4][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[4][8] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[9].mult_inst (.prod({ \prod_terms[4][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[4][9] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[10].mult_inst (.prod({ \prod_terms[4][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[4][10] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[11].mult_inst (.prod({ \prod_terms[4][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[4][11] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[12].mult_inst (.prod({ \prod_terms[4][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[4][12] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[13].mult_inst (.prod({ \prod_terms[4][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[4][13] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[14].mult_inst (.prod({ \prod_terms[4][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[4][14] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[15].mult_inst (.prod({ \prod_terms[4][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[4][15] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[16].mult_inst (.prod({ \prod_terms[4][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[4][16] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[17].mult_inst (.prod({ \prod_terms[4][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[4][17] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[18].mult_inst (.prod({ \prod_terms[4][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[4][18] [4:0] }));
  multiplier9514 \row_iteration[4].prod_calc[19].mult_inst (.prod({ \prod_terms[4][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[4][19] [4:0] }));
  ReLU_19bit \row_iteration[5].relu_inst (.in_data({ \row_sums[5] [18:0] }), .out_data({ \row_output[5] [17:0] }));
  multiplier9514 \row_iteration[5].prod_calc[0].mult_inst (.prod({ \prod_terms[5][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[5][0] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[1].mult_inst (.prod({ \prod_terms[5][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[5][1] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[2].mult_inst (.prod({ \prod_terms[5][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[5][2] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[3].mult_inst (.prod({ \prod_terms[5][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[5][3] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[4].mult_inst (.prod({ \prod_terms[5][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[5][4] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[5].mult_inst (.prod({ \prod_terms[5][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[5][5] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[6].mult_inst (.prod({ \prod_terms[5][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[5][6] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[7].mult_inst (.prod({ \prod_terms[5][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[5][7] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[8].mult_inst (.prod({ \prod_terms[5][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[5][8] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[9].mult_inst (.prod({ \prod_terms[5][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[5][9] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[10].mult_inst (.prod({ \prod_terms[5][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[5][10] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[11].mult_inst (.prod({ \prod_terms[5][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[5][11] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[12].mult_inst (.prod({ \prod_terms[5][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[5][12] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[13].mult_inst (.prod({ \prod_terms[5][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[5][13] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[14].mult_inst (.prod({ \prod_terms[5][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[5][14] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[15].mult_inst (.prod({ \prod_terms[5][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[5][15] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[16].mult_inst (.prod({ \prod_terms[5][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[5][16] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[17].mult_inst (.prod({ \prod_terms[5][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[5][17] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[18].mult_inst (.prod({ \prod_terms[5][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[5][18] [4:0] }));
  multiplier9514 \row_iteration[5].prod_calc[19].mult_inst (.prod({ \prod_terms[5][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[5][19] [4:0] }));
  ReLU_19bit \row_iteration[6].relu_inst (.in_data({ \row_sums[6] [18:0] }), .out_data({ \row_output[6] [17:0] }));
  multiplier9514 \row_iteration[6].prod_calc[0].mult_inst (.prod({ \prod_terms[6][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[6][0] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[1].mult_inst (.prod({ \prod_terms[6][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[6][1] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[2].mult_inst (.prod({ \prod_terms[6][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[6][2] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[3].mult_inst (.prod({ \prod_terms[6][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[6][3] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[4].mult_inst (.prod({ \prod_terms[6][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[6][4] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[5].mult_inst (.prod({ \prod_terms[6][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[6][5] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[6].mult_inst (.prod({ \prod_terms[6][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[6][6] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[7].mult_inst (.prod({ \prod_terms[6][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[6][7] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[8].mult_inst (.prod({ \prod_terms[6][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[6][8] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[9].mult_inst (.prod({ \prod_terms[6][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[6][9] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[10].mult_inst (.prod({ \prod_terms[6][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[6][10] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[11].mult_inst (.prod({ \prod_terms[6][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[6][11] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[12].mult_inst (.prod({ \prod_terms[6][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[6][12] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[13].mult_inst (.prod({ \prod_terms[6][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[6][13] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[14].mult_inst (.prod({ \prod_terms[6][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[6][14] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[15].mult_inst (.prod({ \prod_terms[6][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[6][15] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[16].mult_inst (.prod({ \prod_terms[6][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[6][16] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[17].mult_inst (.prod({ \prod_terms[6][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[6][17] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[18].mult_inst (.prod({ \prod_terms[6][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[6][18] [4:0] }));
  multiplier9514 \row_iteration[6].prod_calc[19].mult_inst (.prod({ \prod_terms[6][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[6][19] [4:0] }));
  ReLU_19bit \row_iteration[7].relu_inst (.in_data({ \row_sums[7] [18:0] }), .out_data({ \row_output[7] [17:0] }));
  multiplier9514 \row_iteration[7].prod_calc[0].mult_inst (.prod({ \prod_terms[7][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[7][0] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[1].mult_inst (.prod({ \prod_terms[7][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[7][1] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[2].mult_inst (.prod({ \prod_terms[7][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[7][2] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[3].mult_inst (.prod({ \prod_terms[7][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[7][3] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[4].mult_inst (.prod({ \prod_terms[7][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[7][4] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[5].mult_inst (.prod({ \prod_terms[7][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[7][5] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[6].mult_inst (.prod({ \prod_terms[7][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[7][6] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[7].mult_inst (.prod({ \prod_terms[7][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[7][7] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[8].mult_inst (.prod({ \prod_terms[7][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[7][8] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[9].mult_inst (.prod({ \prod_terms[7][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[7][9] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[10].mult_inst (.prod({ \prod_terms[7][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[7][10] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[11].mult_inst (.prod({ \prod_terms[7][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[7][11] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[12].mult_inst (.prod({ \prod_terms[7][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[7][12] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[13].mult_inst (.prod({ \prod_terms[7][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[7][13] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[14].mult_inst (.prod({ \prod_terms[7][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[7][14] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[15].mult_inst (.prod({ \prod_terms[7][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[7][15] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[16].mult_inst (.prod({ \prod_terms[7][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[7][16] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[17].mult_inst (.prod({ \prod_terms[7][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[7][17] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[18].mult_inst (.prod({ \prod_terms[7][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[7][18] [4:0] }));
  multiplier9514 \row_iteration[7].prod_calc[19].mult_inst (.prod({ \prod_terms[7][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[7][19] [4:0] }));
  ReLU_19bit \row_iteration[8].relu_inst (.in_data({ \row_sums[8] [18:0] }), .out_data({ \row_output[8] [17:0] }));
  multiplier9514 \row_iteration[8].prod_calc[0].mult_inst (.prod({ \prod_terms[8][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[8][0] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[1].mult_inst (.prod({ \prod_terms[8][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[8][1] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[2].mult_inst (.prod({ \prod_terms[8][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[8][2] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[3].mult_inst (.prod({ \prod_terms[8][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[8][3] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[4].mult_inst (.prod({ \prod_terms[8][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[8][4] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[5].mult_inst (.prod({ \prod_terms[8][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[8][5] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[6].mult_inst (.prod({ \prod_terms[8][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[8][6] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[7].mult_inst (.prod({ \prod_terms[8][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[8][7] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[8].mult_inst (.prod({ \prod_terms[8][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[8][8] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[9].mult_inst (.prod({ \prod_terms[8][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[8][9] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[10].mult_inst (.prod({ \prod_terms[8][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[8][10] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[11].mult_inst (.prod({ \prod_terms[8][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[8][11] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[12].mult_inst (.prod({ \prod_terms[8][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[8][12] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[13].mult_inst (.prod({ \prod_terms[8][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[8][13] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[14].mult_inst (.prod({ \prod_terms[8][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[8][14] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[15].mult_inst (.prod({ \prod_terms[8][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[8][15] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[16].mult_inst (.prod({ \prod_terms[8][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[8][16] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[17].mult_inst (.prod({ \prod_terms[8][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[8][17] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[18].mult_inst (.prod({ \prod_terms[8][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[8][18] [4:0] }));
  multiplier9514 \row_iteration[8].prod_calc[19].mult_inst (.prod({ \prod_terms[8][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[8][19] [4:0] }));
  ReLU_19bit \row_iteration[9].relu_inst (.in_data({ \row_sums[9] [18:0] }), .out_data({ \row_output[9] [17:0] }));
  multiplier9514 \row_iteration[9].prod_calc[0].mult_inst (.prod({ \prod_terms[9][0] [13:0] }), .num1({ in[8:0] }),
     .num2({ \w2[9][0] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[1].mult_inst (.prod({ \prod_terms[9][1] [13:0] }), .num1({ in[17:9] }),
     .num2({ \w2[9][1] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[2].mult_inst (.prod({ \prod_terms[9][2] [13:0] }), .num1({ in[26:18] }),
     .num2({ \w2[9][2] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[3].mult_inst (.prod({ \prod_terms[9][3] [13:0] }), .num1({ in[35:27] }),
     .num2({ \w2[9][3] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[4].mult_inst (.prod({ \prod_terms[9][4] [13:0] }), .num1({ in[44:36] }),
     .num2({ \w2[9][4] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[5].mult_inst (.prod({ \prod_terms[9][5] [13:0] }), .num1({ in[53:45] }),
     .num2({ \w2[9][5] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[6].mult_inst (.prod({ \prod_terms[9][6] [13:0] }), .num1({ in[62:54] }),
     .num2({ \w2[9][6] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[7].mult_inst (.prod({ \prod_terms[9][7] [13:0] }), .num1({ in[71:63] }),
     .num2({ \w2[9][7] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[8].mult_inst (.prod({ \prod_terms[9][8] [13:0] }), .num1({ in[80:72] }),
     .num2({ \w2[9][8] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[9].mult_inst (.prod({ \prod_terms[9][9] [13:0] }), .num1({ in[89:81] }),
     .num2({ \w2[9][9] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[10].mult_inst (.prod({ \prod_terms[9][10] [13:0] }), .num1({ in[98:90] }),
     .num2({ \w2[9][10] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[11].mult_inst (.prod({ \prod_terms[9][11] [13:0] }), .num1({ in[107:99] }),
     .num2({ \w2[9][11] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[12].mult_inst (.prod({ \prod_terms[9][12] [13:0] }), .num1({ in[116:108] }),
     .num2({ \w2[9][12] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[13].mult_inst (.prod({ \prod_terms[9][13] [13:0] }), .num1({ in[125:117] }),
     .num2({ \w2[9][13] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[14].mult_inst (.prod({ \prod_terms[9][14] [13:0] }), .num1({ in[134:126] }),
     .num2({ \w2[9][14] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[15].mult_inst (.prod({ \prod_terms[9][15] [13:0] }), .num1({ in[143:135] }),
     .num2({ \w2[9][15] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[16].mult_inst (.prod({ \prod_terms[9][16] [13:0] }), .num1({ in[152:144] }),
     .num2({ \w2[9][16] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[17].mult_inst (.prod({ \prod_terms[9][17] [13:0] }), .num1({ in[161:153] }),
     .num2({ \w2[9][17] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[18].mult_inst (.prod({ \prod_terms[9][18] [13:0] }), .num1({ in[170:162] }),
     .num2({ \w2[9][18] [4:0] }));
  multiplier9514 \row_iteration[9].prod_calc[19].mult_inst (.prod({ \prod_terms[9][19] [13:0] }), .num1({ in[179:171] }),
     .num2({ \w2[9][19] [4:0] }));
endmodule

module VDW_WMUX4 (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX4_CIM_4 (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX4_CIM_3 (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX4_CIM_2 (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX4_CIM_1 (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_WMUX4_CIM (Z, A, B, S);
// conformal library_module
output [3:0] Z;
input [3:0] A, B;
input S;
  assign Z = S ? B : A;
endmodule

module VDW_GT_u18(Z, A, B);
// conformal library_module
output Z;
input   [17:0] A;
input   [17:0] B;
wire  N$1, N$2, N$3, N$4, N$5, N$6, N$7, N$8, N$9, N$10, N$11, N$12, N$13, N$14, 
    N$15, N$16, N$17, N$18, N$19, N$20, N$21, N$22, N$23, N$24, N$25, N$26, 
    N$27, N$28, N$29, N$30, N$31, N$32, N$33, N$34, N$35, N$36, N$37, N$38, 
    N$39, N$40, N$41, N$42, N$43, N$44, N$45, N$46, N$47, N$48, N$49, N$50, 
    N$51, N$52, N$53, N$54, N$55, N$56, N$57, N$58, N$59, N$60, N$61, N$62, 
    N$63, N$64, N$65, N$66, N$67, N$68, N$69, N$70, N$71, N$72, N$73, N$74, 
    N$75, N$76, N$77, N$78, N$79, N$80, N$81, N$82, N$83, N$84, N$85, N$86, Z;
wire   [17:0] B;
wire   [17:0] A;
  or U$1(Z, N$2, N$1);
  and U$2(N$1, N$4, N$3);
  xnor U$3(N$3, A[17], B[17]);
  and U$4(N$2, N$5, A[17]);
  not U$5(N$5, B[17]);
  or U$6(N$4, N$7, N$6);
  and U$7(N$6, N$9, N$8);
  xnor U$8(N$8, A[16], B[16]);
  and U$9(N$7, N$10, A[16]);
  not U$10(N$10, B[16]);
  or U$11(N$9, N$12, N$11);
  and U$12(N$11, N$14, N$13);
  xnor U$13(N$13, A[15], B[15]);
  and U$14(N$12, N$15, A[15]);
  not U$15(N$15, B[15]);
  or U$16(N$14, N$17, N$16);
  and U$17(N$16, N$19, N$18);
  xnor U$18(N$18, A[14], B[14]);
  and U$19(N$17, N$20, A[14]);
  not U$20(N$20, B[14]);
  or U$21(N$19, N$22, N$21);
  and U$22(N$21, N$24, N$23);
  xnor U$23(N$23, A[13], B[13]);
  and U$24(N$22, N$25, A[13]);
  not U$25(N$25, B[13]);
  or U$26(N$24, N$27, N$26);
  and U$27(N$26, N$29, N$28);
  xnor U$28(N$28, A[12], B[12]);
  and U$29(N$27, N$30, A[12]);
  not U$30(N$30, B[12]);
  or U$31(N$29, N$32, N$31);
  and U$32(N$31, N$34, N$33);
  xnor U$33(N$33, A[11], B[11]);
  and U$34(N$32, N$35, A[11]);
  not U$35(N$35, B[11]);
  or U$36(N$34, N$37, N$36);
  and U$37(N$36, N$39, N$38);
  xnor U$38(N$38, A[10], B[10]);
  and U$39(N$37, N$40, A[10]);
  not U$40(N$40, B[10]);
  or U$41(N$39, N$42, N$41);
  and U$42(N$41, N$44, N$43);
  xnor U$43(N$43, A[9], B[9]);
  and U$44(N$42, N$45, A[9]);
  not U$45(N$45, B[9]);
  or U$46(N$44, N$47, N$46);
  and U$47(N$46, N$49, N$48);
  xnor U$48(N$48, A[8], B[8]);
  and U$49(N$47, N$50, A[8]);
  not U$50(N$50, B[8]);
  or U$51(N$49, N$52, N$51);
  and U$52(N$51, N$54, N$53);
  xnor U$53(N$53, A[7], B[7]);
  and U$54(N$52, N$55, A[7]);
  not U$55(N$55, B[7]);
  or U$56(N$54, N$57, N$56);
  and U$57(N$56, N$59, N$58);
  xnor U$58(N$58, A[6], B[6]);
  and U$59(N$57, N$60, A[6]);
  not U$60(N$60, B[6]);
  or U$61(N$59, N$62, N$61);
  and U$62(N$61, N$64, N$63);
  xnor U$63(N$63, A[5], B[5]);
  and U$64(N$62, N$65, A[5]);
  not U$65(N$65, B[5]);
  or U$66(N$64, N$67, N$66);
  and U$67(N$66, N$69, N$68);
  xnor U$68(N$68, A[4], B[4]);
  and U$69(N$67, N$70, A[4]);
  not U$70(N$70, B[4]);
  or U$71(N$69, N$72, N$71);
  and U$72(N$71, N$74, N$73);
  xnor U$73(N$73, A[3], B[3]);
  and U$74(N$72, N$75, A[3]);
  not U$75(N$75, B[3]);
  or U$76(N$74, N$77, N$76);
  and U$77(N$76, N$79, N$78);
  xnor U$78(N$78, A[2], B[2]);
  and U$79(N$77, N$80, A[2]);
  not U$80(N$80, B[2]);
  or U$81(N$79, N$82, N$81);
  and U$82(N$81, N$84, N$83);
  xnor U$83(N$83, A[1], B[1]);
  and U$84(N$82, N$85, A[1]);
  not U$85(N$85, B[1]);
  and U$86(N$84, N$86, A[0]);
  not U$87(N$86, B[0]);
endmodule

module compare_n_out(a, b, max);
output max;
input   [17:0] a;
input   [17:0] b;
wire  max;
wire   [17:0] b;
wire   [17:0] a;
  VDW_GT_u18 gt_57_21(.Z(max), .A({ a[17:0] }), .B({ b[17:0] }));
endmodule

module find_max_index(data_in, clk, rst_n, max_index, max_value);
input  clk, rst_n;
input   [179:0] data_in;
output  [3:0] max_index;
output  [17:0] max_value;
wire  n132, \stage3[0].gt , \stage2[1].gt , \stage2[0].gt , \stage1[4].gt , 
    \stage1[3].gt , \stage1[2].gt , \stage1[1].gt , \stage1[0].gt , gt_final, 
    rst_n, clk;
wire  N$1, N$2, N$3, N$4;
wire   [3:0] final_index;
wire   [3:0] \stage3_indices[0] ;
wire   [3:0] \stage3_indices[1] ;
wire   [3:0] \stage2_indices[0] ;
wire   [3:0] \stage2_indices[1] ;
wire   [3:0] \stage2_indices[2] ;
wire   [3:0] \stage1_indices[0] ;
wire   [3:0] \stage1_indices[1] ;
wire   [3:0] \stage1_indices[2] ;
wire   [3:0] \stage1_indices[3] ;
wire   [3:0] \stage1_indices[4] ;
wire   [17:0] final_winner;
wire   [17:0] \stage3_winners[0] ;
wire   [17:0] \stage3_winners[1] ;
wire   [17:0] \stage2_winners[0] ;
wire   [17:0] \stage2_winners[1] ;
wire   [17:0] \stage2_winners[2] ;
wire   [17:0] \stage1_winners[0] ;
wire   [17:0] \stage1_winners[1] ;
wire   [17:0] \stage1_winners[2] ;
wire   [17:0] \stage1_winners[3] ;
wire   [17:0] \stage1_winners[4] ;
wire   [17:0] max_value;
wire   [3:0] max_index;
wire   [179:0] data_in;
  assign N$1 = 1'b0;
  assign N$2 = 1'b0;
  assign N$3 = 1'b0;
  assign N$4 = 1'b0;
  assign \stage1_indices[0] [3] = 1'b0;
  assign \stage1_indices[0] [2] = 1'b0;
  assign \stage1_indices[0] [1] = 1'b0;
  assign \stage1_indices[1] [3] = 1'b0;
  assign \stage1_indices[1] [2] = 1'b0;
  assign \stage1_indices[2] [3] = 1'b0;
  assign \stage1_indices[2] [1] = 1'b0;
  assign \stage1_indices[3] [3] = 1'b0;
  assign \stage1_indices[4] [2] = 1'b0;
  assign \stage1_indices[4] [1] = 1'b0;
  assign \stage1_indices[1] [1] = 1'b1;
  assign \stage1_indices[2] [2] = 1'b1;
  assign \stage1_indices[3] [2] = 1'b1;
  assign \stage1_indices[3] [1] = 1'b1;
  assign \stage1_indices[4] [3] = 1'b1;
  VDW_WMUX4 U$1(.Z({ final_index[3:0] }), .A({ \stage3_indices[1] [3:0] }), .B({ \stage3_indices[0] [3:0] }), .S(gt_final));
  VDW_WMUX4 U$2(.Z({ \stage3_indices[0] [3:0] }), .A({ \stage2_indices[0] [3:0] }), .B({ \stage2_indices[1] [3:0] }), .S(\stage3[0].gt ));
  assign \stage3_indices[1] [3] = \stage2_indices[2] [3];
  assign \stage3_indices[1] [2] = \stage2_indices[2] [2];
  assign \stage3_indices[1] [1] = \stage2_indices[2] [1];
  assign \stage3_indices[1] [0] = \stage2_indices[2] [0];
  VDW_WMUX4 U$7(.Z({ \stage2_indices[0] [3:0] }), .A({ \stage1_indices[0] [3:0] }), .B({ \stage1_indices[1] [3:0] }), .S(\stage2[0].gt ));
  VDW_WMUX4 U$8(.Z({ \stage2_indices[1] [3:0] }), .A({ \stage1_indices[2] [3:0] }), .B({ \stage1_indices[3] [3:0] }), .S(\stage2[1].gt ));
  assign \stage2_indices[2] [3] = \stage1_indices[4] [3];
  assign \stage2_indices[2] [2] = \stage1_indices[4] [2];
  assign \stage2_indices[2] [1] = \stage1_indices[4] [1];
  assign \stage2_indices[2] [0] = \stage1_indices[4] [0];
  VDW_WMUX4_CIM_4 U$13(.Z({dummy$0, dummy$1, dummy$2, \stage1_indices[0] [0]}),
     .A({1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b1}), .S(
    \stage1[0].gt ));
  VDW_WMUX4_CIM_3 U$14(.Z({dummy$3, dummy$4, dummy$5, \stage1_indices[1] [0]}),
     .A({1'b0, 1'b0, 1'b1, 1'b0}), .B({1'b0, 1'b0, 1'b1, 1'b1}), .S(
    \stage1[1].gt ));
  VDW_WMUX4_CIM_2 U$15(.Z({dummy$6, dummy$7, dummy$8, \stage1_indices[2] [0]}),
     .A({1'b0, 1'b1, 1'b0, 1'b0}), .B({1'b0, 1'b1, 1'b0, 1'b1}), .S(
    \stage1[2].gt ));
  VDW_WMUX4_CIM_1 U$16(.Z({dummy$9, dummy$10, dummy$11, \stage1_indices[3] [0]}),
     .A({1'b0, 1'b1, 1'b1, 1'b0}), .B({1'b0, 1'b1, 1'b1, 1'b1}), .S(
    \stage1[3].gt ));
  VDW_WMUX4_CIM U$17(.Z({dummy$12, dummy$13, dummy$14, \stage1_indices[4] [0]}),
     .A({1'b1, 1'b0, 1'b0, 1'b0}), .B({1'b1, 1'b0, 1'b0, 1'b1}), .S(
    \stage1[4].gt ));
  VDW_WMUX18 U$18(.Z({ final_winner[17:0] }), .A({ \stage3_winners[1] [17:0] }), .B({ \stage3_winners[0] [17:0] }), .S(gt_final));
  VDW_WMUX18 U$19(.Z({ \stage3_winners[0] [17:0] }), .A({ \stage2_winners[0] [17:0] }), .B({ \stage2_winners[1] [17:0] }), .S(\stage3[0].gt ));
  assign \stage3_winners[1] [17] = \stage2_winners[2] [17];
  assign \stage3_winners[1] [16] = \stage2_winners[2] [16];
  assign \stage3_winners[1] [15] = \stage2_winners[2] [15];
  assign \stage3_winners[1] [14] = \stage2_winners[2] [14];
  assign \stage3_winners[1] [13] = \stage2_winners[2] [13];
  assign \stage3_winners[1] [12] = \stage2_winners[2] [12];
  assign \stage3_winners[1] [11] = \stage2_winners[2] [11];
  assign \stage3_winners[1] [10] = \stage2_winners[2] [10];
  assign \stage3_winners[1] [9] = \stage2_winners[2] [9];
  assign \stage3_winners[1] [8] = \stage2_winners[2] [8];
  assign \stage3_winners[1] [7] = \stage2_winners[2] [7];
  assign \stage3_winners[1] [6] = \stage2_winners[2] [6];
  assign \stage3_winners[1] [5] = \stage2_winners[2] [5];
  assign \stage3_winners[1] [4] = \stage2_winners[2] [4];
  assign \stage3_winners[1] [3] = \stage2_winners[2] [3];
  assign \stage3_winners[1] [2] = \stage2_winners[2] [2];
  assign \stage3_winners[1] [1] = \stage2_winners[2] [1];
  assign \stage3_winners[1] [0] = \stage2_winners[2] [0];
  VDW_WMUX18 U$38(.Z({ \stage2_winners[0] [17:0] }), .A({ \stage1_winners[0] [17:0] }), .B({ \stage1_winners[1] [17:0] }), .S(\stage2[0].gt ));
  VDW_WMUX18 U$39(.Z({ \stage2_winners[1] [17:0] }), .A({ \stage1_winners[2] [17:0] }), .B({ \stage1_winners[3] [17:0] }), .S(\stage2[1].gt ));
  assign \stage2_winners[2] [17] = \stage1_winners[4] [17];
  assign \stage2_winners[2] [16] = \stage1_winners[4] [16];
  assign \stage2_winners[2] [15] = \stage1_winners[4] [15];
  assign \stage2_winners[2] [14] = \stage1_winners[4] [14];
  assign \stage2_winners[2] [13] = \stage1_winners[4] [13];
  assign \stage2_winners[2] [12] = \stage1_winners[4] [12];
  assign \stage2_winners[2] [11] = \stage1_winners[4] [11];
  assign \stage2_winners[2] [10] = \stage1_winners[4] [10];
  assign \stage2_winners[2] [9] = \stage1_winners[4] [9];
  assign \stage2_winners[2] [8] = \stage1_winners[4] [8];
  assign \stage2_winners[2] [7] = \stage1_winners[4] [7];
  assign \stage2_winners[2] [6] = \stage1_winners[4] [6];
  assign \stage2_winners[2] [5] = \stage1_winners[4] [5];
  assign \stage2_winners[2] [4] = \stage1_winners[4] [4];
  assign \stage2_winners[2] [3] = \stage1_winners[4] [3];
  assign \stage2_winners[2] [2] = \stage1_winners[4] [2];
  assign \stage2_winners[2] [1] = \stage1_winners[4] [1];
  assign \stage2_winners[2] [0] = \stage1_winners[4] [0];
  VDW_WMUX18 U$58(.Z({ \stage1_winners[0] [17:0] }), .A({ data_in[17:0] }), .B({ data_in[35:18] }), .S(\stage1[0].gt ));
  VDW_WMUX18 U$59(.Z({ \stage1_winners[1] [17:0] }), .A({ data_in[53:36] }), .B({ data_in[71:54] }), .S(\stage1[1].gt ));
  VDW_WMUX18 U$60(.Z({ \stage1_winners[2] [17:0] }), .A({ data_in[89:72] }), .B({ data_in[107:90] }), .S(\stage1[2].gt ));
  VDW_WMUX18 U$61(.Z({ \stage1_winners[3] [17:0] }), .A({ data_in[125:108] }), .B({ data_in[143:126] }), .S(\stage1[3].gt ));
  VDW_WMUX18 U$62(.Z({ \stage1_winners[4] [17:0] }), .A({ data_in[161:144] }), .B({ data_in[179:162] }), .S(\stage1[4].gt ));
  assign max_value[0] = final_winner[0];
  assign max_value[1] = final_winner[1];
  assign max_value[2] = final_winner[2];
  assign max_value[3] = final_winner[3];
  assign max_value[4] = final_winner[4];
  assign max_value[5] = final_winner[5];
  assign max_value[6] = final_winner[6];
  assign max_value[7] = final_winner[7];
  assign max_value[8] = final_winner[8];
  assign max_value[9] = final_winner[9];
  assign max_value[10] = final_winner[10];
  assign max_value[11] = final_winner[11];
  assign max_value[12] = final_winner[12];
  assign max_value[13] = final_winner[13];
  assign max_value[14] = final_winner[14];
  assign max_value[15] = final_winner[15];
  assign max_value[16] = final_winner[16];
  assign max_value[17] = final_winner[17];
  _HDFF_verplex \max_index_reg[3] (.Q(max_index[3]), .QN( ), .S(N$4), .R(n132)
    , .CK(clk), .D(final_index[3]));
  _HDFF_verplex \max_index_reg[2] (.Q(max_index[2]), .QN( ), .S(N$3), .R(n132)
    , .CK(clk), .D(final_index[2]));
  _HDFF_verplex \max_index_reg[1] (.Q(max_index[1]), .QN( ), .S(N$2), .R(n132)
    , .CK(clk), .D(final_index[1]));
  _HDFF_verplex \max_index_reg[0] (.Q(max_index[0]), .QN( ), .S(N$1), .R(n132)
    , .CK(clk), .D(final_index[0]));
  not U$81(n132, rst_n);
  compare_n_out cmp_final(.a({ \stage3_winners[0] [17:0] }), .b({ \stage3_winners[1] [17:0] }), .max(gt_final));
  compare_n_out \stage1[0].cmp (.a({ data_in[35:18] }), .b({ data_in[17:0] }), .max(\stage1[0].gt ));
  compare_n_out \stage1[1].cmp (.a({ data_in[71:54] }), .b({ data_in[53:36] }), .max(\stage1[1].gt ));
  compare_n_out \stage1[2].cmp (.a({ data_in[107:90] }), .b({ data_in[89:72] }), .max(\stage1[2].gt ));
  compare_n_out \stage1[3].cmp (.a({ data_in[143:126] }), .b({ data_in[125:108] }), .max(\stage1[3].gt ));
  compare_n_out \stage1[4].cmp (.a({ data_in[179:162] }), .b({ data_in[161:144] }), .max(\stage1[4].gt ));
  compare_n_out \stage2[0].cmp (.a({ \stage1_winners[1] [17:0] }), .b({ \stage1_winners[0] [17:0] }), .max(\stage2[0].gt ));
  compare_n_out \stage2[1].cmp (.a({ \stage1_winners[3] [17:0] }), .b({ \stage1_winners[2] [17:0] }), .max(\stage2[1].gt ));
  compare_n_out \stage3[0].cmp (.a({ \stage2_winners[1] [17:0] }), .b({ \stage2_winners[0] [17:0] }), .max(\stage3[0].gt ));
endmodule

module VDW_ONEHOT_SEL_2_1(Z, S, D1, D0);
// conformal library_module
input   [1:0] S;
input   [0:0] D1;
input   [0:0] D0;
output  [0:0] Z;
wire  N$1, N$2;
wire   [0:0] Z;
wire   [1:0] S;
wire   [0:0] D1;
wire   [0:0] D0;
  or U$1(Z[0], N$2, N$1);
  and U$2(N$1, D0[0], S[0]);
  and U$3(N$2, D1[0], S[1]);
endmodule

module decoder_4_to_10(in_val, out_activehigh);
input   [3:0] in_val;
output  [0:9] out_activehigh;
wire  n159_21, n159_20, n158_11, n157_10, n156_9, n155_8, n154_7, n153_6, n152_5, 
    n159_19, n159_18, n158_10, n157_9, n156_8, n155_7, n154_6, n153_5, n152_4, 
    n159_17, n159_16, n158_9, n157_8, n156_7, n155_6, n154_5, n153_4, n159_15, 
    n159_14, n158_8, n157_7, n156_6, n155_5, n154_4, n159_13, n159_12, n158_7, 
    n157_6, n156_5, n155_4, n159_11, n159_10, n158_6, n157_5, n156_4, n159_9, 
    n159_8, n158_5, n157_4, n159_7, n159_6, n158_4, n159_5, n159_4, n159_3, 
    n159_2, n159, n158_2, n158, n157_2, n157, n156_2, n156, n155_2, n155, 
    n154_2, n154, N$1, n153_2, n153, n152_2, n152, N$2, n150_2, n150, n151, 
    N$3;
wire   [0:9] out_activehigh;
wire   [3:0] in_val;
  VDW_ONEHOT_SEL_2_1 U$1(.Z({out_activehigh[0]}), .S({n159_21, n150}), .D1({1'b0}),
     .D0({1'b1}));
  or U$2(n159_21, n159_20, n159_2);
  or U$3(n159_20, n158_11, n159);
  or U$4(n158_11, n157_10, n158);
  or U$5(n157_10, n156_9, n157);
  or U$6(n156_9, n155_8, n156);
  or U$7(n155_8, n154_7, n155);
  or U$8(n154_7, n153_6, n154);
  or U$9(n153_6, n152_5, n153);
  or U$10(n152_5, n151, n152);
  VDW_ONEHOT_SEL_2_1 U$11(.Z({out_activehigh[1]}), .S({n151, n159_19}), .D1({
    1'b1}), .D0({1'b0}));
  or U$12(n159_19, n159_18, n159_2);
  or U$13(n159_18, n158_10, n159);
  or U$14(n158_10, n157_9, n158);
  or U$15(n157_9, n156_8, n157);
  or U$16(n156_8, n155_7, n156);
  or U$17(n155_7, n154_6, n155);
  or U$18(n154_6, n153_5, n154);
  or U$19(n153_5, n152_4, n153);
  or U$20(n152_4, n150, n152);
  VDW_ONEHOT_SEL_2_1 U$21(.Z({out_activehigh[2]}), .S({n159_17, n152}), .D1({
    1'b0}), .D0({1'b1}));
  or U$22(n159_17, n159_16, n159_2);
  or U$23(n159_16, n158_9, n159);
  or U$24(n158_9, n157_8, n158);
  or U$25(n157_8, n156_7, n157);
  or U$26(n156_7, n155_6, n156);
  or U$27(n155_6, n154_5, n155);
  or U$28(n154_5, n153_4, n154);
  or U$29(n153_4, n150_2, n153);
  VDW_ONEHOT_SEL_2_1 U$30(.Z({out_activehigh[3]}), .S({n159_15, n153}), .D1({
    1'b0}), .D0({1'b1}));
  or U$31(n159_15, n159_14, n159_2);
  or U$32(n159_14, n158_8, n159);
  or U$33(n158_8, n157_7, n158);
  or U$34(n157_7, n156_6, n157);
  or U$35(n156_6, n155_5, n156);
  or U$36(n155_5, n154_4, n155);
  or U$37(n154_4, n152_2, n154);
  VDW_ONEHOT_SEL_2_1 U$38(.Z({out_activehigh[4]}), .S({n159_13, n154}), .D1({
    1'b0}), .D0({1'b1}));
  or U$39(n159_13, n159_12, n159_2);
  or U$40(n159_12, n158_7, n159);
  or U$41(n158_7, n157_6, n158);
  or U$42(n157_6, n156_5, n157);
  or U$43(n156_5, n155_4, n156);
  or U$44(n155_4, n153_2, n155);
  VDW_ONEHOT_SEL_2_1 U$45(.Z({out_activehigh[5]}), .S({n159_11, n155}), .D1({
    1'b0}), .D0({1'b1}));
  or U$46(n159_11, n159_10, n159_2);
  or U$47(n159_10, n158_6, n159);
  or U$48(n158_6, n157_5, n158);
  or U$49(n157_5, n156_4, n157);
  or U$50(n156_4, n154_2, n156);
  VDW_ONEHOT_SEL_2_1 U$51(.Z({out_activehigh[6]}), .S({n159_9, n156}), .D1({1'b0}),
     .D0({1'b1}));
  or U$52(n159_9, n159_8, n159_2);
  or U$53(n159_8, n158_5, n159);
  or U$54(n158_5, n157_4, n158);
  or U$55(n157_4, n155_2, n157);
  VDW_ONEHOT_SEL_2_1 U$56(.Z({out_activehigh[7]}), .S({n159_7, n157}), .D1({1'b0}),
     .D0({1'b1}));
  or U$57(n159_7, n159_6, n159_2);
  or U$58(n159_6, n158_4, n159);
  or U$59(n158_4, n156_2, n158);
  VDW_ONEHOT_SEL_2_1 U$60(.Z({out_activehigh[8]}), .S({n159_5, n158}), .D1({1'b0}),
     .D0({1'b1}));
  or U$61(n159_5, n159_4, n159_2);
  or U$62(n159_4, n157_2, n159);
  VDW_ONEHOT_SEL_2_1 U$63(.Z({out_activehigh[9]}), .S({n159_3, n159}), .D1({1'b0}),
     .D0({1'b1}));
  or U$64(n159_3, n158_2, n159_2);
  nor U$65(n159_2, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159);
  nor U$66(n159, N$3, in_val[1], in_val[2], N$1);
  or U$67(n158_2, n157_2, n158);
  nor U$68(n158, in_val[0], in_val[1], in_val[2], N$1);
  or U$69(n157_2, n156_2, n157);
  and U$70(n157, in_val[0], in_val[1], in_val[2], N$1);
  or U$71(n156_2, n155_2, n156);
  and U$72(n156, N$3, in_val[1], in_val[2], N$1);
  or U$73(n155_2, n154_2, n155);
  and U$74(n155, in_val[0], N$2, in_val[2], N$1);
  or U$75(n154_2, n153_2, n154);
  not U$76(N$1, in_val[3]);
  and U$77(n154, N$3, N$2, in_val[2], N$1);
  or U$78(n153_2, n152_2, n153);
  nor U$79(n153, N$3, N$2, in_val[2], in_val[3]);
  or U$80(n152_2, n150_2, n152);
  not U$81(N$2, in_val[1]);
  nor U$82(n152, in_val[0], N$2, in_val[2], in_val[3]);
  or U$83(n150_2, n151, n150);
  nor U$84(n150, in_val[0], in_val[1], in_val[2], in_val[3]);
  not U$85(N$3, in_val[0]);
  nor U$86(n151, N$3, in_val[1], in_val[2], in_val[3]);
endmodule

module mytop(in, clk, rst_n, updown, out_activehigh, done);
input  clk, rst_n, updown;
output done;
input   [127:0] in;
output  [0:9] out_activehigh;
wire  n5893_2, n5900_2, n5900, n5893, done, updown, rst_n, clk;
wire  N$1, N$2, N$3;
wire   [1:0] n5900_3;
wire   [1:0] n5902;
wire   [17:0] max;
wire   [3:0] out;
wire   [179:0] layer2_out;
wire   [1:0] counter;
wire   [179:0] layer1_out;
wire   [0:9] out_activehigh;
wire   [127:0] in;
  assign N$1 = 1'b0;
  assign N$2 = 1'b0;
  assign N$3 = 1'b0;
  _HDFF_verplex \counter_reg[1] (.Q(counter[1]), .QN( ), .S(N$2), .R(n5893_2)
    , .CK(clk), .D(n5900_3[1]));
  _HDFF_verplex \counter_reg[0] (.Q(counter[0]), .QN( ), .S(N$1), .R(n5893_2)
    , .CK(clk), .D(n5900_3[0]));
  VDW_WMUX2 U$1(.Z({ n5900_3[1:0] }), .A({ counter[1:0] }), .B({ n5902[1:0] }), .S(n5900));
  VDW_ADD_2_1_0_CIM add_5902_28(.SUM({ n5902[1:0] }), .A({ counter[1:0] }), .B({1'b0, 1'b1}));
  not U$2(n5893_2, updown);
  _HDFF_verplex done_reg(.Q(done), .QN( ), .S(N$3), .R(n5893), .CK(clk), .D(
    n5900_2));
  _HMUX U$3(.O(n5900_2), .I0(1'b1), .I1(done), .S(n5900));
  VDW_LT_u2_CIM lt_5900_17(.Z(n5900), .A({ counter[1:0] }), .B({1'b1, 1'b1}));
  not U$4(n5893, updown);
  layer1 instanceL1(.clk(clk), .rst_n(rst_n), .updown(updown), .in({ in[127:0] }), .out({ layer1_out[179:0] }));
  layer2 instanceL2(.clk(clk), .rst_n(rst_n), .in({ layer1_out[179:0] }), .out({ layer2_out[179:0] }));
  find_max_index uut(.data_in({ layer2_out[179:0] }), .clk(clk), .rst_n(rst_n), .max_index({ out[3:0] }),
     .max_value({ max[17:0] }));
  decoder_4_to_10 dut(.in_val({ out[3:0] }), .out_activehigh({ out_activehigh[0:9] }));
endmodule

module _HMUX(O, I0, I1, S);
// verplex MUX
output  O;
input   I0, I1, S;
  not  (N1, S);
  and  (N2, S, I1);
  and  (N3, N1, I0);
  or   (O, N2, N3);
endmodule

module _HDFF_verplex(Q, QN, S, R, CK, D);
// verplex DFF
output  Q, QN;
input   S, R, CK, D;
wire   N1;
  DFF_UDP  i0(N1, S, R, CK, D);
  buf  (Q, N1);
  not  (QN, N1);
endmodule

primitive DFF_UDP(Q, S, R, CK, D);
output Q;
input  S, R, CK, D;
reg    Q;
  table
    1  0   ?    ?  :  ?  :  1; // Asserting preset
    *  0   ?    ?  :  1  :  1; // Changing preset
    ?  1   ?    ?  :  ?  :  0; // Asserting reset (dominates preset)
    0  *   ?    ?  :  0  :  0; // Changing reset
    0  ?   (01) 0  :  ?  :  0; // rising clock
    ?  0   (01) 1  :  ?  :  1; // rising clock 
    0  ?   p    0  :  0  :  0; // potential rising clock
    ?  0   p    1  :  1  :  1; // potential rising clock
    0  0   n    ?  :  ?  :  -; // Clock falling register output does not change
    0  0   ?    *  :  ?  :  -; // Changing Data
  endtable
endprimitive

