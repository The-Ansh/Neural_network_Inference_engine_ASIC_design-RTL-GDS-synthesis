`timescale 1ns / 1ns

module adder_5to6 (
    input  signed [4:0] a,
    input  signed [4:0] b,
    output signed [5:0] sum
);
    assign sum = a + b;
endmodule

module adder_6to7 (
    input signed [5:0] a,
    input signed [5:0] b,
    output signed [6:0] sum
);
    assign sum = a + b;
endmodule

module adder_7to8 (
    input signed [6:0] a,
    input signed [6:0] b,
    output signed [7:0] sum
);
    assign sum = a + b;
endmodule

module adder_8to9 (
    input  signed [7:0] a,
    input  signed [7:0] b,
    output signed [8:0] sum
);
    assign sum = a + b;
endmodule

module adder_9to10 (
    input signed [8:0] a,
    input signed [8:0] b,
    output signed [9:0] sum
);
    assign sum = a + b;
endmodule

module adder_10to10 (
    input signed [9:0] a,
    input signed [9:0] b,
    output signed [9:0] sum
);
    wire signed [10:0] result;
    assign result = a + b;
    assign sum = result[9:0];
endmodule

module compare_n_out(
    input  [17:0] a,
    input  [17:0] b,
    output wire  max // 1 if a > b, else 0 (explicitly declared as wire)
);
    // The result of a comparison is already a 1-bit value (1 for true, 0 for false).
    assign max = (a > b);
endmodule

module find_max_index #(
    parameter NUM_INPUTS = 10,
    parameter DATA_WIDTH = 18
)(
    input [179:0] data_in,
    input clk,
    input rst_n,
    output reg [3:0] max_index,
    output wire [17:0] max_value
);
    // Intermediate signals for each stage of the comparator tree
    wire [17:0] stage1_winners [0:4];
    wire [17:0] stage2_winners [0:2];
    wire [17:0] stage3_winners [0:1];
    wire [17:0] final_winner;

    wire [3:0] stage1_indices [0:4];
    wire [3:0] stage2_indices [0:2];
    wire [3:0] stage3_indices [0:1];
    wire [3:0] final_index;

    genvar i;
    generate
        for (i = 0; i < 5; i = i + 1) begin : stage1
            wire gt;
            compare_n_out cmp (
                .a(data_in[(2*i+2)*DATA_WIDTH - 1 : (2*i+1)*DATA_WIDTH]),
                .b(data_in[(2*i+1)*DATA_WIDTH - 1 : (2*i)*DATA_WIDTH]),
                .max(gt)
            );
            assign stage1_winners[i] = gt ? data_in[(2*i+2)*DATA_WIDTH - 1 : (2*i+1)*DATA_WIDTH] : data_in[(2*i+1)*DATA_WIDTH - 1 : (2*i)*DATA_WIDTH];
            assign stage1_indices[i] = gt ? (2*i+1) : (2*i);
        end

        for (i = 0; i < 2; i = i + 1) begin : stage2
            wire gt;
            compare_n_out cmp (
                .a(stage1_winners[2*i+1]),
                .b(stage1_winners[2*i]),
                .max(gt)
            );
            assign stage2_winners[i] = gt ? stage1_winners[2*i+1] : stage1_winners[2*i];
            assign stage2_indices[i] = gt ? stage1_indices[2*i+1] : stage1_indices[2*i];
        end
        assign stage2_winners[2] = stage1_winners[4]; // Carry forward the unpaired winner
        assign stage2_indices[2] = stage1_indices[4];

        for (i = 0; i < 1; i = i + 1) begin : stage3
            wire gt;
            compare_n_out cmp (
                .a(stage2_winners[2*i+1]),
                .b(stage2_winners[2*i]),
                .max(gt)
            );
            assign stage3_winners [i] = gt ? stage2_winners[2*i+1] : stage2_winners[2*i];
            assign stage3_indices[i] = gt ? stage2_indices[2*i+1] : stage2_indices[2*i];
        end
        assign stage3_winners [1] = stage2_winners[2]; // Carry forward the unpaired winner
        assign stage3_indices[1] = stage2_indices[2];
        
        wire gt_final;
        compare_n_out cmp_final (
            .a(stage3_winners[0]),
            .b(stage3_winners[1]),
            .max(gt_final)
        );
        assign final_winner = gt_final ? stage3_winners[0] : stage3_winners[1];
        assign final_index = gt_final ? stage3_indices[0] : stage3_indices[1];
    endgenerate

    assign max_value = final_winner;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            max_index <= 4'b0000;
        else
        max_index <= final_index;
    end
endmodule

module decoder_4_to_10 (
    input  wire [3:0]  in_val,
    output reg  [0:9]  out_activehigh
);

    // This combinational block updates whenever 'in_val' changes.
    always @(*) begin
        // Default to all zeros to avoid latches for unspecified cases
        out_activehigh = 10'b0; 

        case (in_val)
            4'd0: out_activehigh[0] = 1'b1;
            4'd1: out_activehigh[1] = 1'b1;
            4'd2: out_activehigh[2] = 1'b1;
            4'd3: out_activehigh[3] = 1'b1; 
            4'd4: out_activehigh[4] = 1'b1;
            4'd5: out_activehigh[5] = 1'b1;
            4'd6: out_activehigh[6] = 1'b1;
            4'd7: out_activehigh[7] = 1'b1;
            4'd8: out_activehigh[8] = 1'b1;
            4'd9: out_activehigh[9] = 1'b1;
            // A default case is good practice, though not strictly
            // necessary here since we defaulted to zero above.
            default: out_activehigh = 10'b0; 
        endcase
    end

endmodule

module multiplier9514(
    output wire signed [13:0] prod,   // signed output (14 bits)
    input  wire        [8:0] num1,   // unsigned 9-bit input (multiplicand)
    input  wire signed [4:0] num2    // signed 5-bit input (multiplier)
);
    wire [8:0] partial_prods [0:4];
    wire signed [13:0] shifted_pps [0:4];
    wire signed [13:0] intermediate_sums [0:2];
    genvar i;
    generate
        for (i = 0; i < 5; i = i + 1) begin : partial_product_generation
            assign partial_prods[i] = num2[i] ? num1 : 9'b0;
            assign shifted_pps[i] = partial_prods[i] << i;
        end
    endgenerate
    assign intermediate_sums[0] = shifted_pps[0] + shifted_pps[1];
    assign intermediate_sums[1] = intermediate_sums[0] + shifted_pps[2];
    assign intermediate_sums[2] = intermediate_sums[1] + shifted_pps[3];
    assign prod = intermediate_sums[2] - shifted_pps[4];
endmodule

module ReLU_10bit (
    input  wire [9:0] in_data,
    output wire [8:0] out_data
);

    // If the sign bit (in_data[9]) is 0, pass the data through.
    // Otherwise, output 0.
    assign out_data = (in_data[9] == 1'b0) ? in_data[8:0] : 9'd0;

endmodule

module ReLU_19bit(
    //input  wire        clk,
    //input  wire        rst_n,
    input  wire [18:0] in_data,
    output wire  [17:0] out_data
);

    assign out_data = (in_data[18] == 1'b0) ? in_data[17:0] : 18'd0;

    // always @(posedge clk or negedge rst_n) begin
    //     if (!rst_n) begin
    //         out_data <= 18'd0;
    //     end

    //     else begin
    //         if (in_data[18] == 1'b0) begin
    //             // Positive input, pass through
    //             out_data <= in_data[17:0];
    //         end else begin
    //             // Negative input, output zero
    //             out_data <= 18'd0;
    //         end
    //     end
    // end
endmodule

module layer1 #(
    parameter ROWS      = 20,
    parameter COLS      = 256,
    parameter A_WIDTH   = 5
)(
    input clk,
    input rst_n,
    input updown,
    // Input vector 'B' (256x1, 1-bit elements) flattened to a single vector
    input [0:127] in, 
    output [179:0] out
);

    // reg [4:0] A [0:19][0:255];
    // initial begin
    //     $readmemb("w1.mem", A);
    // end
    reg [0:255] B;

wire [4:0] A [0:19][0:255];
assign A[0][0] = 5'b00001;
assign A[0][1] = 5'b00001;
assign A[0][2] = 5'b00000;
assign A[0][3] = 5'b11110;
assign A[0][4] = 5'b00001;
assign A[0][5] = 5'b00001;
assign A[0][6] = 5'b00100;
assign A[0][7] = 5'b11111;
assign A[0][8] = 5'b11111;
assign A[0][9] = 5'b11101;
assign A[0][10] = 5'b00000;
assign A[0][11] = 5'b11110;
assign A[0][12] = 5'b11110;
assign A[0][13] = 5'b00001;
assign A[0][14] = 5'b00001;
assign A[0][15] = 5'b00000;
assign A[0][16] = 5'b11111;
assign A[0][17] = 5'b11110;
assign A[0][18] = 5'b11111;
assign A[0][19] = 5'b00011;
assign A[0][20] = 5'b00000;
assign A[0][21] = 5'b11111;
assign A[0][22] = 5'b00001;
assign A[0][23] = 5'b11111;
assign A[0][24] = 5'b00000;
assign A[0][25] = 5'b00000;
assign A[0][26] = 5'b11110;
assign A[0][27] = 5'b00001;
assign A[0][28] = 5'b11111;
assign A[0][29] = 5'b00001;
assign A[0][30] = 5'b00000;
assign A[0][31] = 5'b00001;
assign A[0][32] = 5'b11111;
assign A[0][33] = 5'b00011;
assign A[0][34] = 5'b11110;
assign A[0][35] = 5'b00010;
assign A[0][36] = 5'b00000;
assign A[0][37] = 5'b11111;
assign A[0][38] = 5'b00000;
assign A[0][39] = 5'b00001;
assign A[0][40] = 5'b00000;
assign A[0][41] = 5'b11111;
assign A[0][42] = 5'b00010;
assign A[0][43] = 5'b11110;
assign A[0][44] = 5'b00000;
assign A[0][45] = 5'b00000;
assign A[0][46] = 5'b00010;
assign A[0][47] = 5'b00010;
assign A[0][48] = 5'b11111;
assign A[0][49] = 5'b11101;
assign A[0][50] = 5'b00000;
assign A[0][51] = 5'b00000;
assign A[0][52] = 5'b00000;
assign A[0][53] = 5'b00000;
assign A[0][54] = 5'b00000;
assign A[0][55] = 5'b00000;
assign A[0][56] = 5'b00001;
assign A[0][57] = 5'b11111;
assign A[0][58] = 5'b11111;
assign A[0][59] = 5'b00001;
assign A[0][60] = 5'b00010;
assign A[0][61] = 5'b00010;
assign A[0][62] = 5'b00000;
assign A[0][63] = 5'b00010;
assign A[0][64] = 5'b00000;
assign A[0][65] = 5'b11111;
assign A[0][66] = 5'b11111;
assign A[0][67] = 5'b11111;
assign A[0][68] = 5'b00001;
assign A[0][69] = 5'b00000;
assign A[0][70] = 5'b11110;
assign A[0][71] = 5'b00010;
assign A[0][72] = 5'b00001;
assign A[0][73] = 5'b00000;
assign A[0][74] = 5'b11111;
assign A[0][75] = 5'b11101;
assign A[0][76] = 5'b00001;
assign A[0][77] = 5'b11110;
assign A[0][78] = 5'b00000;
assign A[0][79] = 5'b00000;
assign A[0][80] = 5'b11101;
assign A[0][81] = 5'b11111;
assign A[0][82] = 5'b00001;
assign A[0][83] = 5'b00010;
assign A[0][84] = 5'b11110;
assign A[0][85] = 5'b11111;
assign A[0][86] = 5'b11111;
assign A[0][87] = 5'b00000;
assign A[0][88] = 5'b00010;
assign A[0][89] = 5'b11110;
assign A[0][90] = 5'b11111;
assign A[0][91] = 5'b00000;
assign A[0][92] = 5'b00001;
assign A[0][93] = 5'b00001;
assign A[0][94] = 5'b11110;
assign A[0][95] = 5'b00010;
assign A[0][96] = 5'b11111;
assign A[0][97] = 5'b11111;
assign A[0][98] = 5'b11111;
assign A[0][99] = 5'b00000;
assign A[0][100] = 5'b00001;
assign A[0][101] = 5'b11111;
assign A[0][102] = 5'b00001;
assign A[0][103] = 5'b00010;
assign A[0][104] = 5'b11101;
assign A[0][105] = 5'b11111;
assign A[0][106] = 5'b11101;
assign A[0][107] = 5'b00000;
assign A[0][108] = 5'b11110;
assign A[0][109] = 5'b00000;
assign A[0][110] = 5'b00000;
assign A[0][111] = 5'b00001;
assign A[0][112] = 5'b11111;
assign A[0][113] = 5'b00000;
assign A[0][114] = 5'b00010;
assign A[0][115] = 5'b11110;
assign A[0][116] = 5'b00000;
assign A[0][117] = 5'b11110;
assign A[0][118] = 5'b11110;
assign A[0][119] = 5'b11101;
assign A[0][120] = 5'b00001;
assign A[0][121] = 5'b11111;
assign A[0][122] = 5'b11111;
assign A[0][123] = 5'b11111;
assign A[0][124] = 5'b00000;
assign A[0][125] = 5'b11111;
assign A[0][126] = 5'b11111;
assign A[0][127] = 5'b00000;
assign A[0][128] = 5'b00001;
assign A[0][129] = 5'b00000;
assign A[0][130] = 5'b00001;
assign A[0][131] = 5'b00000;
assign A[0][132] = 5'b00001;
assign A[0][133] = 5'b00000;
assign A[0][134] = 5'b11111;
assign A[0][135] = 5'b00000;
assign A[0][136] = 5'b00001;
assign A[0][137] = 5'b11100;
assign A[0][138] = 5'b00010;
assign A[0][139] = 5'b00001;
assign A[0][140] = 5'b00000;
assign A[0][141] = 5'b11111;
assign A[0][142] = 5'b11111;
assign A[0][143] = 5'b00000;
assign A[0][144] = 5'b00001;
assign A[0][145] = 5'b11110;
assign A[0][146] = 5'b00011;
assign A[0][147] = 5'b00000;
assign A[0][148] = 5'b00000;
assign A[0][149] = 5'b11110;
assign A[0][150] = 5'b00001;
assign A[0][151] = 5'b11110;
assign A[0][152] = 5'b00000;
assign A[0][153] = 5'b00001;
assign A[0][154] = 5'b11101;
assign A[0][155] = 5'b11111;
assign A[0][156] = 5'b11111;
assign A[0][157] = 5'b11111;
assign A[0][158] = 5'b11111;
assign A[0][159] = 5'b00010;
assign A[0][160] = 5'b00000;
assign A[0][161] = 5'b00000;
assign A[0][162] = 5'b11110;
assign A[0][163] = 5'b00000;
assign A[0][164] = 5'b11110;
assign A[0][165] = 5'b11111;
assign A[0][166] = 5'b00001;
assign A[0][167] = 5'b11101;
assign A[0][168] = 5'b00000;
assign A[0][169] = 5'b11111;
assign A[0][170] = 5'b11111;
assign A[0][171] = 5'b00001;
assign A[0][172] = 5'b11111;
assign A[0][173] = 5'b00000;
assign A[0][174] = 5'b00001;
assign A[0][175] = 5'b11111;
assign A[0][176] = 5'b11111;
assign A[0][177] = 5'b11101;
assign A[0][178] = 5'b00000;
assign A[0][179] = 5'b00001;
assign A[0][180] = 5'b00000;
assign A[0][181] = 5'b00000;
assign A[0][182] = 5'b00000;
assign A[0][183] = 5'b00001;
assign A[0][184] = 5'b11111;
assign A[0][185] = 5'b11110;
assign A[0][186] = 5'b11110;
assign A[0][187] = 5'b00001;
assign A[0][188] = 5'b00000;
assign A[0][189] = 5'b00001;
assign A[0][190] = 5'b11111;
assign A[0][191] = 5'b00010;
assign A[0][192] = 5'b00000;
assign A[0][193] = 5'b11110;
assign A[0][194] = 5'b11110;
assign A[0][195] = 5'b11111;
assign A[0][196] = 5'b00001;
assign A[0][197] = 5'b11100;
assign A[0][198] = 5'b00000;
assign A[0][199] = 5'b11111;
assign A[0][200] = 5'b00010;
assign A[0][201] = 5'b00001;
assign A[0][202] = 5'b00001;
assign A[0][203] = 5'b00001;
assign A[0][204] = 5'b00001;
assign A[0][205] = 5'b11110;
assign A[0][206] = 5'b00000;
assign A[0][207] = 5'b00000;
assign A[0][208] = 5'b11111;
assign A[0][209] = 5'b11110;
assign A[0][210] = 5'b11111;
assign A[0][211] = 5'b11111;
assign A[0][212] = 5'b00001;
assign A[0][213] = 5'b11110;
assign A[0][214] = 5'b00000;
assign A[0][215] = 5'b00000;
assign A[0][216] = 5'b00011;
assign A[0][217] = 5'b00000;
assign A[0][218] = 5'b00000;
assign A[0][219] = 5'b00001;
assign A[0][220] = 5'b11111;
assign A[0][221] = 5'b00000;
assign A[0][222] = 5'b00001;
assign A[0][223] = 5'b00000;
assign A[0][224] = 5'b00011;
assign A[0][225] = 5'b00000;
assign A[0][226] = 5'b11111;
assign A[0][227] = 5'b00001;
assign A[0][228] = 5'b00001;
assign A[0][229] = 5'b00000;
assign A[0][230] = 5'b11101;
assign A[0][231] = 5'b00000;
assign A[0][232] = 5'b11110;
assign A[0][233] = 5'b00001;
assign A[0][234] = 5'b11110;
assign A[0][235] = 5'b00001;
assign A[0][236] = 5'b00000;
assign A[0][237] = 5'b00010;
assign A[0][238] = 5'b00001;
assign A[0][239] = 5'b00010;
assign A[0][240] = 5'b00000;
assign A[0][241] = 5'b11111;
assign A[0][242] = 5'b11111;
assign A[0][243] = 5'b11111;
assign A[0][244] = 5'b00010;
assign A[0][245] = 5'b00001;
assign A[0][246] = 5'b00010;
assign A[0][247] = 5'b00001;
assign A[0][248] = 5'b00011;
assign A[0][249] = 5'b00000;
assign A[0][250] = 5'b11111;
assign A[0][251] = 5'b00000;
assign A[0][252] = 5'b11110;
assign A[0][253] = 5'b00001;
assign A[0][254] = 5'b11110;
assign A[0][255] = 5'b11111;
assign A[1][0] = 5'b00010;
assign A[1][1] = 5'b11110;
assign A[1][2] = 5'b11111;
assign A[1][3] = 5'b00000;
assign A[1][4] = 5'b00000;
assign A[1][5] = 5'b11110;
assign A[1][6] = 5'b00001;
assign A[1][7] = 5'b11111;
assign A[1][8] = 5'b11111;
assign A[1][9] = 5'b00000;
assign A[1][10] = 5'b11110;
assign A[1][11] = 5'b00010;
assign A[1][12] = 5'b00001;
assign A[1][13] = 5'b11101;
assign A[1][14] = 5'b00001;
assign A[1][15] = 5'b00000;
assign A[1][16] = 5'b11111;
assign A[1][17] = 5'b11111;
assign A[1][18] = 5'b00000;
assign A[1][19] = 5'b00010;
assign A[1][20] = 5'b00000;
assign A[1][21] = 5'b11111;
assign A[1][22] = 5'b00000;
assign A[1][23] = 5'b00010;
assign A[1][24] = 5'b11111;
assign A[1][25] = 5'b00000;
assign A[1][26] = 5'b11101;
assign A[1][27] = 5'b00000;
assign A[1][28] = 5'b11111;
assign A[1][29] = 5'b11111;
assign A[1][30] = 5'b00010;
assign A[1][31] = 5'b00000;
assign A[1][32] = 5'b11110;
assign A[1][33] = 5'b11101;
assign A[1][34] = 5'b00000;
assign A[1][35] = 5'b00000;
assign A[1][36] = 5'b00000;
assign A[1][37] = 5'b00000;
assign A[1][38] = 5'b00000;
assign A[1][39] = 5'b11111;
assign A[1][40] = 5'b11110;
assign A[1][41] = 5'b11111;
assign A[1][42] = 5'b00000;
assign A[1][43] = 5'b00000;
assign A[1][44] = 5'b11111;
assign A[1][45] = 5'b11111;
assign A[1][46] = 5'b00000;
assign A[1][47] = 5'b00000;
assign A[1][48] = 5'b11111;
assign A[1][49] = 5'b00011;
assign A[1][50] = 5'b11111;
assign A[1][51] = 5'b11111;
assign A[1][52] = 5'b11101;
assign A[1][53] = 5'b00000;
assign A[1][54] = 5'b00001;
assign A[1][55] = 5'b11111;
assign A[1][56] = 5'b11110;
assign A[1][57] = 5'b00000;
assign A[1][58] = 5'b11111;
assign A[1][59] = 5'b11110;
assign A[1][60] = 5'b11111;
assign A[1][61] = 5'b00001;
assign A[1][62] = 5'b11101;
assign A[1][63] = 5'b00000;
assign A[1][64] = 5'b00000;
assign A[1][65] = 5'b00001;
assign A[1][66] = 5'b11110;
assign A[1][67] = 5'b11110;
assign A[1][68] = 5'b11101;
assign A[1][69] = 5'b00010;
assign A[1][70] = 5'b00001;
assign A[1][71] = 5'b11110;
assign A[1][72] = 5'b00000;
assign A[1][73] = 5'b11111;
assign A[1][74] = 5'b11110;
assign A[1][75] = 5'b00001;
assign A[1][76] = 5'b11110;
assign A[1][77] = 5'b11111;
assign A[1][78] = 5'b11111;
assign A[1][79] = 5'b11101;
assign A[1][80] = 5'b00000;
assign A[1][81] = 5'b11101;
assign A[1][82] = 5'b00001;
assign A[1][83] = 5'b11110;
assign A[1][84] = 5'b11110;
assign A[1][85] = 5'b00001;
assign A[1][86] = 5'b00000;
assign A[1][87] = 5'b00000;
assign A[1][88] = 5'b11111;
assign A[1][89] = 5'b11110;
assign A[1][90] = 5'b00001;
assign A[1][91] = 5'b00001;
assign A[1][92] = 5'b00000;
assign A[1][93] = 5'b00001;
assign A[1][94] = 5'b11111;
assign A[1][95] = 5'b00010;
assign A[1][96] = 5'b11111;
assign A[1][97] = 5'b00000;
assign A[1][98] = 5'b00000;
assign A[1][99] = 5'b00001;
assign A[1][100] = 5'b00010;
assign A[1][101] = 5'b00000;
assign A[1][102] = 5'b00010;
assign A[1][103] = 5'b00010;
assign A[1][104] = 5'b00011;
assign A[1][105] = 5'b11110;
assign A[1][106] = 5'b00001;
assign A[1][107] = 5'b11110;
assign A[1][108] = 5'b00001;
assign A[1][109] = 5'b11111;
assign A[1][110] = 5'b11111;
assign A[1][111] = 5'b11111;
assign A[1][112] = 5'b11111;
assign A[1][113] = 5'b11111;
assign A[1][114] = 5'b11110;
assign A[1][115] = 5'b11111;
assign A[1][116] = 5'b00000;
assign A[1][117] = 5'b00000;
assign A[1][118] = 5'b00001;
assign A[1][119] = 5'b00001;
assign A[1][120] = 5'b00000;
assign A[1][121] = 5'b00000;
assign A[1][122] = 5'b00001;
assign A[1][123] = 5'b11110;
assign A[1][124] = 5'b00000;
assign A[1][125] = 5'b00000;
assign A[1][126] = 5'b00000;
assign A[1][127] = 5'b00000;
assign A[1][128] = 5'b00000;
assign A[1][129] = 5'b00000;
assign A[1][130] = 5'b00001;
assign A[1][131] = 5'b00001;
assign A[1][132] = 5'b11110;
assign A[1][133] = 5'b00001;
assign A[1][134] = 5'b11111;
assign A[1][135] = 5'b11111;
assign A[1][136] = 5'b00000;
assign A[1][137] = 5'b11111;
assign A[1][138] = 5'b00001;
assign A[1][139] = 5'b00000;
assign A[1][140] = 5'b00000;
assign A[1][141] = 5'b00010;
assign A[1][142] = 5'b00000;
assign A[1][143] = 5'b00011;
assign A[1][144] = 5'b00000;
assign A[1][145] = 5'b00010;
assign A[1][146] = 5'b00011;
assign A[1][147] = 5'b11101;
assign A[1][148] = 5'b11101;
assign A[1][149] = 5'b11111;
assign A[1][150] = 5'b00000;
assign A[1][151] = 5'b00011;
assign A[1][152] = 5'b00001;
assign A[1][153] = 5'b00000;
assign A[1][154] = 5'b00010;
assign A[1][155] = 5'b11110;
assign A[1][156] = 5'b11111;
assign A[1][157] = 5'b00001;
assign A[1][158] = 5'b00001;
assign A[1][159] = 5'b00000;
assign A[1][160] = 5'b00010;
assign A[1][161] = 5'b11111;
assign A[1][162] = 5'b11111;
assign A[1][163] = 5'b00000;
assign A[1][164] = 5'b11111;
assign A[1][165] = 5'b00000;
assign A[1][166] = 5'b00010;
assign A[1][167] = 5'b11110;
assign A[1][168] = 5'b00000;
assign A[1][169] = 5'b11110;
assign A[1][170] = 5'b00001;
assign A[1][171] = 5'b11110;
assign A[1][172] = 5'b00000;
assign A[1][173] = 5'b00001;
assign A[1][174] = 5'b00011;
assign A[1][175] = 5'b00000;
assign A[1][176] = 5'b00001;
assign A[1][177] = 5'b11111;
assign A[1][178] = 5'b11111;
assign A[1][179] = 5'b11111;
assign A[1][180] = 5'b00000;
assign A[1][181] = 5'b00000;
assign A[1][182] = 5'b11110;
assign A[1][183] = 5'b00010;
assign A[1][184] = 5'b11111;
assign A[1][185] = 5'b11111;
assign A[1][186] = 5'b11101;
assign A[1][187] = 5'b00011;
assign A[1][188] = 5'b00010;
assign A[1][189] = 5'b11101;
assign A[1][190] = 5'b00011;
assign A[1][191] = 5'b00010;
assign A[1][192] = 5'b00011;
assign A[1][193] = 5'b11111;
assign A[1][194] = 5'b11111;
assign A[1][195] = 5'b00011;
assign A[1][196] = 5'b00011;
assign A[1][197] = 5'b11101;
assign A[1][198] = 5'b00001;
assign A[1][199] = 5'b11111;
assign A[1][200] = 5'b00001;
assign A[1][201] = 5'b00000;
assign A[1][202] = 5'b00001;
assign A[1][203] = 5'b00000;
assign A[1][204] = 5'b11111;
assign A[1][205] = 5'b00000;
assign A[1][206] = 5'b00000;
assign A[1][207] = 5'b11111;
assign A[1][208] = 5'b11111;
assign A[1][209] = 5'b11111;
assign A[1][210] = 5'b11111;
assign A[1][211] = 5'b11111;
assign A[1][212] = 5'b00001;
assign A[1][213] = 5'b00000;
assign A[1][214] = 5'b11110;
assign A[1][215] = 5'b00000;
assign A[1][216] = 5'b11111;
assign A[1][217] = 5'b11110;
assign A[1][218] = 5'b00001;
assign A[1][219] = 5'b11111;
assign A[1][220] = 5'b11111;
assign A[1][221] = 5'b00001;
assign A[1][222] = 5'b00000;
assign A[1][223] = 5'b00001;
assign A[1][224] = 5'b11101;
assign A[1][225] = 5'b11110;
assign A[1][226] = 5'b00000;
assign A[1][227] = 5'b11111;
assign A[1][228] = 5'b00100;
assign A[1][229] = 5'b00000;
assign A[1][230] = 5'b00001;
assign A[1][231] = 5'b11110;
assign A[1][232] = 5'b00010;
assign A[1][233] = 5'b00010;
assign A[1][234] = 5'b00001;
assign A[1][235] = 5'b00000;
assign A[1][236] = 5'b00001;
assign A[1][237] = 5'b11111;
assign A[1][238] = 5'b00011;
assign A[1][239] = 5'b11110;
assign A[1][240] = 5'b11111;
assign A[1][241] = 5'b11101;
assign A[1][242] = 5'b11110;
assign A[1][243] = 5'b11101;
assign A[1][244] = 5'b11111;
assign A[1][245] = 5'b00001;
assign A[1][246] = 5'b00000;
assign A[1][247] = 5'b11111;
assign A[1][248] = 5'b11111;
assign A[1][249] = 5'b00000;
assign A[1][250] = 5'b11111;
assign A[1][251] = 5'b11111;
assign A[1][252] = 5'b11111;
assign A[1][253] = 5'b00001;
assign A[1][254] = 5'b11111;
assign A[1][255] = 5'b11110;
assign A[2][0] = 5'b11010;
assign A[2][1] = 5'b00000;
assign A[2][2] = 5'b11111;
assign A[2][3] = 5'b00000;
assign A[2][4] = 5'b11111;
assign A[2][5] = 5'b11101;
assign A[2][6] = 5'b11111;
assign A[2][7] = 5'b11101;
assign A[2][8] = 5'b00001;
assign A[2][9] = 5'b11110;
assign A[2][10] = 5'b11110;
assign A[2][11] = 5'b11110;
assign A[2][12] = 5'b11111;
assign A[2][13] = 5'b11011;
assign A[2][14] = 5'b11111;
assign A[2][15] = 5'b11111;
assign A[2][16] = 5'b11111;
assign A[2][17] = 5'b11111;
assign A[2][18] = 5'b11110;
assign A[2][19] = 5'b11111;
assign A[2][20] = 5'b11101;
assign A[2][21] = 5'b00010;
assign A[2][22] = 5'b11110;
assign A[2][23] = 5'b00000;
assign A[2][24] = 5'b00000;
assign A[2][25] = 5'b11110;
assign A[2][26] = 5'b00000;
assign A[2][27] = 5'b11110;
assign A[2][28] = 5'b00000;
assign A[2][29] = 5'b00010;
assign A[2][30] = 5'b11111;
assign A[2][31] = 5'b11110;
assign A[2][32] = 5'b11100;
assign A[2][33] = 5'b11111;
assign A[2][34] = 5'b11111;
assign A[2][35] = 5'b11111;
assign A[2][36] = 5'b00000;
assign A[2][37] = 5'b11110;
assign A[2][38] = 5'b00000;
assign A[2][39] = 5'b11111;
assign A[2][40] = 5'b11111;
assign A[2][41] = 5'b00000;
assign A[2][42] = 5'b00001;
assign A[2][43] = 5'b11111;
assign A[2][44] = 5'b11110;
assign A[2][45] = 5'b11101;
assign A[2][46] = 5'b11111;
assign A[2][47] = 5'b00000;
assign A[2][48] = 5'b00001;
assign A[2][49] = 5'b00000;
assign A[2][50] = 5'b00001;
assign A[2][51] = 5'b11111;
assign A[2][52] = 5'b11111;
assign A[2][53] = 5'b00000;
assign A[2][54] = 5'b00001;
assign A[2][55] = 5'b00001;
assign A[2][56] = 5'b00000;
assign A[2][57] = 5'b00001;
assign A[2][58] = 5'b11111;
assign A[2][59] = 5'b00010;
assign A[2][60] = 5'b00001;
assign A[2][61] = 5'b11111;
assign A[2][62] = 5'b11111;
assign A[2][63] = 5'b00001;
assign A[2][64] = 5'b11111;
assign A[2][65] = 5'b00000;
assign A[2][66] = 5'b00010;
assign A[2][67] = 5'b00001;
assign A[2][68] = 5'b00000;
assign A[2][69] = 5'b11111;
assign A[2][70] = 5'b11111;
assign A[2][71] = 5'b00010;
assign A[2][72] = 5'b00001;
assign A[2][73] = 5'b00001;
assign A[2][74] = 5'b11111;
assign A[2][75] = 5'b00000;
assign A[2][76] = 5'b00000;
assign A[2][77] = 5'b00000;
assign A[2][78] = 5'b11111;
assign A[2][79] = 5'b11101;
assign A[2][80] = 5'b11111;
assign A[2][81] = 5'b11110;
assign A[2][82] = 5'b00001;
assign A[2][83] = 5'b11100;
assign A[2][84] = 5'b00010;
assign A[2][85] = 5'b11111;
assign A[2][86] = 5'b00000;
assign A[2][87] = 5'b00000;
assign A[2][88] = 5'b00011;
assign A[2][89] = 5'b00000;
assign A[2][90] = 5'b00011;
assign A[2][91] = 5'b11110;
assign A[2][92] = 5'b00000;
assign A[2][93] = 5'b00001;
assign A[2][94] = 5'b11110;
assign A[2][95] = 5'b11111;
assign A[2][96] = 5'b11110;
assign A[2][97] = 5'b00011;
assign A[2][98] = 5'b11110;
assign A[2][99] = 5'b00001;
assign A[2][100] = 5'b00001;
assign A[2][101] = 5'b11110;
assign A[2][102] = 5'b11111;
assign A[2][103] = 5'b00000;
assign A[2][104] = 5'b00010;
assign A[2][105] = 5'b11111;
assign A[2][106] = 5'b00001;
assign A[2][107] = 5'b00000;
assign A[2][108] = 5'b00001;
assign A[2][109] = 5'b11111;
assign A[2][110] = 5'b00011;
assign A[2][111] = 5'b00000;
assign A[2][112] = 5'b00011;
assign A[2][113] = 5'b11110;
assign A[2][114] = 5'b00010;
assign A[2][115] = 5'b11111;
assign A[2][116] = 5'b00001;
assign A[2][117] = 5'b00001;
assign A[2][118] = 5'b11110;
assign A[2][119] = 5'b00010;
assign A[2][120] = 5'b00000;
assign A[2][121] = 5'b00010;
assign A[2][122] = 5'b00001;
assign A[2][123] = 5'b00000;
assign A[2][124] = 5'b00001;
assign A[2][125] = 5'b00001;
assign A[2][126] = 5'b00000;
assign A[2][127] = 5'b11111;
assign A[2][128] = 5'b11111;
assign A[2][129] = 5'b00011;
assign A[2][130] = 5'b00001;
assign A[2][131] = 5'b00010;
assign A[2][132] = 5'b00001;
assign A[2][133] = 5'b00000;
assign A[2][134] = 5'b11110;
assign A[2][135] = 5'b00000;
assign A[2][136] = 5'b11111;
assign A[2][137] = 5'b00100;
assign A[2][138] = 5'b00001;
assign A[2][139] = 5'b00000;
assign A[2][140] = 5'b11110;
assign A[2][141] = 5'b00001;
assign A[2][142] = 5'b00000;
assign A[2][143] = 5'b11111;
assign A[2][144] = 5'b11101;
assign A[2][145] = 5'b00011;
assign A[2][146] = 5'b11101;
assign A[2][147] = 5'b11111;
assign A[2][148] = 5'b00010;
assign A[2][149] = 5'b00001;
assign A[2][150] = 5'b00000;
assign A[2][151] = 5'b00000;
assign A[2][152] = 5'b00000;
assign A[2][153] = 5'b11111;
assign A[2][154] = 5'b00001;
assign A[2][155] = 5'b00010;
assign A[2][156] = 5'b00001;
assign A[2][157] = 5'b00000;
assign A[2][158] = 5'b00010;
assign A[2][159] = 5'b11101;
assign A[2][160] = 5'b00000;
assign A[2][161] = 5'b00100;
assign A[2][162] = 5'b00000;
assign A[2][163] = 5'b00001;
assign A[2][164] = 5'b11111;
assign A[2][165] = 5'b00001;
assign A[2][166] = 5'b00001;
assign A[2][167] = 5'b00011;
assign A[2][168] = 5'b00010;
assign A[2][169] = 5'b00011;
assign A[2][170] = 5'b00000;
assign A[2][171] = 5'b00001;
assign A[2][172] = 5'b00010;
assign A[2][173] = 5'b11111;
assign A[2][174] = 5'b11110;
assign A[2][175] = 5'b00001;
assign A[2][176] = 5'b11111;
assign A[2][177] = 5'b11110;
assign A[2][178] = 5'b11111;
assign A[2][179] = 5'b11111;
assign A[2][180] = 5'b11110;
assign A[2][181] = 5'b00011;
assign A[2][182] = 5'b00001;
assign A[2][183] = 5'b00001;
assign A[2][184] = 5'b00000;
assign A[2][185] = 5'b00000;
assign A[2][186] = 5'b00001;
assign A[2][187] = 5'b00001;
assign A[2][188] = 5'b00001;
assign A[2][189] = 5'b11111;
assign A[2][190] = 5'b11111;
assign A[2][191] = 5'b00001;
assign A[2][192] = 5'b00010;
assign A[2][193] = 5'b11111;
assign A[2][194] = 5'b00010;
assign A[2][195] = 5'b00010;
assign A[2][196] = 5'b00001;
assign A[2][197] = 5'b00001;
assign A[2][198] = 5'b00000;
assign A[2][199] = 5'b00000;
assign A[2][200] = 5'b11110;
assign A[2][201] = 5'b00011;
assign A[2][202] = 5'b00000;
assign A[2][203] = 5'b00011;
assign A[2][204] = 5'b00001;
assign A[2][205] = 5'b00001;
assign A[2][206] = 5'b00001;
assign A[2][207] = 5'b11111;
assign A[2][208] = 5'b00000;
assign A[2][209] = 5'b00001;
assign A[2][210] = 5'b11110;
assign A[2][211] = 5'b00010;
assign A[2][212] = 5'b00000;
assign A[2][213] = 5'b11111;
assign A[2][214] = 5'b11101;
assign A[2][215] = 5'b11110;
assign A[2][216] = 5'b11111;
assign A[2][217] = 5'b11110;
assign A[2][218] = 5'b11111;
assign A[2][219] = 5'b11110;
assign A[2][220] = 5'b00011;
assign A[2][221] = 5'b00001;
assign A[2][222] = 5'b11111;
assign A[2][223] = 5'b00000;
assign A[2][224] = 5'b11111;
assign A[2][225] = 5'b11111;
assign A[2][226] = 5'b00001;
assign A[2][227] = 5'b11111;
assign A[2][228] = 5'b11100;
assign A[2][229] = 5'b00000;
assign A[2][230] = 5'b11111;
assign A[2][231] = 5'b11110;
assign A[2][232] = 5'b11111;
assign A[2][233] = 5'b11110;
assign A[2][234] = 5'b11100;
assign A[2][235] = 5'b11111;
assign A[2][236] = 5'b11100;
assign A[2][237] = 5'b00000;
assign A[2][238] = 5'b11111;
assign A[2][239] = 5'b00001;
assign A[2][240] = 5'b11111;
assign A[2][241] = 5'b00000;
assign A[2][242] = 5'b11110;
assign A[2][243] = 5'b11101;
assign A[2][244] = 5'b11100;
assign A[2][245] = 5'b11111;
assign A[2][246] = 5'b00000;
assign A[2][247] = 5'b11101;
assign A[2][248] = 5'b00000;
assign A[2][249] = 5'b00000;
assign A[2][250] = 5'b00001;
assign A[2][251] = 5'b00010;
assign A[2][252] = 5'b11111;
assign A[2][253] = 5'b11111;
assign A[2][254] = 5'b11110;
assign A[2][255] = 5'b00000;
assign A[3][0] = 5'b00000;
assign A[3][1] = 5'b00001;
assign A[3][2] = 5'b11111;
assign A[3][3] = 5'b00000;
assign A[3][4] = 5'b00001;
assign A[3][5] = 5'b11110;
assign A[3][6] = 5'b11101;
assign A[3][7] = 5'b11111;
assign A[3][8] = 5'b00010;
assign A[3][9] = 5'b11110;
assign A[3][10] = 5'b11111;
assign A[3][11] = 5'b11111;
assign A[3][12] = 5'b00000;
assign A[3][13] = 5'b11111;
assign A[3][14] = 5'b00010;
assign A[3][15] = 5'b00011;
assign A[3][16] = 5'b11111;
assign A[3][17] = 5'b00000;
assign A[3][18] = 5'b11110;
assign A[3][19] = 5'b00000;
assign A[3][20] = 5'b11110;
assign A[3][21] = 5'b00000;
assign A[3][22] = 5'b00000;
assign A[3][23] = 5'b00000;
assign A[3][24] = 5'b00000;
assign A[3][25] = 5'b00001;
assign A[3][26] = 5'b11110;
assign A[3][27] = 5'b00000;
assign A[3][28] = 5'b00010;
assign A[3][29] = 5'b11110;
assign A[3][30] = 5'b00000;
assign A[3][31] = 5'b00001;
assign A[3][32] = 5'b00000;
assign A[3][33] = 5'b11110;
assign A[3][34] = 5'b11111;
assign A[3][35] = 5'b11111;
assign A[3][36] = 5'b11111;
assign A[3][37] = 5'b11111;
assign A[3][38] = 5'b00001;
assign A[3][39] = 5'b11110;
assign A[3][40] = 5'b00000;
assign A[3][41] = 5'b11111;
assign A[3][42] = 5'b00000;
assign A[3][43] = 5'b11111;
assign A[3][44] = 5'b00001;
assign A[3][45] = 5'b00010;
assign A[3][46] = 5'b00001;
assign A[3][47] = 5'b11110;
assign A[3][48] = 5'b11111;
assign A[3][49] = 5'b11111;
assign A[3][50] = 5'b11111;
assign A[3][51] = 5'b00000;
assign A[3][52] = 5'b11111;
assign A[3][53] = 5'b00010;
assign A[3][54] = 5'b11101;
assign A[3][55] = 5'b11111;
assign A[3][56] = 5'b00011;
assign A[3][57] = 5'b00001;
assign A[3][58] = 5'b00001;
assign A[3][59] = 5'b00000;
assign A[3][60] = 5'b00000;
assign A[3][61] = 5'b00001;
assign A[3][62] = 5'b00000;
assign A[3][63] = 5'b00000;
assign A[3][64] = 5'b00001;
assign A[3][65] = 5'b00010;
assign A[3][66] = 5'b11111;
assign A[3][67] = 5'b11111;
assign A[3][68] = 5'b00001;
assign A[3][69] = 5'b00010;
assign A[3][70] = 5'b00011;
assign A[3][71] = 5'b00000;
assign A[3][72] = 5'b00011;
assign A[3][73] = 5'b11110;
assign A[3][74] = 5'b11100;
assign A[3][75] = 5'b00000;
assign A[3][76] = 5'b00010;
assign A[3][77] = 5'b00001;
assign A[3][78] = 5'b11110;
assign A[3][79] = 5'b00010;
assign A[3][80] = 5'b11111;
assign A[3][81] = 5'b00001;
assign A[3][82] = 5'b00000;
assign A[3][83] = 5'b11111;
assign A[3][84] = 5'b11111;
assign A[3][85] = 5'b00010;
assign A[3][86] = 5'b00001;
assign A[3][87] = 5'b00001;
assign A[3][88] = 5'b00000;
assign A[3][89] = 5'b11110;
assign A[3][90] = 5'b00001;
assign A[3][91] = 5'b00010;
assign A[3][92] = 5'b11111;
assign A[3][93] = 5'b11111;
assign A[3][94] = 5'b00000;
assign A[3][95] = 5'b11111;
assign A[3][96] = 5'b11111;
assign A[3][97] = 5'b00000;
assign A[3][98] = 5'b11111;
assign A[3][99] = 5'b11111;
assign A[3][100] = 5'b11110;
assign A[3][101] = 5'b11111;
assign A[3][102] = 5'b00010;
assign A[3][103] = 5'b00000;
assign A[3][104] = 5'b00001;
assign A[3][105] = 5'b11111;
assign A[3][106] = 5'b00010;
assign A[3][107] = 5'b00000;
assign A[3][108] = 5'b00100;
assign A[3][109] = 5'b00011;
assign A[3][110] = 5'b11101;
assign A[3][111] = 5'b11111;
assign A[3][112] = 5'b00000;
assign A[3][113] = 5'b00001;
assign A[3][114] = 5'b11101;
assign A[3][115] = 5'b11111;
assign A[3][116] = 5'b00000;
assign A[3][117] = 5'b11111;
assign A[3][118] = 5'b00000;
assign A[3][119] = 5'b11111;
assign A[3][120] = 5'b11110;
assign A[3][121] = 5'b00001;
assign A[3][122] = 5'b00000;
assign A[3][123] = 5'b00010;
assign A[3][124] = 5'b00000;
assign A[3][125] = 5'b00000;
assign A[3][126] = 5'b00000;
assign A[3][127] = 5'b00001;
assign A[3][128] = 5'b11111;
assign A[3][129] = 5'b11110;
assign A[3][130] = 5'b11110;
assign A[3][131] = 5'b00000;
assign A[3][132] = 5'b11111;
assign A[3][133] = 5'b00000;
assign A[3][134] = 5'b00000;
assign A[3][135] = 5'b11110;
assign A[3][136] = 5'b00010;
assign A[3][137] = 5'b00001;
assign A[3][138] = 5'b00000;
assign A[3][139] = 5'b00001;
assign A[3][140] = 5'b11110;
assign A[3][141] = 5'b11110;
assign A[3][142] = 5'b11111;
assign A[3][143] = 5'b00000;
assign A[3][144] = 5'b11110;
assign A[3][145] = 5'b00010;
assign A[3][146] = 5'b11111;
assign A[3][147] = 5'b11111;
assign A[3][148] = 5'b00001;
assign A[3][149] = 5'b00011;
assign A[3][150] = 5'b00010;
assign A[3][151] = 5'b11111;
assign A[3][152] = 5'b00001;
assign A[3][153] = 5'b00000;
assign A[3][154] = 5'b00010;
assign A[3][155] = 5'b11111;
assign A[3][156] = 5'b11111;
assign A[3][157] = 5'b11111;
assign A[3][158] = 5'b11110;
assign A[3][159] = 5'b11110;
assign A[3][160] = 5'b11111;
assign A[3][161] = 5'b11101;
assign A[3][162] = 5'b00001;
assign A[3][163] = 5'b00000;
assign A[3][164] = 5'b00001;
assign A[3][165] = 5'b11111;
assign A[3][166] = 5'b00000;
assign A[3][167] = 5'b00000;
assign A[3][168] = 5'b11111;
assign A[3][169] = 5'b00000;
assign A[3][170] = 5'b11101;
assign A[3][171] = 5'b00000;
assign A[3][172] = 5'b00001;
assign A[3][173] = 5'b00000;
assign A[3][174] = 5'b11110;
assign A[3][175] = 5'b11101;
assign A[3][176] = 5'b00000;
assign A[3][177] = 5'b00000;
assign A[3][178] = 5'b00001;
assign A[3][179] = 5'b00010;
assign A[3][180] = 5'b00010;
assign A[3][181] = 5'b00001;
assign A[3][182] = 5'b00000;
assign A[3][183] = 5'b11111;
assign A[3][184] = 5'b11110;
assign A[3][185] = 5'b11111;
assign A[3][186] = 5'b00010;
assign A[3][187] = 5'b00010;
assign A[3][188] = 5'b11111;
assign A[3][189] = 5'b00000;
assign A[3][190] = 5'b00000;
assign A[3][191] = 5'b11110;
assign A[3][192] = 5'b00001;
assign A[3][193] = 5'b00000;
assign A[3][194] = 5'b11110;
assign A[3][195] = 5'b00010;
assign A[3][196] = 5'b00000;
assign A[3][197] = 5'b00010;
assign A[3][198] = 5'b11101;
assign A[3][199] = 5'b00000;
assign A[3][200] = 5'b11111;
assign A[3][201] = 5'b00001;
assign A[3][202] = 5'b00000;
assign A[3][203] = 5'b11110;
assign A[3][204] = 5'b00001;
assign A[3][205] = 5'b11111;
assign A[3][206] = 5'b11110;
assign A[3][207] = 5'b00000;
assign A[3][208] = 5'b00000;
assign A[3][209] = 5'b11111;
assign A[3][210] = 5'b11111;
assign A[3][211] = 5'b00010;
assign A[3][212] = 5'b11111;
assign A[3][213] = 5'b00000;
assign A[3][214] = 5'b11110;
assign A[3][215] = 5'b11111;
assign A[3][216] = 5'b00010;
assign A[3][217] = 5'b00000;
assign A[3][218] = 5'b11111;
assign A[3][219] = 5'b11111;
assign A[3][220] = 5'b11111;
assign A[3][221] = 5'b11111;
assign A[3][222] = 5'b11111;
assign A[3][223] = 5'b00001;
assign A[3][224] = 5'b00001;
assign A[3][225] = 5'b00001;
assign A[3][226] = 5'b11111;
assign A[3][227] = 5'b00000;
assign A[3][228] = 5'b00000;
assign A[3][229] = 5'b11111;
assign A[3][230] = 5'b11110;
assign A[3][231] = 5'b00000;
assign A[3][232] = 5'b00000;
assign A[3][233] = 5'b00001;
assign A[3][234] = 5'b00000;
assign A[3][235] = 5'b00001;
assign A[3][236] = 5'b00000;
assign A[3][237] = 5'b00000;
assign A[3][238] = 5'b11111;
assign A[3][239] = 5'b11111;
assign A[3][240] = 5'b00010;
assign A[3][241] = 5'b00000;
assign A[3][242] = 5'b11101;
assign A[3][243] = 5'b00010;
assign A[3][244] = 5'b00010;
assign A[3][245] = 5'b00000;
assign A[3][246] = 5'b11111;
assign A[3][247] = 5'b00001;
assign A[3][248] = 5'b11111;
assign A[3][249] = 5'b00001;
assign A[3][250] = 5'b00000;
assign A[3][251] = 5'b11110;
assign A[3][252] = 5'b00000;
assign A[3][253] = 5'b00000;
assign A[3][254] = 5'b00000;
assign A[3][255] = 5'b11111;
assign A[4][0] = 5'b11111;
assign A[4][1] = 5'b11111;
assign A[4][2] = 5'b00000;
assign A[4][3] = 5'b00001;
assign A[4][4] = 5'b00000;
assign A[4][5] = 5'b11110;
assign A[4][6] = 5'b11110;
assign A[4][7] = 5'b11111;
assign A[4][8] = 5'b00001;
assign A[4][9] = 5'b11111;
assign A[4][10] = 5'b11111;
assign A[4][11] = 5'b11101;
assign A[4][12] = 5'b00000;
assign A[4][13] = 5'b00000;
assign A[4][14] = 5'b00001;
assign A[4][15] = 5'b00001;
assign A[4][16] = 5'b11111;
assign A[4][17] = 5'b00000;
assign A[4][18] = 5'b00000;
assign A[4][19] = 5'b11111;
assign A[4][20] = 5'b11111;
assign A[4][21] = 5'b00001;
assign A[4][22] = 5'b00000;
assign A[4][23] = 5'b11110;
assign A[4][24] = 5'b00001;
assign A[4][25] = 5'b11111;
assign A[4][26] = 5'b11101;
assign A[4][27] = 5'b00000;
assign A[4][28] = 5'b11111;
assign A[4][29] = 5'b00010;
assign A[4][30] = 5'b00011;
assign A[4][31] = 5'b11101;
assign A[4][32] = 5'b11110;
assign A[4][33] = 5'b11110;
assign A[4][34] = 5'b11110;
assign A[4][35] = 5'b11111;
assign A[4][36] = 5'b00000;
assign A[4][37] = 5'b11101;
assign A[4][38] = 5'b00000;
assign A[4][39] = 5'b11111;
assign A[4][40] = 5'b11110;
assign A[4][41] = 5'b00000;
assign A[4][42] = 5'b11101;
assign A[4][43] = 5'b11110;
assign A[4][44] = 5'b00100;
assign A[4][45] = 5'b00000;
assign A[4][46] = 5'b00001;
assign A[4][47] = 5'b00000;
assign A[4][48] = 5'b11111;
assign A[4][49] = 5'b00010;
assign A[4][50] = 5'b00000;
assign A[4][51] = 5'b11111;
assign A[4][52] = 5'b11110;
assign A[4][53] = 5'b11111;
assign A[4][54] = 5'b11111;
assign A[4][55] = 5'b11100;
assign A[4][56] = 5'b00011;
assign A[4][57] = 5'b00001;
assign A[4][58] = 5'b00001;
assign A[4][59] = 5'b11111;
assign A[4][60] = 5'b11111;
assign A[4][61] = 5'b00010;
assign A[4][62] = 5'b00001;
assign A[4][63] = 5'b00000;
assign A[4][64] = 5'b00010;
assign A[4][65] = 5'b00001;
assign A[4][66] = 5'b11110;
assign A[4][67] = 5'b11110;
assign A[4][68] = 5'b11111;
assign A[4][69] = 5'b11111;
assign A[4][70] = 5'b11100;
assign A[4][71] = 5'b00010;
assign A[4][72] = 5'b00000;
assign A[4][73] = 5'b11111;
assign A[4][74] = 5'b00010;
assign A[4][75] = 5'b00000;
assign A[4][76] = 5'b11110;
assign A[4][77] = 5'b00001;
assign A[4][78] = 5'b11011;
assign A[4][79] = 5'b11111;
assign A[4][80] = 5'b11110;
assign A[4][81] = 5'b00010;
assign A[4][82] = 5'b11111;
assign A[4][83] = 5'b11111;
assign A[4][84] = 5'b11111;
assign A[4][85] = 5'b00010;
assign A[4][86] = 5'b00011;
assign A[4][87] = 5'b00001;
assign A[4][88] = 5'b00000;
assign A[4][89] = 5'b00000;
assign A[4][90] = 5'b00000;
assign A[4][91] = 5'b11110;
assign A[4][92] = 5'b00001;
assign A[4][93] = 5'b00000;
assign A[4][94] = 5'b11110;
assign A[4][95] = 5'b11111;
assign A[4][96] = 5'b11101;
assign A[4][97] = 5'b00001;
assign A[4][98] = 5'b00010;
assign A[4][99] = 5'b00000;
assign A[4][100] = 5'b00000;
assign A[4][101] = 5'b00010;
assign A[4][102] = 5'b00001;
assign A[4][103] = 5'b11110;
assign A[4][104] = 5'b00001;
assign A[4][105] = 5'b00000;
assign A[4][106] = 5'b11110;
assign A[4][107] = 5'b00000;
assign A[4][108] = 5'b00000;
assign A[4][109] = 5'b00000;
assign A[4][110] = 5'b11101;
assign A[4][111] = 5'b11111;
assign A[4][112] = 5'b11111;
assign A[4][113] = 5'b11111;
assign A[4][114] = 5'b00010;
assign A[4][115] = 5'b00000;
assign A[4][116] = 5'b00011;
assign A[4][117] = 5'b00001;
assign A[4][118] = 5'b11111;
assign A[4][119] = 5'b11111;
assign A[4][120] = 5'b00000;
assign A[4][121] = 5'b00000;
assign A[4][122] = 5'b00000;
assign A[4][123] = 5'b00000;
assign A[4][124] = 5'b11110;
assign A[4][125] = 5'b11110;
assign A[4][126] = 5'b11110;
assign A[4][127] = 5'b11101;
assign A[4][128] = 5'b00000;
assign A[4][129] = 5'b11110;
assign A[4][130] = 5'b00000;
assign A[4][131] = 5'b00100;
assign A[4][132] = 5'b00011;
assign A[4][133] = 5'b11111;
assign A[4][134] = 5'b11110;
assign A[4][135] = 5'b00000;
assign A[4][136] = 5'b11110;
assign A[4][137] = 5'b00010;
assign A[4][138] = 5'b00001;
assign A[4][139] = 5'b00000;
assign A[4][140] = 5'b11110;
assign A[4][141] = 5'b00000;
assign A[4][142] = 5'b00001;
assign A[4][143] = 5'b00001;
assign A[4][144] = 5'b11111;
assign A[4][145] = 5'b11111;
assign A[4][146] = 5'b00001;
assign A[4][147] = 5'b00000;
assign A[4][148] = 5'b11110;
assign A[4][149] = 5'b11111;
assign A[4][150] = 5'b11111;
assign A[4][151] = 5'b00000;
assign A[4][152] = 5'b00000;
assign A[4][153] = 5'b00000;
assign A[4][154] = 5'b00001;
assign A[4][155] = 5'b11110;
assign A[4][156] = 5'b00000;
assign A[4][157] = 5'b11111;
assign A[4][158] = 5'b11110;
assign A[4][159] = 5'b00001;
assign A[4][160] = 5'b00010;
assign A[4][161] = 5'b00001;
assign A[4][162] = 5'b00010;
assign A[4][163] = 5'b00010;
assign A[4][164] = 5'b11110;
assign A[4][165] = 5'b00000;
assign A[4][166] = 5'b11111;
assign A[4][167] = 5'b11110;
assign A[4][168] = 5'b11111;
assign A[4][169] = 5'b11110;
assign A[4][170] = 5'b00000;
assign A[4][171] = 5'b00001;
assign A[4][172] = 5'b11111;
assign A[4][173] = 5'b00010;
assign A[4][174] = 5'b11111;
assign A[4][175] = 5'b00001;
assign A[4][176] = 5'b00001;
assign A[4][177] = 5'b00011;
assign A[4][178] = 5'b11111;
assign A[4][179] = 5'b00001;
assign A[4][180] = 5'b11111;
assign A[4][181] = 5'b00000;
assign A[4][182] = 5'b11101;
assign A[4][183] = 5'b11111;
assign A[4][184] = 5'b00000;
assign A[4][185] = 5'b00000;
assign A[4][186] = 5'b00001;
assign A[4][187] = 5'b00001;
assign A[4][188] = 5'b00011;
assign A[4][189] = 5'b00000;
assign A[4][190] = 5'b00010;
assign A[4][191] = 5'b00001;
assign A[4][192] = 5'b11110;
assign A[4][193] = 5'b00000;
assign A[4][194] = 5'b00001;
assign A[4][195] = 5'b00001;
assign A[4][196] = 5'b11110;
assign A[4][197] = 5'b11101;
assign A[4][198] = 5'b00000;
assign A[4][199] = 5'b00010;
assign A[4][200] = 5'b00000;
assign A[4][201] = 5'b00000;
assign A[4][202] = 5'b11111;
assign A[4][203] = 5'b00000;
assign A[4][204] = 5'b11111;
assign A[4][205] = 5'b00011;
assign A[4][206] = 5'b00000;
assign A[4][207] = 5'b00010;
assign A[4][208] = 5'b00001;
assign A[4][209] = 5'b11101;
assign A[4][210] = 5'b11111;
assign A[4][211] = 5'b00001;
assign A[4][212] = 5'b11111;
assign A[4][213] = 5'b00000;
assign A[4][214] = 5'b11111;
assign A[4][215] = 5'b11111;
assign A[4][216] = 5'b00000;
assign A[4][217] = 5'b00011;
assign A[4][218] = 5'b11111;
assign A[4][219] = 5'b00010;
assign A[4][220] = 5'b00010;
assign A[4][221] = 5'b11111;
assign A[4][222] = 5'b00000;
assign A[4][223] = 5'b00010;
assign A[4][224] = 5'b11111;
assign A[4][225] = 5'b11111;
assign A[4][226] = 5'b00001;
assign A[4][227] = 5'b00000;
assign A[4][228] = 5'b00010;
assign A[4][229] = 5'b11111;
assign A[4][230] = 5'b11111;
assign A[4][231] = 5'b00000;
assign A[4][232] = 5'b11111;
assign A[4][233] = 5'b11110;
assign A[4][234] = 5'b11111;
assign A[4][235] = 5'b00001;
assign A[4][236] = 5'b00000;
assign A[4][237] = 5'b00001;
assign A[4][238] = 5'b11110;
assign A[4][239] = 5'b00010;
assign A[4][240] = 5'b00011;
assign A[4][241] = 5'b00000;
assign A[4][242] = 5'b00001;
assign A[4][243] = 5'b11111;
assign A[4][244] = 5'b11111;
assign A[4][245] = 5'b00001;
assign A[4][246] = 5'b00001;
assign A[4][247] = 5'b00011;
assign A[4][248] = 5'b11111;
assign A[4][249] = 5'b11111;
assign A[4][250] = 5'b00000;
assign A[4][251] = 5'b00001;
assign A[4][252] = 5'b00001;
assign A[4][253] = 5'b00001;
assign A[4][254] = 5'b11111;
assign A[4][255] = 5'b00001;
assign A[5][0] = 5'b11110;
assign A[5][1] = 5'b00000;
assign A[5][2] = 5'b11111;
assign A[5][3] = 5'b11111;
assign A[5][4] = 5'b00000;
assign A[5][5] = 5'b11111;
assign A[5][6] = 5'b11111;
assign A[5][7] = 5'b11111;
assign A[5][8] = 5'b11111;
assign A[5][9] = 5'b00000;
assign A[5][10] = 5'b11111;
assign A[5][11] = 5'b11111;
assign A[5][12] = 5'b11101;
assign A[5][13] = 5'b11101;
assign A[5][14] = 5'b11111;
assign A[5][15] = 5'b11110;
assign A[5][16] = 5'b11111;
assign A[5][17] = 5'b00001;
assign A[5][18] = 5'b11111;
assign A[5][19] = 5'b00010;
assign A[5][20] = 5'b00001;
assign A[5][21] = 5'b00000;
assign A[5][22] = 5'b00010;
assign A[5][23] = 5'b11111;
assign A[5][24] = 5'b11110;
assign A[5][25] = 5'b11111;
assign A[5][26] = 5'b11111;
assign A[5][27] = 5'b00000;
assign A[5][28] = 5'b00000;
assign A[5][29] = 5'b11111;
assign A[5][30] = 5'b11111;
assign A[5][31] = 5'b11111;
assign A[5][32] = 5'b00000;
assign A[5][33] = 5'b00000;
assign A[5][34] = 5'b11111;
assign A[5][35] = 5'b00001;
assign A[5][36] = 5'b00000;
assign A[5][37] = 5'b00001;
assign A[5][38] = 5'b00010;
assign A[5][39] = 5'b00011;
assign A[5][40] = 5'b11111;
assign A[5][41] = 5'b11110;
assign A[5][42] = 5'b11011;
assign A[5][43] = 5'b11110;
assign A[5][44] = 5'b11101;
assign A[5][45] = 5'b11110;
assign A[5][46] = 5'b00000;
assign A[5][47] = 5'b00000;
assign A[5][48] = 5'b00000;
assign A[5][49] = 5'b11111;
assign A[5][50] = 5'b11111;
assign A[5][51] = 5'b00010;
assign A[5][52] = 5'b11111;
assign A[5][53] = 5'b00001;
assign A[5][54] = 5'b00010;
assign A[5][55] = 5'b00000;
assign A[5][56] = 5'b00000;
assign A[5][57] = 5'b00000;
assign A[5][58] = 5'b11111;
assign A[5][59] = 5'b11111;
assign A[5][60] = 5'b11110;
assign A[5][61] = 5'b00000;
assign A[5][62] = 5'b00001;
assign A[5][63] = 5'b00010;
assign A[5][64] = 5'b00010;
assign A[5][65] = 5'b11111;
assign A[5][66] = 5'b00000;
assign A[5][67] = 5'b00001;
assign A[5][68] = 5'b00001;
assign A[5][69] = 5'b00001;
assign A[5][70] = 5'b00011;
assign A[5][71] = 5'b11110;
assign A[5][72] = 5'b11111;
assign A[5][73] = 5'b11110;
assign A[5][74] = 5'b00011;
assign A[5][75] = 5'b11111;
assign A[5][76] = 5'b11111;
assign A[5][77] = 5'b00000;
assign A[5][78] = 5'b11111;
assign A[5][79] = 5'b00000;
assign A[5][80] = 5'b00000;
assign A[5][81] = 5'b00000;
assign A[5][82] = 5'b11110;
assign A[5][83] = 5'b11111;
assign A[5][84] = 5'b00010;
assign A[5][85] = 5'b00001;
assign A[5][86] = 5'b00001;
assign A[5][87] = 5'b00001;
assign A[5][88] = 5'b00001;
assign A[5][89] = 5'b11110;
assign A[5][90] = 5'b11110;
assign A[5][91] = 5'b11110;
assign A[5][92] = 5'b00001;
assign A[5][93] = 5'b00000;
assign A[5][94] = 5'b00000;
assign A[5][95] = 5'b11111;
assign A[5][96] = 5'b00001;
assign A[5][97] = 5'b00000;
assign A[5][98] = 5'b11111;
assign A[5][99] = 5'b00011;
assign A[5][100] = 5'b00001;
assign A[5][101] = 5'b11111;
assign A[5][102] = 5'b00001;
assign A[5][103] = 5'b00010;
assign A[5][104] = 5'b00000;
assign A[5][105] = 5'b00000;
assign A[5][106] = 5'b00000;
assign A[5][107] = 5'b11110;
assign A[5][108] = 5'b11101;
assign A[5][109] = 5'b00000;
assign A[5][110] = 5'b00011;
assign A[5][111] = 5'b00001;
assign A[5][112] = 5'b00000;
assign A[5][113] = 5'b11111;
assign A[5][114] = 5'b00010;
assign A[5][115] = 5'b00000;
assign A[5][116] = 5'b00000;
assign A[5][117] = 5'b00000;
assign A[5][118] = 5'b00011;
assign A[5][119] = 5'b00000;
assign A[5][120] = 5'b11111;
assign A[5][121] = 5'b11101;
assign A[5][122] = 5'b00000;
assign A[5][123] = 5'b00000;
assign A[5][124] = 5'b11110;
assign A[5][125] = 5'b11111;
assign A[5][126] = 5'b11111;
assign A[5][127] = 5'b11111;
assign A[5][128] = 5'b00001;
assign A[5][129] = 5'b11111;
assign A[5][130] = 5'b00010;
assign A[5][131] = 5'b00000;
assign A[5][132] = 5'b00001;
assign A[5][133] = 5'b11111;
assign A[5][134] = 5'b00001;
assign A[5][135] = 5'b00000;
assign A[5][136] = 5'b00000;
assign A[5][137] = 5'b11110;
assign A[5][138] = 5'b00000;
assign A[5][139] = 5'b11110;
assign A[5][140] = 5'b11101;
assign A[5][141] = 5'b11110;
assign A[5][142] = 5'b11110;
assign A[5][143] = 5'b00001;
assign A[5][144] = 5'b11100;
assign A[5][145] = 5'b00000;
assign A[5][146] = 5'b11101;
assign A[5][147] = 5'b11111;
assign A[5][148] = 5'b00000;
assign A[5][149] = 5'b00010;
assign A[5][150] = 5'b00000;
assign A[5][151] = 5'b00001;
assign A[5][152] = 5'b11101;
assign A[5][153] = 5'b00001;
assign A[5][154] = 5'b11101;
assign A[5][155] = 5'b11110;
assign A[5][156] = 5'b11111;
assign A[5][157] = 5'b11111;
assign A[5][158] = 5'b00000;
assign A[5][159] = 5'b11111;
assign A[5][160] = 5'b11110;
assign A[5][161] = 5'b11111;
assign A[5][162] = 5'b11110;
assign A[5][163] = 5'b11111;
assign A[5][164] = 5'b00000;
assign A[5][165] = 5'b00001;
assign A[5][166] = 5'b00010;
assign A[5][167] = 5'b11110;
assign A[5][168] = 5'b00000;
assign A[5][169] = 5'b00011;
assign A[5][170] = 5'b11111;
assign A[5][171] = 5'b11111;
assign A[5][172] = 5'b00000;
assign A[5][173] = 5'b00001;
assign A[5][174] = 5'b11111;
assign A[5][175] = 5'b11101;
assign A[5][176] = 5'b11111;
assign A[5][177] = 5'b11110;
assign A[5][178] = 5'b00001;
assign A[5][179] = 5'b00001;
assign A[5][180] = 5'b11110;
assign A[5][181] = 5'b00010;
assign A[5][182] = 5'b00010;
assign A[5][183] = 5'b00001;
assign A[5][184] = 5'b11111;
assign A[5][185] = 5'b00001;
assign A[5][186] = 5'b00000;
assign A[5][187] = 5'b00010;
assign A[5][188] = 5'b00001;
assign A[5][189] = 5'b00010;
assign A[5][190] = 5'b00001;
assign A[5][191] = 5'b11101;
assign A[5][192] = 5'b11100;
assign A[5][193] = 5'b00001;
assign A[5][194] = 5'b00000;
assign A[5][195] = 5'b00000;
assign A[5][196] = 5'b00011;
assign A[5][197] = 5'b00001;
assign A[5][198] = 5'b00001;
assign A[5][199] = 5'b00000;
assign A[5][200] = 5'b00001;
assign A[5][201] = 5'b00001;
assign A[5][202] = 5'b11110;
assign A[5][203] = 5'b00001;
assign A[5][204] = 5'b00000;
assign A[5][205] = 5'b11111;
assign A[5][206] = 5'b11110;
assign A[5][207] = 5'b00000;
assign A[5][208] = 5'b11111;
assign A[5][209] = 5'b11110;
assign A[5][210] = 5'b11110;
assign A[5][211] = 5'b00000;
assign A[5][212] = 5'b00100;
assign A[5][213] = 5'b00000;
assign A[5][214] = 5'b11111;
assign A[5][215] = 5'b00001;
assign A[5][216] = 5'b11110;
assign A[5][217] = 5'b00001;
assign A[5][218] = 5'b00000;
assign A[5][219] = 5'b00010;
assign A[5][220] = 5'b00000;
assign A[5][221] = 5'b11110;
assign A[5][222] = 5'b00001;
assign A[5][223] = 5'b11110;
assign A[5][224] = 5'b00001;
assign A[5][225] = 5'b00001;
assign A[5][226] = 5'b11111;
assign A[5][227] = 5'b11111;
assign A[5][228] = 5'b11111;
assign A[5][229] = 5'b00000;
assign A[5][230] = 5'b11111;
assign A[5][231] = 5'b11111;
assign A[5][232] = 5'b00001;
assign A[5][233] = 5'b00011;
assign A[5][234] = 5'b00010;
assign A[5][235] = 5'b11110;
assign A[5][236] = 5'b11110;
assign A[5][237] = 5'b11101;
assign A[5][238] = 5'b11111;
assign A[5][239] = 5'b00000;
assign A[5][240] = 5'b11101;
assign A[5][241] = 5'b11110;
assign A[5][242] = 5'b11110;
assign A[5][243] = 5'b11110;
assign A[5][244] = 5'b00001;
assign A[5][245] = 5'b11111;
assign A[5][246] = 5'b00001;
assign A[5][247] = 5'b00000;
assign A[5][248] = 5'b11111;
assign A[5][249] = 5'b00000;
assign A[5][250] = 5'b00001;
assign A[5][251] = 5'b00001;
assign A[5][252] = 5'b00001;
assign A[5][253] = 5'b00000;
assign A[5][254] = 5'b11111;
assign A[5][255] = 5'b11111;
assign A[6][0] = 5'b00010;
assign A[6][1] = 5'b00001;
assign A[6][2] = 5'b11111;
assign A[6][3] = 5'b00000;
assign A[6][4] = 5'b00000;
assign A[6][5] = 5'b00000;
assign A[6][6] = 5'b00000;
assign A[6][7] = 5'b11101;
assign A[6][8] = 5'b00011;
assign A[6][9] = 5'b00001;
assign A[6][10] = 5'b00011;
assign A[6][11] = 5'b00011;
assign A[6][12] = 5'b00010;
assign A[6][13] = 5'b11110;
assign A[6][14] = 5'b11110;
assign A[6][15] = 5'b11110;
assign A[6][16] = 5'b11111;
assign A[6][17] = 5'b00001;
assign A[6][18] = 5'b00000;
assign A[6][19] = 5'b00000;
assign A[6][20] = 5'b00000;
assign A[6][21] = 5'b00001;
assign A[6][22] = 5'b00000;
assign A[6][23] = 5'b00010;
assign A[6][24] = 5'b00001;
assign A[6][25] = 5'b11110;
assign A[6][26] = 5'b00100;
assign A[6][27] = 5'b00000;
assign A[6][28] = 5'b11101;
assign A[6][29] = 5'b00000;
assign A[6][30] = 5'b11111;
assign A[6][31] = 5'b00001;
assign A[6][32] = 5'b11111;
assign A[6][33] = 5'b00010;
assign A[6][34] = 5'b00001;
assign A[6][35] = 5'b00001;
assign A[6][36] = 5'b00000;
assign A[6][37] = 5'b00001;
assign A[6][38] = 5'b00000;
assign A[6][39] = 5'b00000;
assign A[6][40] = 5'b00001;
assign A[6][41] = 5'b11101;
assign A[6][42] = 5'b00000;
assign A[6][43] = 5'b00001;
assign A[6][44] = 5'b00000;
assign A[6][45] = 5'b11111;
assign A[6][46] = 5'b00011;
assign A[6][47] = 5'b11111;
assign A[6][48] = 5'b11111;
assign A[6][49] = 5'b00011;
assign A[6][50] = 5'b00000;
assign A[6][51] = 5'b00010;
assign A[6][52] = 5'b00001;
assign A[6][53] = 5'b00001;
assign A[6][54] = 5'b00000;
assign A[6][55] = 5'b00000;
assign A[6][56] = 5'b00001;
assign A[6][57] = 5'b11111;
assign A[6][58] = 5'b11111;
assign A[6][59] = 5'b11111;
assign A[6][60] = 5'b00011;
assign A[6][61] = 5'b00001;
assign A[6][62] = 5'b00000;
assign A[6][63] = 5'b00010;
assign A[6][64] = 5'b00001;
assign A[6][65] = 5'b00011;
assign A[6][66] = 5'b00011;
assign A[6][67] = 5'b00001;
assign A[6][68] = 5'b00000;
assign A[6][69] = 5'b00001;
assign A[6][70] = 5'b00000;
assign A[6][71] = 5'b00011;
assign A[6][72] = 5'b00000;
assign A[6][73] = 5'b11111;
assign A[6][74] = 5'b00000;
assign A[6][75] = 5'b00001;
assign A[6][76] = 5'b00001;
assign A[6][77] = 5'b00001;
assign A[6][78] = 5'b00000;
assign A[6][79] = 5'b00100;
assign A[6][80] = 5'b00000;
assign A[6][81] = 5'b00011;
assign A[6][82] = 5'b00010;
assign A[6][83] = 5'b00001;
assign A[6][84] = 5'b00010;
assign A[6][85] = 5'b00011;
assign A[6][86] = 5'b00011;
assign A[6][87] = 5'b11110;
assign A[6][88] = 5'b00000;
assign A[6][89] = 5'b00000;
assign A[6][90] = 5'b11110;
assign A[6][91] = 5'b11101;
assign A[6][92] = 5'b00001;
assign A[6][93] = 5'b00010;
assign A[6][94] = 5'b11111;
assign A[6][95] = 5'b00000;
assign A[6][96] = 5'b00010;
assign A[6][97] = 5'b00001;
assign A[6][98] = 5'b00010;
assign A[6][99] = 5'b11111;
assign A[6][100] = 5'b00010;
assign A[6][101] = 5'b00001;
assign A[6][102] = 5'b00001;
assign A[6][103] = 5'b00000;
assign A[6][104] = 5'b00000;
assign A[6][105] = 5'b00011;
assign A[6][106] = 5'b00001;
assign A[6][107] = 5'b00010;
assign A[6][108] = 5'b00000;
assign A[6][109] = 5'b00010;
assign A[6][110] = 5'b00010;
assign A[6][111] = 5'b00001;
assign A[6][112] = 5'b00001;
assign A[6][113] = 5'b00010;
assign A[6][114] = 5'b00011;
assign A[6][115] = 5'b00001;
assign A[6][116] = 5'b00000;
assign A[6][117] = 5'b00010;
assign A[6][118] = 5'b11111;
assign A[6][119] = 5'b00001;
assign A[6][120] = 5'b11111;
assign A[6][121] = 5'b00011;
assign A[6][122] = 5'b11110;
assign A[6][123] = 5'b00000;
assign A[6][124] = 5'b00000;
assign A[6][125] = 5'b11111;
assign A[6][126] = 5'b11111;
assign A[6][127] = 5'b00010;
assign A[6][128] = 5'b11111;
assign A[6][129] = 5'b00010;
assign A[6][130] = 5'b00000;
assign A[6][131] = 5'b00001;
assign A[6][132] = 5'b00010;
assign A[6][133] = 5'b11111;
assign A[6][134] = 5'b00000;
assign A[6][135] = 5'b11110;
assign A[6][136] = 5'b00001;
assign A[6][137] = 5'b00000;
assign A[6][138] = 5'b11110;
assign A[6][139] = 5'b00010;
assign A[6][140] = 5'b11110;
assign A[6][141] = 5'b00000;
assign A[6][142] = 5'b00001;
assign A[6][143] = 5'b00010;
assign A[6][144] = 5'b00011;
assign A[6][145] = 5'b11111;
assign A[6][146] = 5'b00001;
assign A[6][147] = 5'b00000;
assign A[6][148] = 5'b11111;
assign A[6][149] = 5'b00000;
assign A[6][150] = 5'b11111;
assign A[6][151] = 5'b11111;
assign A[6][152] = 5'b00000;
assign A[6][153] = 5'b11110;
assign A[6][154] = 5'b00001;
assign A[6][155] = 5'b00010;
assign A[6][156] = 5'b00001;
assign A[6][157] = 5'b11110;
assign A[6][158] = 5'b11111;
assign A[6][159] = 5'b00001;
assign A[6][160] = 5'b00001;
assign A[6][161] = 5'b11111;
assign A[6][162] = 5'b00000;
assign A[6][163] = 5'b11111;
assign A[6][164] = 5'b11110;
assign A[6][165] = 5'b00001;
assign A[6][166] = 5'b00000;
assign A[6][167] = 5'b00001;
assign A[6][168] = 5'b00001;
assign A[6][169] = 5'b00000;
assign A[6][170] = 5'b11101;
assign A[6][171] = 5'b00011;
assign A[6][172] = 5'b00011;
assign A[6][173] = 5'b00010;
assign A[6][174] = 5'b00000;
assign A[6][175] = 5'b11111;
assign A[6][176] = 5'b00000;
assign A[6][177] = 5'b11111;
assign A[6][178] = 5'b11111;
assign A[6][179] = 5'b11100;
assign A[6][180] = 5'b11100;
assign A[6][181] = 5'b00000;
assign A[6][182] = 5'b11110;
assign A[6][183] = 5'b11100;
assign A[6][184] = 5'b00001;
assign A[6][185] = 5'b00010;
assign A[6][186] = 5'b00000;
assign A[6][187] = 5'b11110;
assign A[6][188] = 5'b11110;
assign A[6][189] = 5'b00001;
assign A[6][190] = 5'b11111;
assign A[6][191] = 5'b00001;
assign A[6][192] = 5'b00000;
assign A[6][193] = 5'b11111;
assign A[6][194] = 5'b11101;
assign A[6][195] = 5'b00001;
assign A[6][196] = 5'b11110;
assign A[6][197] = 5'b11110;
assign A[6][198] = 5'b11110;
assign A[6][199] = 5'b00000;
assign A[6][200] = 5'b00001;
assign A[6][201] = 5'b11111;
assign A[6][202] = 5'b00000;
assign A[6][203] = 5'b11111;
assign A[6][204] = 5'b11111;
assign A[6][205] = 5'b11110;
assign A[6][206] = 5'b00001;
assign A[6][207] = 5'b00010;
assign A[6][208] = 5'b00001;
assign A[6][209] = 5'b00001;
assign A[6][210] = 5'b11111;
assign A[6][211] = 5'b00010;
assign A[6][212] = 5'b00000;
assign A[6][213] = 5'b00010;
assign A[6][214] = 5'b00000;
assign A[6][215] = 5'b11110;
assign A[6][216] = 5'b00000;
assign A[6][217] = 5'b11111;
assign A[6][218] = 5'b11111;
assign A[6][219] = 5'b00000;
assign A[6][220] = 5'b00001;
assign A[6][221] = 5'b11110;
assign A[6][222] = 5'b11101;
assign A[6][223] = 5'b11111;
assign A[6][224] = 5'b00000;
assign A[6][225] = 5'b00001;
assign A[6][226] = 5'b11111;
assign A[6][227] = 5'b11111;
assign A[6][228] = 5'b11111;
assign A[6][229] = 5'b11101;
assign A[6][230] = 5'b00001;
assign A[6][231] = 5'b11101;
assign A[6][232] = 5'b00000;
assign A[6][233] = 5'b11111;
assign A[6][234] = 5'b11101;
assign A[6][235] = 5'b00000;
assign A[6][236] = 5'b00000;
assign A[6][237] = 5'b11110;
assign A[6][238] = 5'b11101;
assign A[6][239] = 5'b11110;
assign A[6][240] = 5'b00001;
assign A[6][241] = 5'b00001;
assign A[6][242] = 5'b00001;
assign A[6][243] = 5'b00001;
assign A[6][244] = 5'b11111;
assign A[6][245] = 5'b00000;
assign A[6][246] = 5'b00011;
assign A[6][247] = 5'b11111;
assign A[6][248] = 5'b00000;
assign A[6][249] = 5'b00000;
assign A[6][250] = 5'b00001;
assign A[6][251] = 5'b00010;
assign A[6][252] = 5'b11110;
assign A[6][253] = 5'b00010;
assign A[6][254] = 5'b11111;
assign A[6][255] = 5'b11101;
assign A[7][0] = 5'b11111;
assign A[7][1] = 5'b11111;
assign A[7][2] = 5'b00000;
assign A[7][3] = 5'b00000;
assign A[7][4] = 5'b11110;
assign A[7][5] = 5'b00000;
assign A[7][6] = 5'b00010;
assign A[7][7] = 5'b00001;
assign A[7][8] = 5'b11110;
assign A[7][9] = 5'b11111;
assign A[7][10] = 5'b00001;
assign A[7][11] = 5'b11111;
assign A[7][12] = 5'b00010;
assign A[7][13] = 5'b11111;
assign A[7][14] = 5'b11111;
assign A[7][15] = 5'b00010;
assign A[7][16] = 5'b00001;
assign A[7][17] = 5'b00001;
assign A[7][18] = 5'b11110;
assign A[7][19] = 5'b00000;
assign A[7][20] = 5'b00000;
assign A[7][21] = 5'b11110;
assign A[7][22] = 5'b11111;
assign A[7][23] = 5'b00001;
assign A[7][24] = 5'b00001;
assign A[7][25] = 5'b00100;
assign A[7][26] = 5'b11101;
assign A[7][27] = 5'b00000;
assign A[7][28] = 5'b00001;
assign A[7][29] = 5'b11101;
assign A[7][30] = 5'b00000;
assign A[7][31] = 5'b00010;
assign A[7][32] = 5'b00000;
assign A[7][33] = 5'b00000;
assign A[7][34] = 5'b00000;
assign A[7][35] = 5'b00001;
assign A[7][36] = 5'b00000;
assign A[7][37] = 5'b00000;
assign A[7][38] = 5'b11110;
assign A[7][39] = 5'b11101;
assign A[7][40] = 5'b11111;
assign A[7][41] = 5'b11110;
assign A[7][42] = 5'b11110;
assign A[7][43] = 5'b11111;
assign A[7][44] = 5'b00001;
assign A[7][45] = 5'b00001;
assign A[7][46] = 5'b11111;
assign A[7][47] = 5'b00001;
assign A[7][48] = 5'b00001;
assign A[7][49] = 5'b11110;
assign A[7][50] = 5'b00010;
assign A[7][51] = 5'b11101;
assign A[7][52] = 5'b00001;
assign A[7][53] = 5'b00000;
assign A[7][54] = 5'b00000;
assign A[7][55] = 5'b00001;
assign A[7][56] = 5'b11111;
assign A[7][57] = 5'b11100;
assign A[7][58] = 5'b11011;
assign A[7][59] = 5'b11110;
assign A[7][60] = 5'b00000;
assign A[7][61] = 5'b00000;
assign A[7][62] = 5'b11101;
assign A[7][63] = 5'b11110;
assign A[7][64] = 5'b11110;
assign A[7][65] = 5'b00010;
assign A[7][66] = 5'b00001;
assign A[7][67] = 5'b11111;
assign A[7][68] = 5'b00001;
assign A[7][69] = 5'b11111;
assign A[7][70] = 5'b11110;
assign A[7][71] = 5'b00001;
assign A[7][72] = 5'b00001;
assign A[7][73] = 5'b11101;
assign A[7][74] = 5'b11011;
assign A[7][75] = 5'b11101;
assign A[7][76] = 5'b11110;
assign A[7][77] = 5'b11101;
assign A[7][78] = 5'b11110;
assign A[7][79] = 5'b00000;
assign A[7][80] = 5'b11111;
assign A[7][81] = 5'b11110;
assign A[7][82] = 5'b11111;
assign A[7][83] = 5'b11110;
assign A[7][84] = 5'b11110;
assign A[7][85] = 5'b00001;
assign A[7][86] = 5'b00101;
assign A[7][87] = 5'b00001;
assign A[7][88] = 5'b00001;
assign A[7][89] = 5'b00000;
assign A[7][90] = 5'b00000;
assign A[7][91] = 5'b00000;
assign A[7][92] = 5'b11111;
assign A[7][93] = 5'b11110;
assign A[7][94] = 5'b11100;
assign A[7][95] = 5'b11101;
assign A[7][96] = 5'b00000;
assign A[7][97] = 5'b11111;
assign A[7][98] = 5'b11110;
assign A[7][99] = 5'b11111;
assign A[7][100] = 5'b00001;
assign A[7][101] = 5'b00001;
assign A[7][102] = 5'b00101;
assign A[7][103] = 5'b11111;
assign A[7][104] = 5'b00001;
assign A[7][105] = 5'b00000;
assign A[7][106] = 5'b00000;
assign A[7][107] = 5'b00010;
assign A[7][108] = 5'b00000;
assign A[7][109] = 5'b11110;
assign A[7][110] = 5'b00000;
assign A[7][111] = 5'b11011;
assign A[7][112] = 5'b00000;
assign A[7][113] = 5'b11111;
assign A[7][114] = 5'b00001;
assign A[7][115] = 5'b00000;
assign A[7][116] = 5'b00000;
assign A[7][117] = 5'b00001;
assign A[7][118] = 5'b00001;
assign A[7][119] = 5'b00000;
assign A[7][120] = 5'b00001;
assign A[7][121] = 5'b11111;
assign A[7][122] = 5'b00000;
assign A[7][123] = 5'b00000;
assign A[7][124] = 5'b00100;
assign A[7][125] = 5'b00000;
assign A[7][126] = 5'b11110;
assign A[7][127] = 5'b11111;
assign A[7][128] = 5'b00010;
assign A[7][129] = 5'b11110;
assign A[7][130] = 5'b00011;
assign A[7][131] = 5'b00000;
assign A[7][132] = 5'b00000;
assign A[7][133] = 5'b00001;
assign A[7][134] = 5'b00001;
assign A[7][135] = 5'b00011;
assign A[7][136] = 5'b00001;
assign A[7][137] = 5'b00000;
assign A[7][138] = 5'b00010;
assign A[7][139] = 5'b00000;
assign A[7][140] = 5'b00000;
assign A[7][141] = 5'b00000;
assign A[7][142] = 5'b11111;
assign A[7][143] = 5'b11111;
assign A[7][144] = 5'b00001;
assign A[7][145] = 5'b00010;
assign A[7][146] = 5'b11101;
assign A[7][147] = 5'b00000;
assign A[7][148] = 5'b00000;
assign A[7][149] = 5'b00001;
assign A[7][150] = 5'b00001;
assign A[7][151] = 5'b00001;
assign A[7][152] = 5'b00001;
assign A[7][153] = 5'b00001;
assign A[7][154] = 5'b00010;
assign A[7][155] = 5'b00000;
assign A[7][156] = 5'b00001;
assign A[7][157] = 5'b00001;
assign A[7][158] = 5'b11111;
assign A[7][159] = 5'b00001;
assign A[7][160] = 5'b00000;
assign A[7][161] = 5'b00001;
assign A[7][162] = 5'b00001;
assign A[7][163] = 5'b00010;
assign A[7][164] = 5'b00000;
assign A[7][165] = 5'b00010;
assign A[7][166] = 5'b00010;
assign A[7][167] = 5'b11111;
assign A[7][168] = 5'b00010;
assign A[7][169] = 5'b00010;
assign A[7][170] = 5'b11111;
assign A[7][171] = 5'b00001;
assign A[7][172] = 5'b00000;
assign A[7][173] = 5'b00011;
assign A[7][174] = 5'b00001;
assign A[7][175] = 5'b00000;
assign A[7][176] = 5'b00001;
assign A[7][177] = 5'b00101;
assign A[7][178] = 5'b00001;
assign A[7][179] = 5'b00001;
assign A[7][180] = 5'b11111;
assign A[7][181] = 5'b11111;
assign A[7][182] = 5'b00000;
assign A[7][183] = 5'b00001;
assign A[7][184] = 5'b00001;
assign A[7][185] = 5'b00001;
assign A[7][186] = 5'b00001;
assign A[7][187] = 5'b00000;
assign A[7][188] = 5'b00010;
assign A[7][189] = 5'b00000;
assign A[7][190] = 5'b00011;
assign A[7][191] = 5'b00001;
assign A[7][192] = 5'b00011;
assign A[7][193] = 5'b00101;
assign A[7][194] = 5'b00001;
assign A[7][195] = 5'b00000;
assign A[7][196] = 5'b00011;
assign A[7][197] = 5'b11111;
assign A[7][198] = 5'b11110;
assign A[7][199] = 5'b00001;
assign A[7][200] = 5'b00000;
assign A[7][201] = 5'b11101;
assign A[7][202] = 5'b00001;
assign A[7][203] = 5'b00010;
assign A[7][204] = 5'b00000;
assign A[7][205] = 5'b00001;
assign A[7][206] = 5'b00001;
assign A[7][207] = 5'b00100;
assign A[7][208] = 5'b00001;
assign A[7][209] = 5'b00000;
assign A[7][210] = 5'b11111;
assign A[7][211] = 5'b11111;
assign A[7][212] = 5'b11111;
assign A[7][213] = 5'b00000;
assign A[7][214] = 5'b11111;
assign A[7][215] = 5'b11110;
assign A[7][216] = 5'b00001;
assign A[7][217] = 5'b00000;
assign A[7][218] = 5'b11101;
assign A[7][219] = 5'b11111;
assign A[7][220] = 5'b00001;
assign A[7][221] = 5'b11011;
assign A[7][222] = 5'b00001;
assign A[7][223] = 5'b00000;
assign A[7][224] = 5'b11110;
assign A[7][225] = 5'b11111;
assign A[7][226] = 5'b11110;
assign A[7][227] = 5'b00010;
assign A[7][228] = 5'b00011;
assign A[7][229] = 5'b00001;
assign A[7][230] = 5'b00000;
assign A[7][231] = 5'b00100;
assign A[7][232] = 5'b00000;
assign A[7][233] = 5'b11111;
assign A[7][234] = 5'b00010;
assign A[7][235] = 5'b00000;
assign A[7][236] = 5'b00000;
assign A[7][237] = 5'b00000;
assign A[7][238] = 5'b11101;
assign A[7][239] = 5'b11101;
assign A[7][240] = 5'b11110;
assign A[7][241] = 5'b00010;
assign A[7][242] = 5'b00000;
assign A[7][243] = 5'b00010;
assign A[7][244] = 5'b00001;
assign A[7][245] = 5'b00000;
assign A[7][246] = 5'b00001;
assign A[7][247] = 5'b00001;
assign A[7][248] = 5'b00001;
assign A[7][249] = 5'b11110;
assign A[7][250] = 5'b00010;
assign A[7][251] = 5'b00010;
assign A[7][252] = 5'b00000;
assign A[7][253] = 5'b11111;
assign A[7][254] = 5'b11101;
assign A[7][255] = 5'b11101;
assign A[8][0] = 5'b00011;
assign A[8][1] = 5'b00001;
assign A[8][2] = 5'b00010;
assign A[8][3] = 5'b11111;
assign A[8][4] = 5'b00001;
assign A[8][5] = 5'b00000;
assign A[8][6] = 5'b00000;
assign A[8][7] = 5'b11110;
assign A[8][8] = 5'b00001;
assign A[8][9] = 5'b00001;
assign A[8][10] = 5'b11110;
assign A[8][11] = 5'b00001;
assign A[8][12] = 5'b00000;
assign A[8][13] = 5'b00010;
assign A[8][14] = 5'b11111;
assign A[8][15] = 5'b00000;
assign A[8][16] = 5'b11111;
assign A[8][17] = 5'b00000;
assign A[8][18] = 5'b00000;
assign A[8][19] = 5'b00010;
assign A[8][20] = 5'b00010;
assign A[8][21] = 5'b11110;
assign A[8][22] = 5'b11110;
assign A[8][23] = 5'b11111;
assign A[8][24] = 5'b00001;
assign A[8][25] = 5'b11111;
assign A[8][26] = 5'b00000;
assign A[8][27] = 5'b11111;
assign A[8][28] = 5'b00010;
assign A[8][29] = 5'b11110;
assign A[8][30] = 5'b11101;
assign A[8][31] = 5'b00000;
assign A[8][32] = 5'b00010;
assign A[8][33] = 5'b00000;
assign A[8][34] = 5'b11111;
assign A[8][35] = 5'b00000;
assign A[8][36] = 5'b00001;
assign A[8][37] = 5'b00001;
assign A[8][38] = 5'b00001;
assign A[8][39] = 5'b00001;
assign A[8][40] = 5'b00001;
assign A[8][41] = 5'b11111;
assign A[8][42] = 5'b11111;
assign A[8][43] = 5'b00000;
assign A[8][44] = 5'b11101;
assign A[8][45] = 5'b11101;
assign A[8][46] = 5'b00001;
assign A[8][47] = 5'b11111;
assign A[8][48] = 5'b00011;
assign A[8][49] = 5'b00010;
assign A[8][50] = 5'b00000;
assign A[8][51] = 5'b00010;
assign A[8][52] = 5'b00000;
assign A[8][53] = 5'b00010;
assign A[8][54] = 5'b00001;
assign A[8][55] = 5'b11101;
assign A[8][56] = 5'b11111;
assign A[8][57] = 5'b11110;
assign A[8][58] = 5'b11111;
assign A[8][59] = 5'b11110;
assign A[8][60] = 5'b00000;
assign A[8][61] = 5'b11111;
assign A[8][62] = 5'b11110;
assign A[8][63] = 5'b11110;
assign A[8][64] = 5'b11101;
assign A[8][65] = 5'b00011;
assign A[8][66] = 5'b00000;
assign A[8][67] = 5'b11111;
assign A[8][68] = 5'b00001;
assign A[8][69] = 5'b00001;
assign A[8][70] = 5'b00000;
assign A[8][71] = 5'b11101;
assign A[8][72] = 5'b11100;
assign A[8][73] = 5'b11100;
assign A[8][74] = 5'b00000;
assign A[8][75] = 5'b11111;
assign A[8][76] = 5'b11101;
assign A[8][77] = 5'b11110;
assign A[8][78] = 5'b11110;
assign A[8][79] = 5'b00001;
assign A[8][80] = 5'b11110;
assign A[8][81] = 5'b11110;
assign A[8][82] = 5'b11110;
assign A[8][83] = 5'b11110;
assign A[8][84] = 5'b11101;
assign A[8][85] = 5'b00000;
assign A[8][86] = 5'b11110;
assign A[8][87] = 5'b00000;
assign A[8][88] = 5'b00001;
assign A[8][89] = 5'b11111;
assign A[8][90] = 5'b00001;
assign A[8][91] = 5'b11101;
assign A[8][92] = 5'b11110;
assign A[8][93] = 5'b00010;
assign A[8][94] = 5'b11011;
assign A[8][95] = 5'b00001;
assign A[8][96] = 5'b11110;
assign A[8][97] = 5'b11110;
assign A[8][98] = 5'b11111;
assign A[8][99] = 5'b00000;
assign A[8][100] = 5'b11101;
assign A[8][101] = 5'b00000;
assign A[8][102] = 5'b00000;
assign A[8][103] = 5'b11111;
assign A[8][104] = 5'b11110;
assign A[8][105] = 5'b11111;
assign A[8][106] = 5'b11111;
assign A[8][107] = 5'b00000;
assign A[8][108] = 5'b00000;
assign A[8][109] = 5'b00001;
assign A[8][110] = 5'b11111;
assign A[8][111] = 5'b11101;
assign A[8][112] = 5'b00001;
assign A[8][113] = 5'b11110;
assign A[8][114] = 5'b11110;
assign A[8][115] = 5'b00001;
assign A[8][116] = 5'b00000;
assign A[8][117] = 5'b00001;
assign A[8][118] = 5'b11110;
assign A[8][119] = 5'b00001;
assign A[8][120] = 5'b11110;
assign A[8][121] = 5'b11111;
assign A[8][122] = 5'b00001;
assign A[8][123] = 5'b00000;
assign A[8][124] = 5'b00001;
assign A[8][125] = 5'b11110;
assign A[8][126] = 5'b11111;
assign A[8][127] = 5'b00000;
assign A[8][128] = 5'b00010;
assign A[8][129] = 5'b00001;
assign A[8][130] = 5'b00001;
assign A[8][131] = 5'b00011;
assign A[8][132] = 5'b11110;
assign A[8][133] = 5'b00000;
assign A[8][134] = 5'b00001;
assign A[8][135] = 5'b00000;
assign A[8][136] = 5'b00001;
assign A[8][137] = 5'b11101;
assign A[8][138] = 5'b00001;
assign A[8][139] = 5'b11111;
assign A[8][140] = 5'b11110;
assign A[8][141] = 5'b00001;
assign A[8][142] = 5'b11110;
assign A[8][143] = 5'b00010;
assign A[8][144] = 5'b00001;
assign A[8][145] = 5'b00010;
assign A[8][146] = 5'b00001;
assign A[8][147] = 5'b00010;
assign A[8][148] = 5'b00011;
assign A[8][149] = 5'b00001;
assign A[8][150] = 5'b11110;
assign A[8][151] = 5'b11111;
assign A[8][152] = 5'b00010;
assign A[8][153] = 5'b00000;
assign A[8][154] = 5'b00010;
assign A[8][155] = 5'b00000;
assign A[8][156] = 5'b00001;
assign A[8][157] = 5'b00001;
assign A[8][158] = 5'b11100;
assign A[8][159] = 5'b11111;
assign A[8][160] = 5'b00010;
assign A[8][161] = 5'b00100;
assign A[8][162] = 5'b00011;
assign A[8][163] = 5'b00001;
assign A[8][164] = 5'b00011;
assign A[8][165] = 5'b00001;
assign A[8][166] = 5'b00100;
assign A[8][167] = 5'b00000;
assign A[8][168] = 5'b00001;
assign A[8][169] = 5'b00010;
assign A[8][170] = 5'b11111;
assign A[8][171] = 5'b11111;
assign A[8][172] = 5'b11111;
assign A[8][173] = 5'b11110;
assign A[8][174] = 5'b00000;
assign A[8][175] = 5'b00001;
assign A[8][176] = 5'b11111;
assign A[8][177] = 5'b00100;
assign A[8][178] = 5'b00001;
assign A[8][179] = 5'b00010;
assign A[8][180] = 5'b00011;
assign A[8][181] = 5'b00011;
assign A[8][182] = 5'b00011;
assign A[8][183] = 5'b00000;
assign A[8][184] = 5'b11110;
assign A[8][185] = 5'b00000;
assign A[8][186] = 5'b11111;
assign A[8][187] = 5'b11110;
assign A[8][188] = 5'b11100;
assign A[8][189] = 5'b00000;
assign A[8][190] = 5'b11110;
assign A[8][191] = 5'b11101;
assign A[8][192] = 5'b00001;
assign A[8][193] = 5'b00100;
assign A[8][194] = 5'b00000;
assign A[8][195] = 5'b00011;
assign A[8][196] = 5'b00001;
assign A[8][197] = 5'b00001;
assign A[8][198] = 5'b00011;
assign A[8][199] = 5'b11111;
assign A[8][200] = 5'b00010;
assign A[8][201] = 5'b00001;
assign A[8][202] = 5'b00000;
assign A[8][203] = 5'b11111;
assign A[8][204] = 5'b00010;
assign A[8][205] = 5'b11110;
assign A[8][206] = 5'b11111;
assign A[8][207] = 5'b00001;
assign A[8][208] = 5'b00100;
assign A[8][209] = 5'b00001;
assign A[8][210] = 5'b11111;
assign A[8][211] = 5'b00001;
assign A[8][212] = 5'b00000;
assign A[8][213] = 5'b00000;
assign A[8][214] = 5'b00000;
assign A[8][215] = 5'b11111;
assign A[8][216] = 5'b00001;
assign A[8][217] = 5'b00000;
assign A[8][218] = 5'b00001;
assign A[8][219] = 5'b00000;
assign A[8][220] = 5'b11111;
assign A[8][221] = 5'b11111;
assign A[8][222] = 5'b11111;
assign A[8][223] = 5'b11101;
assign A[8][224] = 5'b00001;
assign A[8][225] = 5'b11111;
assign A[8][226] = 5'b00001;
assign A[8][227] = 5'b00001;
assign A[8][228] = 5'b11111;
assign A[8][229] = 5'b00001;
assign A[8][230] = 5'b00011;
assign A[8][231] = 5'b11110;
assign A[8][232] = 5'b11111;
assign A[8][233] = 5'b00001;
assign A[8][234] = 5'b00001;
assign A[8][235] = 5'b11110;
assign A[8][236] = 5'b00001;
assign A[8][237] = 5'b11111;
assign A[8][238] = 5'b11110;
assign A[8][239] = 5'b00010;
assign A[8][240] = 5'b11101;
assign A[8][241] = 5'b00001;
assign A[8][242] = 5'b00000;
assign A[8][243] = 5'b11110;
assign A[8][244] = 5'b00000;
assign A[8][245] = 5'b00000;
assign A[8][246] = 5'b00000;
assign A[8][247] = 5'b00010;
assign A[8][248] = 5'b00000;
assign A[8][249] = 5'b00000;
assign A[8][250] = 5'b00010;
assign A[8][251] = 5'b00001;
assign A[8][252] = 5'b11111;
assign A[8][253] = 5'b00100;
assign A[8][254] = 5'b00000;
assign A[8][255] = 5'b00000;
assign A[9][0] = 5'b00100;
assign A[9][1] = 5'b00000;
assign A[9][2] = 5'b00010;
assign A[9][3] = 5'b00011;
assign A[9][4] = 5'b11111;
assign A[9][5] = 5'b00010;
assign A[9][6] = 5'b11110;
assign A[9][7] = 5'b00101;
assign A[9][8] = 5'b00001;
assign A[9][9] = 5'b00000;
assign A[9][10] = 5'b00001;
assign A[9][11] = 5'b11111;
assign A[9][12] = 5'b00000;
assign A[9][13] = 5'b00000;
assign A[9][14] = 5'b11111;
assign A[9][15] = 5'b00000;
assign A[9][16] = 5'b00010;
assign A[9][17] = 5'b00010;
assign A[9][18] = 5'b11110;
assign A[9][19] = 5'b00010;
assign A[9][20] = 5'b00000;
assign A[9][21] = 5'b00001;
assign A[9][22] = 5'b00001;
assign A[9][23] = 5'b00000;
assign A[9][24] = 5'b00000;
assign A[9][25] = 5'b11110;
assign A[9][26] = 5'b11111;
assign A[9][27] = 5'b00000;
assign A[9][28] = 5'b00000;
assign A[9][29] = 5'b11110;
assign A[9][30] = 5'b00100;
assign A[9][31] = 5'b00000;
assign A[9][32] = 5'b11111;
assign A[9][33] = 5'b00010;
assign A[9][34] = 5'b00001;
assign A[9][35] = 5'b00000;
assign A[9][36] = 5'b00001;
assign A[9][37] = 5'b00000;
assign A[9][38] = 5'b00010;
assign A[9][39] = 5'b00010;
assign A[9][40] = 5'b00000;
assign A[9][41] = 5'b00000;
assign A[9][42] = 5'b11111;
assign A[9][43] = 5'b00010;
assign A[9][44] = 5'b00000;
assign A[9][45] = 5'b00010;
assign A[9][46] = 5'b00010;
assign A[9][47] = 5'b00010;
assign A[9][48] = 5'b11111;
assign A[9][49] = 5'b11110;
assign A[9][50] = 5'b00010;
assign A[9][51] = 5'b00000;
assign A[9][52] = 5'b11110;
assign A[9][53] = 5'b00000;
assign A[9][54] = 5'b11111;
assign A[9][55] = 5'b00001;
assign A[9][56] = 5'b00010;
assign A[9][57] = 5'b00010;
assign A[9][58] = 5'b11111;
assign A[9][59] = 5'b00000;
assign A[9][60] = 5'b00010;
assign A[9][61] = 5'b00001;
assign A[9][62] = 5'b00010;
assign A[9][63] = 5'b00000;
assign A[9][64] = 5'b11111;
assign A[9][65] = 5'b11101;
assign A[9][66] = 5'b11110;
assign A[9][67] = 5'b00000;
assign A[9][68] = 5'b11111;
assign A[9][69] = 5'b00001;
assign A[9][70] = 5'b11110;
assign A[9][71] = 5'b00010;
assign A[9][72] = 5'b00011;
assign A[9][73] = 5'b00000;
assign A[9][74] = 5'b00011;
assign A[9][75] = 5'b00001;
assign A[9][76] = 5'b00011;
assign A[9][77] = 5'b00010;
assign A[9][78] = 5'b00000;
assign A[9][79] = 5'b00001;
assign A[9][80] = 5'b11110;
assign A[9][81] = 5'b11110;
assign A[9][82] = 5'b00011;
assign A[9][83] = 5'b00000;
assign A[9][84] = 5'b11110;
assign A[9][85] = 5'b00000;
assign A[9][86] = 5'b00010;
assign A[9][87] = 5'b00001;
assign A[9][88] = 5'b00001;
assign A[9][89] = 5'b00000;
assign A[9][90] = 5'b00000;
assign A[9][91] = 5'b11111;
assign A[9][92] = 5'b00000;
assign A[9][93] = 5'b11110;
assign A[9][94] = 5'b11110;
assign A[9][95] = 5'b00001;
assign A[9][96] = 5'b00000;
assign A[9][97] = 5'b11110;
assign A[9][98] = 5'b11101;
assign A[9][99] = 5'b00000;
assign A[9][100] = 5'b00010;
assign A[9][101] = 5'b00010;
assign A[9][102] = 5'b00001;
assign A[9][103] = 5'b00001;
assign A[9][104] = 5'b00000;
assign A[9][105] = 5'b00001;
assign A[9][106] = 5'b00001;
assign A[9][107] = 5'b00000;
assign A[9][108] = 5'b00010;
assign A[9][109] = 5'b00000;
assign A[9][110] = 5'b11110;
assign A[9][111] = 5'b00000;
assign A[9][112] = 5'b00000;
assign A[9][113] = 5'b00010;
assign A[9][114] = 5'b00001;
assign A[9][115] = 5'b00000;
assign A[9][116] = 5'b00001;
assign A[9][117] = 5'b00000;
assign A[9][118] = 5'b00001;
assign A[9][119] = 5'b00001;
assign A[9][120] = 5'b00010;
assign A[9][121] = 5'b00001;
assign A[9][122] = 5'b00000;
assign A[9][123] = 5'b00010;
assign A[9][124] = 5'b00011;
assign A[9][125] = 5'b00000;
assign A[9][126] = 5'b11110;
assign A[9][127] = 5'b00001;
assign A[9][128] = 5'b11110;
assign A[9][129] = 5'b11110;
assign A[9][130] = 5'b00001;
assign A[9][131] = 5'b00001;
assign A[9][132] = 5'b00000;
assign A[9][133] = 5'b11111;
assign A[9][134] = 5'b00010;
assign A[9][135] = 5'b11111;
assign A[9][136] = 5'b00000;
assign A[9][137] = 5'b00010;
assign A[9][138] = 5'b00001;
assign A[9][139] = 5'b00001;
assign A[9][140] = 5'b11111;
assign A[9][141] = 5'b00001;
assign A[9][142] = 5'b00000;
assign A[9][143] = 5'b00011;
assign A[9][144] = 5'b00000;
assign A[9][145] = 5'b00000;
assign A[9][146] = 5'b11101;
assign A[9][147] = 5'b00000;
assign A[9][148] = 5'b11110;
assign A[9][149] = 5'b00010;
assign A[9][150] = 5'b00001;
assign A[9][151] = 5'b00001;
assign A[9][152] = 5'b11111;
assign A[9][153] = 5'b00010;
assign A[9][154] = 5'b00001;
assign A[9][155] = 5'b00001;
assign A[9][156] = 5'b00011;
assign A[9][157] = 5'b11111;
assign A[9][158] = 5'b00000;
assign A[9][159] = 5'b00011;
assign A[9][160] = 5'b00000;
assign A[9][161] = 5'b11111;
assign A[9][162] = 5'b00000;
assign A[9][163] = 5'b11101;
assign A[9][164] = 5'b11111;
assign A[9][165] = 5'b00000;
assign A[9][166] = 5'b00001;
assign A[9][167] = 5'b00000;
assign A[9][168] = 5'b00010;
assign A[9][169] = 5'b11110;
assign A[9][170] = 5'b00001;
assign A[9][171] = 5'b00000;
assign A[9][172] = 5'b00001;
assign A[9][173] = 5'b00010;
assign A[9][174] = 5'b00001;
assign A[9][175] = 5'b00010;
assign A[9][176] = 5'b11101;
assign A[9][177] = 5'b11110;
assign A[9][178] = 5'b11111;
assign A[9][179] = 5'b11111;
assign A[9][180] = 5'b00001;
assign A[9][181] = 5'b11110;
assign A[9][182] = 5'b11100;
assign A[9][183] = 5'b00010;
assign A[9][184] = 5'b00010;
assign A[9][185] = 5'b00001;
assign A[9][186] = 5'b00000;
assign A[9][187] = 5'b11110;
assign A[9][188] = 5'b11111;
assign A[9][189] = 5'b00000;
assign A[9][190] = 5'b11111;
assign A[9][191] = 5'b00001;
assign A[9][192] = 5'b11110;
assign A[9][193] = 5'b11110;
assign A[9][194] = 5'b00000;
assign A[9][195] = 5'b11111;
assign A[9][196] = 5'b11111;
assign A[9][197] = 5'b00011;
assign A[9][198] = 5'b11111;
assign A[9][199] = 5'b11110;
assign A[9][200] = 5'b11110;
assign A[9][201] = 5'b11111;
assign A[9][202] = 5'b11110;
assign A[9][203] = 5'b00001;
assign A[9][204] = 5'b11111;
assign A[9][205] = 5'b00001;
assign A[9][206] = 5'b11111;
assign A[9][207] = 5'b00000;
assign A[9][208] = 5'b11111;
assign A[9][209] = 5'b00011;
assign A[9][210] = 5'b11110;
assign A[9][211] = 5'b11110;
assign A[9][212] = 5'b11110;
assign A[9][213] = 5'b11110;
assign A[9][214] = 5'b11110;
assign A[9][215] = 5'b11110;
assign A[9][216] = 5'b11111;
assign A[9][217] = 5'b11101;
assign A[9][218] = 5'b11111;
assign A[9][219] = 5'b00010;
assign A[9][220] = 5'b11111;
assign A[9][221] = 5'b11101;
assign A[9][222] = 5'b00001;
assign A[9][223] = 5'b11111;
assign A[9][224] = 5'b00001;
assign A[9][225] = 5'b11111;
assign A[9][226] = 5'b11101;
assign A[9][227] = 5'b11101;
assign A[9][228] = 5'b11111;
assign A[9][229] = 5'b11111;
assign A[9][230] = 5'b11101;
assign A[9][231] = 5'b11111;
assign A[9][232] = 5'b11110;
assign A[9][233] = 5'b11110;
assign A[9][234] = 5'b11100;
assign A[9][235] = 5'b11111;
assign A[9][236] = 5'b00001;
assign A[9][237] = 5'b00000;
assign A[9][238] = 5'b11110;
assign A[9][239] = 5'b11111;
assign A[9][240] = 5'b11111;
assign A[9][241] = 5'b11101;
assign A[9][242] = 5'b00010;
assign A[9][243] = 5'b00000;
assign A[9][244] = 5'b11110;
assign A[9][245] = 5'b11011;
assign A[9][246] = 5'b11111;
assign A[9][247] = 5'b11111;
assign A[9][248] = 5'b11111;
assign A[9][249] = 5'b00000;
assign A[9][250] = 5'b11110;
assign A[9][251] = 5'b11111;
assign A[9][252] = 5'b11111;
assign A[9][253] = 5'b11011;
assign A[9][254] = 5'b11101;
assign A[9][255] = 5'b00010;
assign A[10][0] = 5'b11110;
assign A[10][1] = 5'b00001;
assign A[10][2] = 5'b11111;
assign A[10][3] = 5'b11111;
assign A[10][4] = 5'b11110;
assign A[10][5] = 5'b11101;
assign A[10][6] = 5'b11111;
assign A[10][7] = 5'b00001;
assign A[10][8] = 5'b11110;
assign A[10][9] = 5'b00000;
assign A[10][10] = 5'b11111;
assign A[10][11] = 5'b00000;
assign A[10][12] = 5'b11111;
assign A[10][13] = 5'b00000;
assign A[10][14] = 5'b00000;
assign A[10][15] = 5'b00001;
assign A[10][16] = 5'b11111;
assign A[10][17] = 5'b00001;
assign A[10][18] = 5'b11110;
assign A[10][19] = 5'b11111;
assign A[10][20] = 5'b00010;
assign A[10][21] = 5'b00001;
assign A[10][22] = 5'b00000;
assign A[10][23] = 5'b11111;
assign A[10][24] = 5'b11111;
assign A[10][25] = 5'b11110;
assign A[10][26] = 5'b00000;
assign A[10][27] = 5'b11111;
assign A[10][28] = 5'b00001;
assign A[10][29] = 5'b11111;
assign A[10][30] = 5'b00001;
assign A[10][31] = 5'b00000;
assign A[10][32] = 5'b11110;
assign A[10][33] = 5'b00001;
assign A[10][34] = 5'b00000;
assign A[10][35] = 5'b11110;
assign A[10][36] = 5'b00000;
assign A[10][37] = 5'b00010;
assign A[10][38] = 5'b11110;
assign A[10][39] = 5'b11110;
assign A[10][40] = 5'b00001;
assign A[10][41] = 5'b00001;
assign A[10][42] = 5'b11110;
assign A[10][43] = 5'b11111;
assign A[10][44] = 5'b11111;
assign A[10][45] = 5'b00000;
assign A[10][46] = 5'b11111;
assign A[10][47] = 5'b00000;
assign A[10][48] = 5'b11111;
assign A[10][49] = 5'b11111;
assign A[10][50] = 5'b00000;
assign A[10][51] = 5'b00010;
assign A[10][52] = 5'b00010;
assign A[10][53] = 5'b00010;
assign A[10][54] = 5'b00000;
assign A[10][55] = 5'b11110;
assign A[10][56] = 5'b00001;
assign A[10][57] = 5'b11101;
assign A[10][58] = 5'b00000;
assign A[10][59] = 5'b00000;
assign A[10][60] = 5'b00001;
assign A[10][61] = 5'b11111;
assign A[10][62] = 5'b00000;
assign A[10][63] = 5'b11110;
assign A[10][64] = 5'b00000;
assign A[10][65] = 5'b00001;
assign A[10][66] = 5'b00001;
assign A[10][67] = 5'b11111;
assign A[10][68] = 5'b00000;
assign A[10][69] = 5'b00000;
assign A[10][70] = 5'b00001;
assign A[10][71] = 5'b00000;
assign A[10][72] = 5'b11111;
assign A[10][73] = 5'b11110;
assign A[10][74] = 5'b00000;
assign A[10][75] = 5'b00010;
assign A[10][76] = 5'b11111;
assign A[10][77] = 5'b00000;
assign A[10][78] = 5'b00010;
assign A[10][79] = 5'b00001;
assign A[10][80] = 5'b00001;
assign A[10][81] = 5'b00000;
assign A[10][82] = 5'b00001;
assign A[10][83] = 5'b11111;
assign A[10][84] = 5'b11111;
assign A[10][85] = 5'b11110;
assign A[10][86] = 5'b00001;
assign A[10][87] = 5'b00000;
assign A[10][88] = 5'b00000;
assign A[10][89] = 5'b00000;
assign A[10][90] = 5'b00000;
assign A[10][91] = 5'b00001;
assign A[10][92] = 5'b11111;
assign A[10][93] = 5'b00000;
assign A[10][94] = 5'b00001;
assign A[10][95] = 5'b00001;
assign A[10][96] = 5'b00010;
assign A[10][97] = 5'b11111;
assign A[10][98] = 5'b00001;
assign A[10][99] = 5'b00000;
assign A[10][100] = 5'b00000;
assign A[10][101] = 5'b00011;
assign A[10][102] = 5'b00011;
assign A[10][103] = 5'b11111;
assign A[10][104] = 5'b00000;
assign A[10][105] = 5'b00000;
assign A[10][106] = 5'b11110;
assign A[10][107] = 5'b11101;
assign A[10][108] = 5'b11111;
assign A[10][109] = 5'b11111;
assign A[10][110] = 5'b11101;
assign A[10][111] = 5'b00000;
assign A[10][112] = 5'b11110;
assign A[10][113] = 5'b00000;
assign A[10][114] = 5'b00001;
assign A[10][115] = 5'b11101;
assign A[10][116] = 5'b00001;
assign A[10][117] = 5'b11111;
assign A[10][118] = 5'b11111;
assign A[10][119] = 5'b11111;
assign A[10][120] = 5'b00001;
assign A[10][121] = 5'b11111;
assign A[10][122] = 5'b11101;
assign A[10][123] = 5'b11111;
assign A[10][124] = 5'b00010;
assign A[10][125] = 5'b00001;
assign A[10][126] = 5'b00001;
assign A[10][127] = 5'b00001;
assign A[10][128] = 5'b00001;
assign A[10][129] = 5'b00000;
assign A[10][130] = 5'b00000;
assign A[10][131] = 5'b00001;
assign A[10][132] = 5'b00000;
assign A[10][133] = 5'b00001;
assign A[10][134] = 5'b00001;
assign A[10][135] = 5'b11111;
assign A[10][136] = 5'b11110;
assign A[10][137] = 5'b00000;
assign A[10][138] = 5'b00000;
assign A[10][139] = 5'b00010;
assign A[10][140] = 5'b11110;
assign A[10][141] = 5'b00000;
assign A[10][142] = 5'b00001;
assign A[10][143] = 5'b00000;
assign A[10][144] = 5'b11111;
assign A[10][145] = 5'b11101;
assign A[10][146] = 5'b11111;
assign A[10][147] = 5'b11111;
assign A[10][148] = 5'b00000;
assign A[10][149] = 5'b11111;
assign A[10][150] = 5'b11111;
assign A[10][151] = 5'b00001;
assign A[10][152] = 5'b00010;
assign A[10][153] = 5'b00000;
assign A[10][154] = 5'b00000;
assign A[10][155] = 5'b00001;
assign A[10][156] = 5'b00000;
assign A[10][157] = 5'b00010;
assign A[10][158] = 5'b00000;
assign A[10][159] = 5'b00010;
assign A[10][160] = 5'b00000;
assign A[10][161] = 5'b00000;
assign A[10][162] = 5'b00010;
assign A[10][163] = 5'b00011;
assign A[10][164] = 5'b00000;
assign A[10][165] = 5'b11111;
assign A[10][166] = 5'b00010;
assign A[10][167] = 5'b00001;
assign A[10][168] = 5'b11101;
assign A[10][169] = 5'b00000;
assign A[10][170] = 5'b11111;
assign A[10][171] = 5'b00001;
assign A[10][172] = 5'b11110;
assign A[10][173] = 5'b00000;
assign A[10][174] = 5'b00000;
assign A[10][175] = 5'b11111;
assign A[10][176] = 5'b00000;
assign A[10][177] = 5'b00001;
assign A[10][178] = 5'b11111;
assign A[10][179] = 5'b00010;
assign A[10][180] = 5'b11111;
assign A[10][181] = 5'b11110;
assign A[10][182] = 5'b11111;
assign A[10][183] = 5'b11111;
assign A[10][184] = 5'b00000;
assign A[10][185] = 5'b00000;
assign A[10][186] = 5'b11101;
assign A[10][187] = 5'b11110;
assign A[10][188] = 5'b00001;
assign A[10][189] = 5'b00001;
assign A[10][190] = 5'b00001;
assign A[10][191] = 5'b00000;
assign A[10][192] = 5'b00000;
assign A[10][193] = 5'b00001;
assign A[10][194] = 5'b11111;
assign A[10][195] = 5'b00001;
assign A[10][196] = 5'b11110;
assign A[10][197] = 5'b11110;
assign A[10][198] = 5'b00001;
assign A[10][199] = 5'b00000;
assign A[10][200] = 5'b11111;
assign A[10][201] = 5'b00000;
assign A[10][202] = 5'b11111;
assign A[10][203] = 5'b00001;
assign A[10][204] = 5'b00001;
assign A[10][205] = 5'b00000;
assign A[10][206] = 5'b00001;
assign A[10][207] = 5'b00001;
assign A[10][208] = 5'b00001;
assign A[10][209] = 5'b11110;
assign A[10][210] = 5'b11111;
assign A[10][211] = 5'b11111;
assign A[10][212] = 5'b00010;
assign A[10][213] = 5'b11111;
assign A[10][214] = 5'b00000;
assign A[10][215] = 5'b00010;
assign A[10][216] = 5'b11110;
assign A[10][217] = 5'b00000;
assign A[10][218] = 5'b00000;
assign A[10][219] = 5'b00010;
assign A[10][220] = 5'b00011;
assign A[10][221] = 5'b11111;
assign A[10][222] = 5'b00000;
assign A[10][223] = 5'b00010;
assign A[10][224] = 5'b00001;
assign A[10][225] = 5'b00000;
assign A[10][226] = 5'b00010;
assign A[10][227] = 5'b11111;
assign A[10][228] = 5'b00010;
assign A[10][229] = 5'b11111;
assign A[10][230] = 5'b00001;
assign A[10][231] = 5'b11111;
assign A[10][232] = 5'b11110;
assign A[10][233] = 5'b11110;
assign A[10][234] = 5'b00000;
assign A[10][235] = 5'b00000;
assign A[10][236] = 5'b11101;
assign A[10][237] = 5'b00000;
assign A[10][238] = 5'b00000;
assign A[10][239] = 5'b11111;
assign A[10][240] = 5'b11111;
assign A[10][241] = 5'b00001;
assign A[10][242] = 5'b00001;
assign A[10][243] = 5'b00001;
assign A[10][244] = 5'b11111;
assign A[10][245] = 5'b00000;
assign A[10][246] = 5'b11111;
assign A[10][247] = 5'b00001;
assign A[10][248] = 5'b11110;
assign A[10][249] = 5'b00000;
assign A[10][250] = 5'b11111;
assign A[10][251] = 5'b11111;
assign A[10][252] = 5'b00001;
assign A[10][253] = 5'b11111;
assign A[10][254] = 5'b00000;
assign A[10][255] = 5'b00000;
assign A[11][0] = 5'b00100;
assign A[11][1] = 5'b11110;
assign A[11][2] = 5'b11111;
assign A[11][3] = 5'b00000;
assign A[11][4] = 5'b11111;
assign A[11][5] = 5'b11101;
assign A[11][6] = 5'b00000;
assign A[11][7] = 5'b00001;
assign A[11][8] = 5'b11011;
assign A[11][9] = 5'b11110;
assign A[11][10] = 5'b00000;
assign A[11][11] = 5'b11101;
assign A[11][12] = 5'b11110;
assign A[11][13] = 5'b00001;
assign A[11][14] = 5'b11110;
assign A[11][15] = 5'b00001;
assign A[11][16] = 5'b11101;
assign A[11][17] = 5'b00000;
assign A[11][18] = 5'b11111;
assign A[11][19] = 5'b00000;
assign A[11][20] = 5'b11111;
assign A[11][21] = 5'b11111;
assign A[11][22] = 5'b11011;
assign A[11][23] = 5'b11111;
assign A[11][24] = 5'b11101;
assign A[11][25] = 5'b11111;
assign A[11][26] = 5'b00000;
assign A[11][27] = 5'b00010;
assign A[11][28] = 5'b00000;
assign A[11][29] = 5'b11111;
assign A[11][30] = 5'b00010;
assign A[11][31] = 5'b11111;
assign A[11][32] = 5'b11110;
assign A[11][33] = 5'b11111;
assign A[11][34] = 5'b00001;
assign A[11][35] = 5'b11111;
assign A[11][36] = 5'b11111;
assign A[11][37] = 5'b00010;
assign A[11][38] = 5'b00000;
assign A[11][39] = 5'b00000;
assign A[11][40] = 5'b11110;
assign A[11][41] = 5'b11110;
assign A[11][42] = 5'b00000;
assign A[11][43] = 5'b00000;
assign A[11][44] = 5'b00010;
assign A[11][45] = 5'b00001;
assign A[11][46] = 5'b11101;
assign A[11][47] = 5'b00000;
assign A[11][48] = 5'b00000;
assign A[11][49] = 5'b11111;
assign A[11][50] = 5'b11101;
assign A[11][51] = 5'b00000;
assign A[11][52] = 5'b00001;
assign A[11][53] = 5'b00000;
assign A[11][54] = 5'b00000;
assign A[11][55] = 5'b11110;
assign A[11][56] = 5'b00010;
assign A[11][57] = 5'b00001;
assign A[11][58] = 5'b00001;
assign A[11][59] = 5'b11111;
assign A[11][60] = 5'b11011;
assign A[11][61] = 5'b11111;
assign A[11][62] = 5'b11110;
assign A[11][63] = 5'b11011;
assign A[11][64] = 5'b00000;
assign A[11][65] = 5'b11110;
assign A[11][66] = 5'b11111;
assign A[11][67] = 5'b00000;
assign A[11][68] = 5'b00010;
assign A[11][69] = 5'b00010;
assign A[11][70] = 5'b00001;
assign A[11][71] = 5'b11101;
assign A[11][72] = 5'b00000;
assign A[11][73] = 5'b00100;
assign A[11][74] = 5'b11110;
assign A[11][75] = 5'b11110;
assign A[11][76] = 5'b11101;
assign A[11][77] = 5'b11110;
assign A[11][78] = 5'b11111;
assign A[11][79] = 5'b11110;
assign A[11][80] = 5'b00001;
assign A[11][81] = 5'b00010;
assign A[11][82] = 5'b00000;
assign A[11][83] = 5'b11111;
assign A[11][84] = 5'b00001;
assign A[11][85] = 5'b11110;
assign A[11][86] = 5'b11111;
assign A[11][87] = 5'b00000;
assign A[11][88] = 5'b11111;
assign A[11][89] = 5'b11100;
assign A[11][90] = 5'b11111;
assign A[11][91] = 5'b11101;
assign A[11][92] = 5'b11100;
assign A[11][93] = 5'b00000;
assign A[11][94] = 5'b11101;
assign A[11][95] = 5'b00000;
assign A[11][96] = 5'b00010;
assign A[11][97] = 5'b00010;
assign A[11][98] = 5'b11110;
assign A[11][99] = 5'b11111;
assign A[11][100] = 5'b00011;
assign A[11][101] = 5'b11101;
assign A[11][102] = 5'b11110;
assign A[11][103] = 5'b11111;
assign A[11][104] = 5'b11111;
assign A[11][105] = 5'b11111;
assign A[11][106] = 5'b00000;
assign A[11][107] = 5'b11101;
assign A[11][108] = 5'b00010;
assign A[11][109] = 5'b00000;
assign A[11][110] = 5'b11110;
assign A[11][111] = 5'b00000;
assign A[11][112] = 5'b00001;
assign A[11][113] = 5'b00000;
assign A[11][114] = 5'b00001;
assign A[11][115] = 5'b00010;
assign A[11][116] = 5'b00001;
assign A[11][117] = 5'b00001;
assign A[11][118] = 5'b11111;
assign A[11][119] = 5'b00000;
assign A[11][120] = 5'b00001;
assign A[11][121] = 5'b11111;
assign A[11][122] = 5'b00001;
assign A[11][123] = 5'b11111;
assign A[11][124] = 5'b00100;
assign A[11][125] = 5'b00000;
assign A[11][126] = 5'b11101;
assign A[11][127] = 5'b11110;
assign A[11][128] = 5'b00011;
assign A[11][129] = 5'b00100;
assign A[11][130] = 5'b00000;
assign A[11][131] = 5'b11111;
assign A[11][132] = 5'b00001;
assign A[11][133] = 5'b11111;
assign A[11][134] = 5'b00001;
assign A[11][135] = 5'b00000;
assign A[11][136] = 5'b00010;
assign A[11][137] = 5'b00010;
assign A[11][138] = 5'b11111;
assign A[11][139] = 5'b00001;
assign A[11][140] = 5'b11110;
assign A[11][141] = 5'b00011;
assign A[11][142] = 5'b00010;
assign A[11][143] = 5'b00010;
assign A[11][144] = 5'b00000;
assign A[11][145] = 5'b00011;
assign A[11][146] = 5'b00101;
assign A[11][147] = 5'b00010;
assign A[11][148] = 5'b00001;
assign A[11][149] = 5'b11111;
assign A[11][150] = 5'b11110;
assign A[11][151] = 5'b00010;
assign A[11][152] = 5'b00001;
assign A[11][153] = 5'b11110;
assign A[11][154] = 5'b00000;
assign A[11][155] = 5'b00010;
assign A[11][156] = 5'b11111;
assign A[11][157] = 5'b00010;
assign A[11][158] = 5'b11111;
assign A[11][159] = 5'b00001;
assign A[11][160] = 5'b11111;
assign A[11][161] = 5'b00111;
assign A[11][162] = 5'b00001;
assign A[11][163] = 5'b00010;
assign A[11][164] = 5'b11110;
assign A[11][165] = 5'b11111;
assign A[11][166] = 5'b11111;
assign A[11][167] = 5'b00011;
assign A[11][168] = 5'b00011;
assign A[11][169] = 5'b00001;
assign A[11][170] = 5'b00100;
assign A[11][171] = 5'b00001;
assign A[11][172] = 5'b00001;
assign A[11][173] = 5'b00010;
assign A[11][174] = 5'b00010;
assign A[11][175] = 5'b00010;
assign A[11][176] = 5'b00010;
assign A[11][177] = 5'b00010;
assign A[11][178] = 5'b00000;
assign A[11][179] = 5'b00001;
assign A[11][180] = 5'b00010;
assign A[11][181] = 5'b00001;
assign A[11][182] = 5'b11111;
assign A[11][183] = 5'b00001;
assign A[11][184] = 5'b00000;
assign A[11][185] = 5'b00010;
assign A[11][186] = 5'b00000;
assign A[11][187] = 5'b00010;
assign A[11][188] = 5'b11111;
assign A[11][189] = 5'b00010;
assign A[11][190] = 5'b00001;
assign A[11][191] = 5'b00000;
assign A[11][192] = 5'b00000;
assign A[11][193] = 5'b00001;
assign A[11][194] = 5'b00011;
assign A[11][195] = 5'b00001;
assign A[11][196] = 5'b00001;
assign A[11][197] = 5'b00010;
assign A[11][198] = 5'b11110;
assign A[11][199] = 5'b00011;
assign A[11][200] = 5'b11110;
assign A[11][201] = 5'b00000;
assign A[11][202] = 5'b00010;
assign A[11][203] = 5'b00000;
assign A[11][204] = 5'b00000;
assign A[11][205] = 5'b11111;
assign A[11][206] = 5'b00000;
assign A[11][207] = 5'b00001;
assign A[11][208] = 5'b00001;
assign A[11][209] = 5'b11111;
assign A[11][210] = 5'b11111;
assign A[11][211] = 5'b00001;
assign A[11][212] = 5'b11100;
assign A[11][213] = 5'b11111;
assign A[11][214] = 5'b00000;
assign A[11][215] = 5'b00001;
assign A[11][216] = 5'b11111;
assign A[11][217] = 5'b00001;
assign A[11][218] = 5'b11110;
assign A[11][219] = 5'b00000;
assign A[11][220] = 5'b11111;
assign A[11][221] = 5'b00001;
assign A[11][222] = 5'b11101;
assign A[11][223] = 5'b11111;
assign A[11][224] = 5'b00001;
assign A[11][225] = 5'b00001;
assign A[11][226] = 5'b11110;
assign A[11][227] = 5'b11111;
assign A[11][228] = 5'b00000;
assign A[11][229] = 5'b00011;
assign A[11][230] = 5'b11110;
assign A[11][231] = 5'b00000;
assign A[11][232] = 5'b00000;
assign A[11][233] = 5'b11111;
assign A[11][234] = 5'b00000;
assign A[11][235] = 5'b00001;
assign A[11][236] = 5'b00000;
assign A[11][237] = 5'b00000;
assign A[11][238] = 5'b11111;
assign A[11][239] = 5'b11110;
assign A[11][240] = 5'b11111;
assign A[11][241] = 5'b11111;
assign A[11][242] = 5'b00001;
assign A[11][243] = 5'b11111;
assign A[11][244] = 5'b11101;
assign A[11][245] = 5'b11111;
assign A[11][246] = 5'b11111;
assign A[11][247] = 5'b00001;
assign A[11][248] = 5'b00000;
assign A[11][249] = 5'b00000;
assign A[11][250] = 5'b00000;
assign A[11][251] = 5'b11110;
assign A[11][252] = 5'b11111;
assign A[11][253] = 5'b00000;
assign A[11][254] = 5'b11110;
assign A[11][255] = 5'b11111;
assign A[12][0] = 5'b00001;
assign A[12][1] = 5'b11110;
assign A[12][2] = 5'b11110;
assign A[12][3] = 5'b00000;
assign A[12][4] = 5'b00001;
assign A[12][5] = 5'b00010;
assign A[12][6] = 5'b11110;
assign A[12][7] = 5'b00000;
assign A[12][8] = 5'b11101;
assign A[12][9] = 5'b11111;
assign A[12][10] = 5'b11110;
assign A[12][11] = 5'b11111;
assign A[12][12] = 5'b00000;
assign A[12][13] = 5'b00010;
assign A[12][14] = 5'b00001;
assign A[12][15] = 5'b11111;
assign A[12][16] = 5'b11111;
assign A[12][17] = 5'b11111;
assign A[12][18] = 5'b11111;
assign A[12][19] = 5'b00000;
assign A[12][20] = 5'b00000;
assign A[12][21] = 5'b00001;
assign A[12][22] = 5'b11111;
assign A[12][23] = 5'b00001;
assign A[12][24] = 5'b00000;
assign A[12][25] = 5'b11111;
assign A[12][26] = 5'b11111;
assign A[12][27] = 5'b00001;
assign A[12][28] = 5'b00000;
assign A[12][29] = 5'b00001;
assign A[12][30] = 5'b11110;
assign A[12][31] = 5'b11110;
assign A[12][32] = 5'b00001;
assign A[12][33] = 5'b00001;
assign A[12][34] = 5'b00000;
assign A[12][35] = 5'b00000;
assign A[12][36] = 5'b00000;
assign A[12][37] = 5'b00001;
assign A[12][38] = 5'b00000;
assign A[12][39] = 5'b11111;
assign A[12][40] = 5'b11111;
assign A[12][41] = 5'b00001;
assign A[12][42] = 5'b00001;
assign A[12][43] = 5'b00001;
assign A[12][44] = 5'b11111;
assign A[12][45] = 5'b00000;
assign A[12][46] = 5'b00010;
assign A[12][47] = 5'b11111;
assign A[12][48] = 5'b11111;
assign A[12][49] = 5'b00001;
assign A[12][50] = 5'b11101;
assign A[12][51] = 5'b11110;
assign A[12][52] = 5'b00001;
assign A[12][53] = 5'b00011;
assign A[12][54] = 5'b11110;
assign A[12][55] = 5'b00001;
assign A[12][56] = 5'b00010;
assign A[12][57] = 5'b00000;
assign A[12][58] = 5'b00001;
assign A[12][59] = 5'b11111;
assign A[12][60] = 5'b11111;
assign A[12][61] = 5'b00000;
assign A[12][62] = 5'b00010;
assign A[12][63] = 5'b00001;
assign A[12][64] = 5'b00011;
assign A[12][65] = 5'b00000;
assign A[12][66] = 5'b00001;
assign A[12][67] = 5'b00000;
assign A[12][68] = 5'b00001;
assign A[12][69] = 5'b00011;
assign A[12][70] = 5'b11110;
assign A[12][71] = 5'b11101;
assign A[12][72] = 5'b00001;
assign A[12][73] = 5'b00000;
assign A[12][74] = 5'b11101;
assign A[12][75] = 5'b11111;
assign A[12][76] = 5'b11111;
assign A[12][77] = 5'b00001;
assign A[12][78] = 5'b11110;
assign A[12][79] = 5'b11111;
assign A[12][80] = 5'b00001;
assign A[12][81] = 5'b11110;
assign A[12][82] = 5'b11111;
assign A[12][83] = 5'b11110;
assign A[12][84] = 5'b00011;
assign A[12][85] = 5'b00010;
assign A[12][86] = 5'b00001;
assign A[12][87] = 5'b11111;
assign A[12][88] = 5'b00001;
assign A[12][89] = 5'b00000;
assign A[12][90] = 5'b00001;
assign A[12][91] = 5'b11111;
assign A[12][92] = 5'b11110;
assign A[12][93] = 5'b11111;
assign A[12][94] = 5'b00001;
assign A[12][95] = 5'b11111;
assign A[12][96] = 5'b11111;
assign A[12][97] = 5'b00000;
assign A[12][98] = 5'b11111;
assign A[12][99] = 5'b00000;
assign A[12][100] = 5'b11110;
assign A[12][101] = 5'b11111;
assign A[12][102] = 5'b00001;
assign A[12][103] = 5'b00000;
assign A[12][104] = 5'b00001;
assign A[12][105] = 5'b00010;
assign A[12][106] = 5'b11110;
assign A[12][107] = 5'b00000;
assign A[12][108] = 5'b00001;
assign A[12][109] = 5'b00000;
assign A[12][110] = 5'b00001;
assign A[12][111] = 5'b00010;
assign A[12][112] = 5'b00001;
assign A[12][113] = 5'b00010;
assign A[12][114] = 5'b00010;
assign A[12][115] = 5'b11110;
assign A[12][116] = 5'b11101;
assign A[12][117] = 5'b00001;
assign A[12][118] = 5'b11111;
assign A[12][119] = 5'b00000;
assign A[12][120] = 5'b00010;
assign A[12][121] = 5'b00001;
assign A[12][122] = 5'b11101;
assign A[12][123] = 5'b11111;
assign A[12][124] = 5'b11110;
assign A[12][125] = 5'b11110;
assign A[12][126] = 5'b00010;
assign A[12][127] = 5'b11110;
assign A[12][128] = 5'b11101;
assign A[12][129] = 5'b11110;
assign A[12][130] = 5'b11111;
assign A[12][131] = 5'b11111;
assign A[12][132] = 5'b11110;
assign A[12][133] = 5'b00000;
assign A[12][134] = 5'b00011;
assign A[12][135] = 5'b00010;
assign A[12][136] = 5'b00000;
assign A[12][137] = 5'b00000;
assign A[12][138] = 5'b00000;
assign A[12][139] = 5'b00000;
assign A[12][140] = 5'b00011;
assign A[12][141] = 5'b00011;
assign A[12][142] = 5'b00001;
assign A[12][143] = 5'b00010;
assign A[12][144] = 5'b00001;
assign A[12][145] = 5'b00000;
assign A[12][146] = 5'b00001;
assign A[12][147] = 5'b00001;
assign A[12][148] = 5'b11111;
assign A[12][149] = 5'b00000;
assign A[12][150] = 5'b00100;
assign A[12][151] = 5'b00011;
assign A[12][152] = 5'b11111;
assign A[12][153] = 5'b00010;
assign A[12][154] = 5'b00010;
assign A[12][155] = 5'b11101;
assign A[12][156] = 5'b00001;
assign A[12][157] = 5'b00000;
assign A[12][158] = 5'b11110;
assign A[12][159] = 5'b00000;
assign A[12][160] = 5'b00001;
assign A[12][161] = 5'b00000;
assign A[12][162] = 5'b00000;
assign A[12][163] = 5'b11110;
assign A[12][164] = 5'b00010;
assign A[12][165] = 5'b00010;
assign A[12][166] = 5'b00000;
assign A[12][167] = 5'b00010;
assign A[12][168] = 5'b00001;
assign A[12][169] = 5'b00000;
assign A[12][170] = 5'b00010;
assign A[12][171] = 5'b00000;
assign A[12][172] = 5'b11111;
assign A[12][173] = 5'b11111;
assign A[12][174] = 5'b00000;
assign A[12][175] = 5'b00000;
assign A[12][176] = 5'b11110;
assign A[12][177] = 5'b11111;
assign A[12][178] = 5'b00001;
assign A[12][179] = 5'b11110;
assign A[12][180] = 5'b11111;
assign A[12][181] = 5'b11111;
assign A[12][182] = 5'b00000;
assign A[12][183] = 5'b00000;
assign A[12][184] = 5'b00000;
assign A[12][185] = 5'b00010;
assign A[12][186] = 5'b00000;
assign A[12][187] = 5'b11110;
assign A[12][188] = 5'b00010;
assign A[12][189] = 5'b11111;
assign A[12][190] = 5'b11101;
assign A[12][191] = 5'b11111;
assign A[12][192] = 5'b00010;
assign A[12][193] = 5'b00000;
assign A[12][194] = 5'b00001;
assign A[12][195] = 5'b00001;
assign A[12][196] = 5'b11101;
assign A[12][197] = 5'b00000;
assign A[12][198] = 5'b00010;
assign A[12][199] = 5'b11111;
assign A[12][200] = 5'b00001;
assign A[12][201] = 5'b00000;
assign A[12][202] = 5'b00001;
assign A[12][203] = 5'b11111;
assign A[12][204] = 5'b00000;
assign A[12][205] = 5'b11110;
assign A[12][206] = 5'b11111;
assign A[12][207] = 5'b00011;
assign A[12][208] = 5'b00000;
assign A[12][209] = 5'b00000;
assign A[12][210] = 5'b11101;
assign A[12][211] = 5'b00000;
assign A[12][212] = 5'b00000;
assign A[12][213] = 5'b11110;
assign A[12][214] = 5'b00001;
assign A[12][215] = 5'b11111;
assign A[12][216] = 5'b00000;
assign A[12][217] = 5'b00001;
assign A[12][218] = 5'b11110;
assign A[12][219] = 5'b11111;
assign A[12][220] = 5'b00010;
assign A[12][221] = 5'b00011;
assign A[12][222] = 5'b00000;
assign A[12][223] = 5'b11111;
assign A[12][224] = 5'b00001;
assign A[12][225] = 5'b11111;
assign A[12][226] = 5'b11111;
assign A[12][227] = 5'b00001;
assign A[12][228] = 5'b00000;
assign A[12][229] = 5'b11111;
assign A[12][230] = 5'b00000;
assign A[12][231] = 5'b11111;
assign A[12][232] = 5'b11101;
assign A[12][233] = 5'b00001;
assign A[12][234] = 5'b11110;
assign A[12][235] = 5'b00001;
assign A[12][236] = 5'b11111;
assign A[12][237] = 5'b11110;
assign A[12][238] = 5'b00000;
assign A[12][239] = 5'b11110;
assign A[12][240] = 5'b11111;
assign A[12][241] = 5'b00000;
assign A[12][242] = 5'b00010;
assign A[12][243] = 5'b00001;
assign A[12][244] = 5'b00001;
assign A[12][245] = 5'b00000;
assign A[12][246] = 5'b00000;
assign A[12][247] = 5'b00000;
assign A[12][248] = 5'b00000;
assign A[12][249] = 5'b11110;
assign A[12][250] = 5'b00010;
assign A[12][251] = 5'b00100;
assign A[12][252] = 5'b11111;
assign A[12][253] = 5'b11110;
assign A[12][254] = 5'b00000;
assign A[12][255] = 5'b00000;
assign A[13][0] = 5'b00000;
assign A[13][1] = 5'b11111;
assign A[13][2] = 5'b11111;
assign A[13][3] = 5'b00001;
assign A[13][4] = 5'b00100;
assign A[13][5] = 5'b11110;
assign A[13][6] = 5'b00001;
assign A[13][7] = 5'b11111;
assign A[13][8] = 5'b00001;
assign A[13][9] = 5'b00001;
assign A[13][10] = 5'b00000;
assign A[13][11] = 5'b11111;
assign A[13][12] = 5'b00001;
assign A[13][13] = 5'b11111;
assign A[13][14] = 5'b00001;
assign A[13][15] = 5'b00001;
assign A[13][16] = 5'b11110;
assign A[13][17] = 5'b11110;
assign A[13][18] = 5'b00000;
assign A[13][19] = 5'b11111;
assign A[13][20] = 5'b11110;
assign A[13][21] = 5'b00001;
assign A[13][22] = 5'b00001;
assign A[13][23] = 5'b00000;
assign A[13][24] = 5'b00000;
assign A[13][25] = 5'b00000;
assign A[13][26] = 5'b11110;
assign A[13][27] = 5'b11111;
assign A[13][28] = 5'b00010;
assign A[13][29] = 5'b00000;
assign A[13][30] = 5'b00001;
assign A[13][31] = 5'b00001;
assign A[13][32] = 5'b00011;
assign A[13][33] = 5'b00001;
assign A[13][34] = 5'b00000;
assign A[13][35] = 5'b00000;
assign A[13][36] = 5'b11100;
assign A[13][37] = 5'b11111;
assign A[13][38] = 5'b00000;
assign A[13][39] = 5'b00000;
assign A[13][40] = 5'b00000;
assign A[13][41] = 5'b00001;
assign A[13][42] = 5'b00001;
assign A[13][43] = 5'b00001;
assign A[13][44] = 5'b00001;
assign A[13][45] = 5'b00000;
assign A[13][46] = 5'b11111;
assign A[13][47] = 5'b00000;
assign A[13][48] = 5'b00010;
assign A[13][49] = 5'b00000;
assign A[13][50] = 5'b00001;
assign A[13][51] = 5'b00011;
assign A[13][52] = 5'b00010;
assign A[13][53] = 5'b00000;
assign A[13][54] = 5'b11110;
assign A[13][55] = 5'b00000;
assign A[13][56] = 5'b11111;
assign A[13][57] = 5'b11111;
assign A[13][58] = 5'b00000;
assign A[13][59] = 5'b11110;
assign A[13][60] = 5'b11101;
assign A[13][61] = 5'b00001;
assign A[13][62] = 5'b00001;
assign A[13][63] = 5'b00011;
assign A[13][64] = 5'b00001;
assign A[13][65] = 5'b00001;
assign A[13][66] = 5'b00000;
assign A[13][67] = 5'b11110;
assign A[13][68] = 5'b00001;
assign A[13][69] = 5'b00001;
assign A[13][70] = 5'b11101;
assign A[13][71] = 5'b00000;
assign A[13][72] = 5'b00011;
assign A[13][73] = 5'b11111;
assign A[13][74] = 5'b00000;
assign A[13][75] = 5'b00001;
assign A[13][76] = 5'b00000;
assign A[13][77] = 5'b00001;
assign A[13][78] = 5'b00000;
assign A[13][79] = 5'b11110;
assign A[13][80] = 5'b00000;
assign A[13][81] = 5'b11111;
assign A[13][82] = 5'b00011;
assign A[13][83] = 5'b00001;
assign A[13][84] = 5'b11110;
assign A[13][85] = 5'b11110;
assign A[13][86] = 5'b00000;
assign A[13][87] = 5'b11110;
assign A[13][88] = 5'b00001;
assign A[13][89] = 5'b00001;
assign A[13][90] = 5'b11110;
assign A[13][91] = 5'b11111;
assign A[13][92] = 5'b00010;
assign A[13][93] = 5'b00010;
assign A[13][94] = 5'b00001;
assign A[13][95] = 5'b00001;
assign A[13][96] = 5'b00000;
assign A[13][97] = 5'b11101;
assign A[13][98] = 5'b00001;
assign A[13][99] = 5'b00010;
assign A[13][100] = 5'b00000;
assign A[13][101] = 5'b00001;
assign A[13][102] = 5'b00001;
assign A[13][103] = 5'b11110;
assign A[13][104] = 5'b11111;
assign A[13][105] = 5'b00000;
assign A[13][106] = 5'b11111;
assign A[13][107] = 5'b00001;
assign A[13][108] = 5'b00001;
assign A[13][109] = 5'b11111;
assign A[13][110] = 5'b00000;
assign A[13][111] = 5'b00000;
assign A[13][112] = 5'b00001;
assign A[13][113] = 5'b11111;
assign A[13][114] = 5'b11111;
assign A[13][115] = 5'b00000;
assign A[13][116] = 5'b00000;
assign A[13][117] = 5'b11111;
assign A[13][118] = 5'b11111;
assign A[13][119] = 5'b00001;
assign A[13][120] = 5'b11111;
assign A[13][121] = 5'b00001;
assign A[13][122] = 5'b00000;
assign A[13][123] = 5'b00001;
assign A[13][124] = 5'b00000;
assign A[13][125] = 5'b00001;
assign A[13][126] = 5'b11111;
assign A[13][127] = 5'b00001;
assign A[13][128] = 5'b00010;
assign A[13][129] = 5'b00000;
assign A[13][130] = 5'b11110;
assign A[13][131] = 5'b00010;
assign A[13][132] = 5'b00000;
assign A[13][133] = 5'b00001;
assign A[13][134] = 5'b11110;
assign A[13][135] = 5'b11111;
assign A[13][136] = 5'b00000;
assign A[13][137] = 5'b11111;
assign A[13][138] = 5'b00000;
assign A[13][139] = 5'b11110;
assign A[13][140] = 5'b11111;
assign A[13][141] = 5'b11110;
assign A[13][142] = 5'b00000;
assign A[13][143] = 5'b11011;
assign A[13][144] = 5'b00001;
assign A[13][145] = 5'b00000;
assign A[13][146] = 5'b11111;
assign A[13][147] = 5'b00000;
assign A[13][148] = 5'b11110;
assign A[13][149] = 5'b00000;
assign A[13][150] = 5'b00010;
assign A[13][151] = 5'b00000;
assign A[13][152] = 5'b00010;
assign A[13][153] = 5'b00010;
assign A[13][154] = 5'b00000;
assign A[13][155] = 5'b00000;
assign A[13][156] = 5'b00001;
assign A[13][157] = 5'b00010;
assign A[13][158] = 5'b00001;
assign A[13][159] = 5'b11110;
assign A[13][160] = 5'b00001;
assign A[13][161] = 5'b00010;
assign A[13][162] = 5'b11111;
assign A[13][163] = 5'b00000;
assign A[13][164] = 5'b00000;
assign A[13][165] = 5'b00001;
assign A[13][166] = 5'b11111;
assign A[13][167] = 5'b00011;
assign A[13][168] = 5'b11111;
assign A[13][169] = 5'b11111;
assign A[13][170] = 5'b00000;
assign A[13][171] = 5'b11111;
assign A[13][172] = 5'b11110;
assign A[13][173] = 5'b00001;
assign A[13][174] = 5'b11111;
assign A[13][175] = 5'b00010;
assign A[13][176] = 5'b00010;
assign A[13][177] = 5'b00000;
assign A[13][178] = 5'b00000;
assign A[13][179] = 5'b00001;
assign A[13][180] = 5'b00001;
assign A[13][181] = 5'b00010;
assign A[13][182] = 5'b00001;
assign A[13][183] = 5'b00000;
assign A[13][184] = 5'b00010;
assign A[13][185] = 5'b00000;
assign A[13][186] = 5'b11111;
assign A[13][187] = 5'b11110;
assign A[13][188] = 5'b00000;
assign A[13][189] = 5'b11111;
assign A[13][190] = 5'b00000;
assign A[13][191] = 5'b00010;
assign A[13][192] = 5'b00011;
assign A[13][193] = 5'b11110;
assign A[13][194] = 5'b00001;
assign A[13][195] = 5'b00010;
assign A[13][196] = 5'b00000;
assign A[13][197] = 5'b00000;
assign A[13][198] = 5'b00001;
assign A[13][199] = 5'b00001;
assign A[13][200] = 5'b00000;
assign A[13][201] = 5'b00001;
assign A[13][202] = 5'b00001;
assign A[13][203] = 5'b11111;
assign A[13][204] = 5'b00001;
assign A[13][205] = 5'b00011;
assign A[13][206] = 5'b00000;
assign A[13][207] = 5'b11111;
assign A[13][208] = 5'b00010;
assign A[13][209] = 5'b00000;
assign A[13][210] = 5'b00010;
assign A[13][211] = 5'b11111;
assign A[13][212] = 5'b00000;
assign A[13][213] = 5'b00010;
assign A[13][214] = 5'b00000;
assign A[13][215] = 5'b11111;
assign A[13][216] = 5'b11111;
assign A[13][217] = 5'b00011;
assign A[13][218] = 5'b00000;
assign A[13][219] = 5'b00000;
assign A[13][220] = 5'b00011;
assign A[13][221] = 5'b00000;
assign A[13][222] = 5'b11111;
assign A[13][223] = 5'b11111;
assign A[13][224] = 5'b00010;
assign A[13][225] = 5'b11111;
assign A[13][226] = 5'b11110;
assign A[13][227] = 5'b00000;
assign A[13][228] = 5'b11111;
assign A[13][229] = 5'b00010;
assign A[13][230] = 5'b00010;
assign A[13][231] = 5'b00011;
assign A[13][232] = 5'b00000;
assign A[13][233] = 5'b00011;
assign A[13][234] = 5'b00000;
assign A[13][235] = 5'b00001;
assign A[13][236] = 5'b11111;
assign A[13][237] = 5'b11111;
assign A[13][238] = 5'b00000;
assign A[13][239] = 5'b11110;
assign A[13][240] = 5'b00000;
assign A[13][241] = 5'b11111;
assign A[13][242] = 5'b11110;
assign A[13][243] = 5'b00000;
assign A[13][244] = 5'b00010;
assign A[13][245] = 5'b00001;
assign A[13][246] = 5'b00010;
assign A[13][247] = 5'b11110;
assign A[13][248] = 5'b00001;
assign A[13][249] = 5'b11111;
assign A[13][250] = 5'b00001;
assign A[13][251] = 5'b00001;
assign A[13][252] = 5'b11110;
assign A[13][253] = 5'b11111;
assign A[13][254] = 5'b00001;
assign A[13][255] = 5'b00000;
assign A[14][0] = 5'b00001;
assign A[14][1] = 5'b11100;
assign A[14][2] = 5'b00000;
assign A[14][3] = 5'b11111;
assign A[14][4] = 5'b11111;
assign A[14][5] = 5'b00010;
assign A[14][6] = 5'b00001;
assign A[14][7] = 5'b00010;
assign A[14][8] = 5'b00001;
assign A[14][9] = 5'b00000;
assign A[14][10] = 5'b11111;
assign A[14][11] = 5'b11111;
assign A[14][12] = 5'b11111;
assign A[14][13] = 5'b00000;
assign A[14][14] = 5'b00000;
assign A[14][15] = 5'b11101;
assign A[14][16] = 5'b00000;
assign A[14][17] = 5'b00011;
assign A[14][18] = 5'b00001;
assign A[14][19] = 5'b11111;
assign A[14][20] = 5'b00000;
assign A[14][21] = 5'b11101;
assign A[14][22] = 5'b00000;
assign A[14][23] = 5'b00001;
assign A[14][24] = 5'b00011;
assign A[14][25] = 5'b00000;
assign A[14][26] = 5'b00000;
assign A[14][27] = 5'b00010;
assign A[14][28] = 5'b00000;
assign A[14][29] = 5'b00000;
assign A[14][30] = 5'b11110;
assign A[14][31] = 5'b00000;
assign A[14][32] = 5'b11111;
assign A[14][33] = 5'b00100;
assign A[14][34] = 5'b11111;
assign A[14][35] = 5'b11110;
assign A[14][36] = 5'b11111;
assign A[14][37] = 5'b00010;
assign A[14][38] = 5'b11111;
assign A[14][39] = 5'b00010;
assign A[14][40] = 5'b11111;
assign A[14][41] = 5'b00000;
assign A[14][42] = 5'b11110;
assign A[14][43] = 5'b00000;
assign A[14][44] = 5'b11110;
assign A[14][45] = 5'b11101;
assign A[14][46] = 5'b11110;
assign A[14][47] = 5'b00001;
assign A[14][48] = 5'b00001;
assign A[14][49] = 5'b00011;
assign A[14][50] = 5'b00011;
assign A[14][51] = 5'b11110;
assign A[14][52] = 5'b00001;
assign A[14][53] = 5'b00000;
assign A[14][54] = 5'b00001;
assign A[14][55] = 5'b11101;
assign A[14][56] = 5'b00001;
assign A[14][57] = 5'b11110;
assign A[14][58] = 5'b00000;
assign A[14][59] = 5'b11111;
assign A[14][60] = 5'b11111;
assign A[14][61] = 5'b11111;
assign A[14][62] = 5'b00001;
assign A[14][63] = 5'b00010;
assign A[14][64] = 5'b00001;
assign A[14][65] = 5'b00010;
assign A[14][66] = 5'b00001;
assign A[14][67] = 5'b00000;
assign A[14][68] = 5'b00001;
assign A[14][69] = 5'b00001;
assign A[14][70] = 5'b00000;
assign A[14][71] = 5'b00000;
assign A[14][72] = 5'b11111;
assign A[14][73] = 5'b00001;
assign A[14][74] = 5'b11110;
assign A[14][75] = 5'b00010;
assign A[14][76] = 5'b11111;
assign A[14][77] = 5'b11110;
assign A[14][78] = 5'b00000;
assign A[14][79] = 5'b11111;
assign A[14][80] = 5'b11110;
assign A[14][81] = 5'b00000;
assign A[14][82] = 5'b00100;
assign A[14][83] = 5'b00000;
assign A[14][84] = 5'b00000;
assign A[14][85] = 5'b00000;
assign A[14][86] = 5'b00100;
assign A[14][87] = 5'b11101;
assign A[14][88] = 5'b00001;
assign A[14][89] = 5'b00000;
assign A[14][90] = 5'b00000;
assign A[14][91] = 5'b00000;
assign A[14][92] = 5'b00000;
assign A[14][93] = 5'b00000;
assign A[14][94] = 5'b00001;
assign A[14][95] = 5'b11111;
assign A[14][96] = 5'b11111;
assign A[14][97] = 5'b00000;
assign A[14][98] = 5'b00001;
assign A[14][99] = 5'b11101;
assign A[14][100] = 5'b00000;
assign A[14][101] = 5'b11111;
assign A[14][102] = 5'b00010;
assign A[14][103] = 5'b11101;
assign A[14][104] = 5'b00000;
assign A[14][105] = 5'b11111;
assign A[14][106] = 5'b11111;
assign A[14][107] = 5'b00001;
assign A[14][108] = 5'b00000;
assign A[14][109] = 5'b00001;
assign A[14][110] = 5'b00001;
assign A[14][111] = 5'b11110;
assign A[14][112] = 5'b11110;
assign A[14][113] = 5'b00001;
assign A[14][114] = 5'b11101;
assign A[14][115] = 5'b00001;
assign A[14][116] = 5'b11111;
assign A[14][117] = 5'b00001;
assign A[14][118] = 5'b11111;
assign A[14][119] = 5'b00000;
assign A[14][120] = 5'b00000;
assign A[14][121] = 5'b00000;
assign A[14][122] = 5'b00000;
assign A[14][123] = 5'b00001;
assign A[14][124] = 5'b00001;
assign A[14][125] = 5'b11110;
assign A[14][126] = 5'b00010;
assign A[14][127] = 5'b00000;
assign A[14][128] = 5'b00001;
assign A[14][129] = 5'b11111;
assign A[14][130] = 5'b00000;
assign A[14][131] = 5'b11101;
assign A[14][132] = 5'b00001;
assign A[14][133] = 5'b11111;
assign A[14][134] = 5'b11111;
assign A[14][135] = 5'b11111;
assign A[14][136] = 5'b00000;
assign A[14][137] = 5'b11110;
assign A[14][138] = 5'b00100;
assign A[14][139] = 5'b00001;
assign A[14][140] = 5'b00000;
assign A[14][141] = 5'b11111;
assign A[14][142] = 5'b11111;
assign A[14][143] = 5'b00000;
assign A[14][144] = 5'b00000;
assign A[14][145] = 5'b11111;
assign A[14][146] = 5'b11111;
assign A[14][147] = 5'b11111;
assign A[14][148] = 5'b00000;
assign A[14][149] = 5'b11111;
assign A[14][150] = 5'b11111;
assign A[14][151] = 5'b11111;
assign A[14][152] = 5'b00000;
assign A[14][153] = 5'b00001;
assign A[14][154] = 5'b11111;
assign A[14][155] = 5'b00010;
assign A[14][156] = 5'b00001;
assign A[14][157] = 5'b11110;
assign A[14][158] = 5'b00000;
assign A[14][159] = 5'b11111;
assign A[14][160] = 5'b00001;
assign A[14][161] = 5'b00010;
assign A[14][162] = 5'b00000;
assign A[14][163] = 5'b00000;
assign A[14][164] = 5'b11110;
assign A[14][165] = 5'b00001;
assign A[14][166] = 5'b00000;
assign A[14][167] = 5'b00000;
assign A[14][168] = 5'b00000;
assign A[14][169] = 5'b00001;
assign A[14][170] = 5'b00000;
assign A[14][171] = 5'b11111;
assign A[14][172] = 5'b00000;
assign A[14][173] = 5'b00011;
assign A[14][174] = 5'b00001;
assign A[14][175] = 5'b00001;
assign A[14][176] = 5'b00000;
assign A[14][177] = 5'b00001;
assign A[14][178] = 5'b11111;
assign A[14][179] = 5'b00000;
assign A[14][180] = 5'b00010;
assign A[14][181] = 5'b00001;
assign A[14][182] = 5'b11111;
assign A[14][183] = 5'b11100;
assign A[14][184] = 5'b00000;
assign A[14][185] = 5'b11111;
assign A[14][186] = 5'b00000;
assign A[14][187] = 5'b00010;
assign A[14][188] = 5'b00000;
assign A[14][189] = 5'b11111;
assign A[14][190] = 5'b00010;
assign A[14][191] = 5'b00001;
assign A[14][192] = 5'b00000;
assign A[14][193] = 5'b11110;
assign A[14][194] = 5'b11111;
assign A[14][195] = 5'b00011;
assign A[14][196] = 5'b00001;
assign A[14][197] = 5'b00000;
assign A[14][198] = 5'b00011;
assign A[14][199] = 5'b00000;
assign A[14][200] = 5'b11110;
assign A[14][201] = 5'b11111;
assign A[14][202] = 5'b00001;
assign A[14][203] = 5'b00011;
assign A[14][204] = 5'b00001;
assign A[14][205] = 5'b00001;
assign A[14][206] = 5'b11111;
assign A[14][207] = 5'b11111;
assign A[14][208] = 5'b00011;
assign A[14][209] = 5'b11111;
assign A[14][210] = 5'b11101;
assign A[14][211] = 5'b00000;
assign A[14][212] = 5'b00000;
assign A[14][213] = 5'b11101;
assign A[14][214] = 5'b11111;
assign A[14][215] = 5'b00000;
assign A[14][216] = 5'b00001;
assign A[14][217] = 5'b00000;
assign A[14][218] = 5'b00010;
assign A[14][219] = 5'b00001;
assign A[14][220] = 5'b11111;
assign A[14][221] = 5'b11111;
assign A[14][222] = 5'b00000;
assign A[14][223] = 5'b00001;
assign A[14][224] = 5'b11101;
assign A[14][225] = 5'b11111;
assign A[14][226] = 5'b00000;
assign A[14][227] = 5'b11111;
assign A[14][228] = 5'b00001;
assign A[14][229] = 5'b00001;
assign A[14][230] = 5'b11111;
assign A[14][231] = 5'b11111;
assign A[14][232] = 5'b11111;
assign A[14][233] = 5'b00001;
assign A[14][234] = 5'b00001;
assign A[14][235] = 5'b11111;
assign A[14][236] = 5'b11111;
assign A[14][237] = 5'b00000;
assign A[14][238] = 5'b11111;
assign A[14][239] = 5'b11111;
assign A[14][240] = 5'b00001;
assign A[14][241] = 5'b11110;
assign A[14][242] = 5'b00000;
assign A[14][243] = 5'b00010;
assign A[14][244] = 5'b00000;
assign A[14][245] = 5'b00000;
assign A[14][246] = 5'b11111;
assign A[14][247] = 5'b00000;
assign A[14][248] = 5'b11110;
assign A[14][249] = 5'b11011;
assign A[14][250] = 5'b00001;
assign A[14][251] = 5'b11111;
assign A[14][252] = 5'b11111;
assign A[14][253] = 5'b00010;
assign A[14][254] = 5'b00011;
assign A[14][255] = 5'b00011;
assign A[15][0] = 5'b00000;
assign A[15][1] = 5'b00010;
assign A[15][2] = 5'b00010;
assign A[15][3] = 5'b11110;
assign A[15][4] = 5'b00000;
assign A[15][5] = 5'b00000;
assign A[15][6] = 5'b00000;
assign A[15][7] = 5'b11111;
assign A[15][8] = 5'b00000;
assign A[15][9] = 5'b00001;
assign A[15][10] = 5'b11110;
assign A[15][11] = 5'b11111;
assign A[15][12] = 5'b11111;
assign A[15][13] = 5'b11110;
assign A[15][14] = 5'b00000;
assign A[15][15] = 5'b11111;
assign A[15][16] = 5'b11111;
assign A[15][17] = 5'b11111;
assign A[15][18] = 5'b11111;
assign A[15][19] = 5'b11111;
assign A[15][20] = 5'b00001;
assign A[15][21] = 5'b11110;
assign A[15][22] = 5'b11110;
assign A[15][23] = 5'b00000;
assign A[15][24] = 5'b11111;
assign A[15][25] = 5'b00000;
assign A[15][26] = 5'b11110;
assign A[15][27] = 5'b11111;
assign A[15][28] = 5'b11110;
assign A[15][29] = 5'b00001;
assign A[15][30] = 5'b00000;
assign A[15][31] = 5'b11111;
assign A[15][32] = 5'b11110;
assign A[15][33] = 5'b00001;
assign A[15][34] = 5'b11110;
assign A[15][35] = 5'b00001;
assign A[15][36] = 5'b11110;
assign A[15][37] = 5'b11111;
assign A[15][38] = 5'b11110;
assign A[15][39] = 5'b00000;
assign A[15][40] = 5'b00001;
assign A[15][41] = 5'b00001;
assign A[15][42] = 5'b11101;
assign A[15][43] = 5'b11110;
assign A[15][44] = 5'b11111;
assign A[15][45] = 5'b11111;
assign A[15][46] = 5'b00000;
assign A[15][47] = 5'b00010;
assign A[15][48] = 5'b00000;
assign A[15][49] = 5'b00010;
assign A[15][50] = 5'b00010;
assign A[15][51] = 5'b00000;
assign A[15][52] = 5'b11111;
assign A[15][53] = 5'b11111;
assign A[15][54] = 5'b00010;
assign A[15][55] = 5'b11111;
assign A[15][56] = 5'b00001;
assign A[15][57] = 5'b00001;
assign A[15][58] = 5'b00100;
assign A[15][59] = 5'b11111;
assign A[15][60] = 5'b00001;
assign A[15][61] = 5'b11110;
assign A[15][62] = 5'b00000;
assign A[15][63] = 5'b00000;
assign A[15][64] = 5'b11111;
assign A[15][65] = 5'b00001;
assign A[15][66] = 5'b00000;
assign A[15][67] = 5'b00001;
assign A[15][68] = 5'b00000;
assign A[15][69] = 5'b11111;
assign A[15][70] = 5'b00010;
assign A[15][71] = 5'b00010;
assign A[15][72] = 5'b11111;
assign A[15][73] = 5'b11110;
assign A[15][74] = 5'b11101;
assign A[15][75] = 5'b00001;
assign A[15][76] = 5'b11111;
assign A[15][77] = 5'b00000;
assign A[15][78] = 5'b00001;
assign A[15][79] = 5'b00000;
assign A[15][80] = 5'b00001;
assign A[15][81] = 5'b11101;
assign A[15][82] = 5'b00000;
assign A[15][83] = 5'b11110;
assign A[15][84] = 5'b00000;
assign A[15][85] = 5'b00010;
assign A[15][86] = 5'b11110;
assign A[15][87] = 5'b00000;
assign A[15][88] = 5'b00000;
assign A[15][89] = 5'b00000;
assign A[15][90] = 5'b00000;
assign A[15][91] = 5'b00001;
assign A[15][92] = 5'b00001;
assign A[15][93] = 5'b11110;
assign A[15][94] = 5'b00001;
assign A[15][95] = 5'b00000;
assign A[15][96] = 5'b00001;
assign A[15][97] = 5'b11111;
assign A[15][98] = 5'b00001;
assign A[15][99] = 5'b00011;
assign A[15][100] = 5'b11101;
assign A[15][101] = 5'b00011;
assign A[15][102] = 5'b00001;
assign A[15][103] = 5'b11111;
assign A[15][104] = 5'b00001;
assign A[15][105] = 5'b11110;
assign A[15][106] = 5'b00001;
assign A[15][107] = 5'b11111;
assign A[15][108] = 5'b11111;
assign A[15][109] = 5'b00001;
assign A[15][110] = 5'b00000;
assign A[15][111] = 5'b11110;
assign A[15][112] = 5'b00000;
assign A[15][113] = 5'b11111;
assign A[15][114] = 5'b11111;
assign A[15][115] = 5'b00010;
assign A[15][116] = 5'b00000;
assign A[15][117] = 5'b11111;
assign A[15][118] = 5'b00001;
assign A[15][119] = 5'b11111;
assign A[15][120] = 5'b00000;
assign A[15][121] = 5'b00000;
assign A[15][122] = 5'b00000;
assign A[15][123] = 5'b00000;
assign A[15][124] = 5'b00000;
assign A[15][125] = 5'b11101;
assign A[15][126] = 5'b00010;
assign A[15][127] = 5'b00001;
assign A[15][128] = 5'b11111;
assign A[15][129] = 5'b00000;
assign A[15][130] = 5'b11111;
assign A[15][131] = 5'b11111;
assign A[15][132] = 5'b11110;
assign A[15][133] = 5'b11111;
assign A[15][134] = 5'b11110;
assign A[15][135] = 5'b11110;
assign A[15][136] = 5'b00000;
assign A[15][137] = 5'b00001;
assign A[15][138] = 5'b00000;
assign A[15][139] = 5'b11110;
assign A[15][140] = 5'b00011;
assign A[15][141] = 5'b00001;
assign A[15][142] = 5'b00000;
assign A[15][143] = 5'b11110;
assign A[15][144] = 5'b11111;
assign A[15][145] = 5'b11110;
assign A[15][146] = 5'b00001;
assign A[15][147] = 5'b00000;
assign A[15][148] = 5'b11111;
assign A[15][149] = 5'b00000;
assign A[15][150] = 5'b00000;
assign A[15][151] = 5'b11111;
assign A[15][152] = 5'b11110;
assign A[15][153] = 5'b11111;
assign A[15][154] = 5'b11101;
assign A[15][155] = 5'b00000;
assign A[15][156] = 5'b00100;
assign A[15][157] = 5'b00000;
assign A[15][158] = 5'b11111;
assign A[15][159] = 5'b00001;
assign A[15][160] = 5'b00001;
assign A[15][161] = 5'b00000;
assign A[15][162] = 5'b11111;
assign A[15][163] = 5'b11111;
assign A[15][164] = 5'b00000;
assign A[15][165] = 5'b00001;
assign A[15][166] = 5'b00001;
assign A[15][167] = 5'b00000;
assign A[15][168] = 5'b00000;
assign A[15][169] = 5'b11101;
assign A[15][170] = 5'b00010;
assign A[15][171] = 5'b00000;
assign A[15][172] = 5'b11110;
assign A[15][173] = 5'b11101;
assign A[15][174] = 5'b11111;
assign A[15][175] = 5'b00001;
assign A[15][176] = 5'b11111;
assign A[15][177] = 5'b11110;
assign A[15][178] = 5'b11110;
assign A[15][179] = 5'b11111;
assign A[15][180] = 5'b00001;
assign A[15][181] = 5'b11110;
assign A[15][182] = 5'b11111;
assign A[15][183] = 5'b00000;
assign A[15][184] = 5'b00001;
assign A[15][185] = 5'b00001;
assign A[15][186] = 5'b11111;
assign A[15][187] = 5'b00000;
assign A[15][188] = 5'b00001;
assign A[15][189] = 5'b11101;
assign A[15][190] = 5'b00010;
assign A[15][191] = 5'b00000;
assign A[15][192] = 5'b00001;
assign A[15][193] = 5'b00001;
assign A[15][194] = 5'b00000;
assign A[15][195] = 5'b11111;
assign A[15][196] = 5'b11111;
assign A[15][197] = 5'b00000;
assign A[15][198] = 5'b11110;
assign A[15][199] = 5'b11111;
assign A[15][200] = 5'b11111;
assign A[15][201] = 5'b00000;
assign A[15][202] = 5'b00010;
assign A[15][203] = 5'b00000;
assign A[15][204] = 5'b11111;
assign A[15][205] = 5'b11111;
assign A[15][206] = 5'b11111;
assign A[15][207] = 5'b00000;
assign A[15][208] = 5'b00000;
assign A[15][209] = 5'b00001;
assign A[15][210] = 5'b00001;
assign A[15][211] = 5'b00000;
assign A[15][212] = 5'b11111;
assign A[15][213] = 5'b11110;
assign A[15][214] = 5'b00010;
assign A[15][215] = 5'b11111;
assign A[15][216] = 5'b00001;
assign A[15][217] = 5'b00001;
assign A[15][218] = 5'b11111;
assign A[15][219] = 5'b00001;
assign A[15][220] = 5'b11110;
assign A[15][221] = 5'b11111;
assign A[15][222] = 5'b11110;
assign A[15][223] = 5'b11111;
assign A[15][224] = 5'b00000;
assign A[15][225] = 5'b00011;
assign A[15][226] = 5'b00000;
assign A[15][227] = 5'b00010;
assign A[15][228] = 5'b00000;
assign A[15][229] = 5'b11111;
assign A[15][230] = 5'b00000;
assign A[15][231] = 5'b00000;
assign A[15][232] = 5'b11111;
assign A[15][233] = 5'b00001;
assign A[15][234] = 5'b11111;
assign A[15][235] = 5'b00000;
assign A[15][236] = 5'b00000;
assign A[15][237] = 5'b00010;
assign A[15][238] = 5'b11111;
assign A[15][239] = 5'b00000;
assign A[15][240] = 5'b00010;
assign A[15][241] = 5'b00001;
assign A[15][242] = 5'b00010;
assign A[15][243] = 5'b11110;
assign A[15][244] = 5'b00000;
assign A[15][245] = 5'b11111;
assign A[15][246] = 5'b00001;
assign A[15][247] = 5'b00000;
assign A[15][248] = 5'b11101;
assign A[15][249] = 5'b00000;
assign A[15][250] = 5'b00010;
assign A[15][251] = 5'b00001;
assign A[15][252] = 5'b00001;
assign A[15][253] = 5'b00000;
assign A[15][254] = 5'b00001;
assign A[15][255] = 5'b11111;
assign A[16][0] = 5'b00000;
assign A[16][1] = 5'b00000;
assign A[16][2] = 5'b11111;
assign A[16][3] = 5'b11110;
assign A[16][4] = 5'b00000;
assign A[16][5] = 5'b00010;
assign A[16][6] = 5'b11110;
assign A[16][7] = 5'b11111;
assign A[16][8] = 5'b11111;
assign A[16][9] = 5'b00010;
assign A[16][10] = 5'b11111;
assign A[16][11] = 5'b00000;
assign A[16][12] = 5'b00011;
assign A[16][13] = 5'b11110;
assign A[16][14] = 5'b11100;
assign A[16][15] = 5'b11110;
assign A[16][16] = 5'b00011;
assign A[16][17] = 5'b00000;
assign A[16][18] = 5'b11111;
assign A[16][19] = 5'b11101;
assign A[16][20] = 5'b11111;
assign A[16][21] = 5'b11110;
assign A[16][22] = 5'b11111;
assign A[16][23] = 5'b11110;
assign A[16][24] = 5'b11111;
assign A[16][25] = 5'b00000;
assign A[16][26] = 5'b11111;
assign A[16][27] = 5'b00001;
assign A[16][28] = 5'b11101;
assign A[16][29] = 5'b00000;
assign A[16][30] = 5'b00001;
assign A[16][31] = 5'b00000;
assign A[16][32] = 5'b00000;
assign A[16][33] = 5'b00001;
assign A[16][34] = 5'b00000;
assign A[16][35] = 5'b00000;
assign A[16][36] = 5'b11110;
assign A[16][37] = 5'b11111;
assign A[16][38] = 5'b00000;
assign A[16][39] = 5'b00001;
assign A[16][40] = 5'b00000;
assign A[16][41] = 5'b11110;
assign A[16][42] = 5'b11111;
assign A[16][43] = 5'b11110;
assign A[16][44] = 5'b11110;
assign A[16][45] = 5'b11110;
assign A[16][46] = 5'b00010;
assign A[16][47] = 5'b11110;
assign A[16][48] = 5'b00000;
assign A[16][49] = 5'b00000;
assign A[16][50] = 5'b00001;
assign A[16][51] = 5'b00010;
assign A[16][52] = 5'b00001;
assign A[16][53] = 5'b11111;
assign A[16][54] = 5'b00010;
assign A[16][55] = 5'b11111;
assign A[16][56] = 5'b11111;
assign A[16][57] = 5'b00001;
assign A[16][58] = 5'b11111;
assign A[16][59] = 5'b11111;
assign A[16][60] = 5'b00001;
assign A[16][61] = 5'b11111;
assign A[16][62] = 5'b11111;
assign A[16][63] = 5'b00001;
assign A[16][64] = 5'b00001;
assign A[16][65] = 5'b11110;
assign A[16][66] = 5'b11110;
assign A[16][67] = 5'b11111;
assign A[16][68] = 5'b00000;
assign A[16][69] = 5'b11111;
assign A[16][70] = 5'b00000;
assign A[16][71] = 5'b11111;
assign A[16][72] = 5'b00000;
assign A[16][73] = 5'b11111;
assign A[16][74] = 5'b00011;
assign A[16][75] = 5'b00000;
assign A[16][76] = 5'b00101;
assign A[16][77] = 5'b11111;
assign A[16][78] = 5'b00001;
assign A[16][79] = 5'b11111;
assign A[16][80] = 5'b11110;
assign A[16][81] = 5'b00001;
assign A[16][82] = 5'b11111;
assign A[16][83] = 5'b11101;
assign A[16][84] = 5'b11111;
assign A[16][85] = 5'b11101;
assign A[16][86] = 5'b11111;
assign A[16][87] = 5'b00010;
assign A[16][88] = 5'b00001;
assign A[16][89] = 5'b11110;
assign A[16][90] = 5'b00000;
assign A[16][91] = 5'b11110;
assign A[16][92] = 5'b00010;
assign A[16][93] = 5'b00001;
assign A[16][94] = 5'b11111;
assign A[16][95] = 5'b00000;
assign A[16][96] = 5'b00001;
assign A[16][97] = 5'b00001;
assign A[16][98] = 5'b00000;
assign A[16][99] = 5'b00001;
assign A[16][100] = 5'b00001;
assign A[16][101] = 5'b00010;
assign A[16][102] = 5'b11100;
assign A[16][103] = 5'b11111;
assign A[16][104] = 5'b00000;
assign A[16][105] = 5'b00001;
assign A[16][106] = 5'b11110;
assign A[16][107] = 5'b00011;
assign A[16][108] = 5'b00001;
assign A[16][109] = 5'b00001;
assign A[16][110] = 5'b00001;
assign A[16][111] = 5'b11110;
assign A[16][112] = 5'b00000;
assign A[16][113] = 5'b00000;
assign A[16][114] = 5'b11111;
assign A[16][115] = 5'b11111;
assign A[16][116] = 5'b00000;
assign A[16][117] = 5'b00010;
assign A[16][118] = 5'b11110;
assign A[16][119] = 5'b00000;
assign A[16][120] = 5'b11111;
assign A[16][121] = 5'b00001;
assign A[16][122] = 5'b00000;
assign A[16][123] = 5'b11111;
assign A[16][124] = 5'b00011;
assign A[16][125] = 5'b00001;
assign A[16][126] = 5'b11110;
assign A[16][127] = 5'b11111;
assign A[16][128] = 5'b00000;
assign A[16][129] = 5'b00010;
assign A[16][130] = 5'b00010;
assign A[16][131] = 5'b11111;
assign A[16][132] = 5'b00001;
assign A[16][133] = 5'b00000;
assign A[16][134] = 5'b00001;
assign A[16][135] = 5'b11110;
assign A[16][136] = 5'b00000;
assign A[16][137] = 5'b00000;
assign A[16][138] = 5'b00000;
assign A[16][139] = 5'b11110;
assign A[16][140] = 5'b11111;
assign A[16][141] = 5'b11110;
assign A[16][142] = 5'b11111;
assign A[16][143] = 5'b11111;
assign A[16][144] = 5'b00000;
assign A[16][145] = 5'b00001;
assign A[16][146] = 5'b00000;
assign A[16][147] = 5'b00011;
assign A[16][148] = 5'b00000;
assign A[16][149] = 5'b00000;
assign A[16][150] = 5'b00001;
assign A[16][151] = 5'b11101;
assign A[16][152] = 5'b00001;
assign A[16][153] = 5'b11110;
assign A[16][154] = 5'b00000;
assign A[16][155] = 5'b00001;
assign A[16][156] = 5'b11111;
assign A[16][157] = 5'b11110;
assign A[16][158] = 5'b11111;
assign A[16][159] = 5'b11110;
assign A[16][160] = 5'b00010;
assign A[16][161] = 5'b00000;
assign A[16][162] = 5'b00010;
assign A[16][163] = 5'b00000;
assign A[16][164] = 5'b00010;
assign A[16][165] = 5'b11111;
assign A[16][166] = 5'b11110;
assign A[16][167] = 5'b00010;
assign A[16][168] = 5'b00010;
assign A[16][169] = 5'b00000;
assign A[16][170] = 5'b00010;
assign A[16][171] = 5'b11111;
assign A[16][172] = 5'b00000;
assign A[16][173] = 5'b11110;
assign A[16][174] = 5'b11111;
assign A[16][175] = 5'b00010;
assign A[16][176] = 5'b00001;
assign A[16][177] = 5'b00010;
assign A[16][178] = 5'b11110;
assign A[16][179] = 5'b00001;
assign A[16][180] = 5'b00000;
assign A[16][181] = 5'b00011;
assign A[16][182] = 5'b00001;
assign A[16][183] = 5'b00000;
assign A[16][184] = 5'b11110;
assign A[16][185] = 5'b11111;
assign A[16][186] = 5'b00001;
assign A[16][187] = 5'b00000;
assign A[16][188] = 5'b00000;
assign A[16][189] = 5'b11111;
assign A[16][190] = 5'b11110;
assign A[16][191] = 5'b00001;
assign A[16][192] = 5'b11111;
assign A[16][193] = 5'b00000;
assign A[16][194] = 5'b11110;
assign A[16][195] = 5'b00010;
assign A[16][196] = 5'b11110;
assign A[16][197] = 5'b00000;
assign A[16][198] = 5'b11111;
assign A[16][199] = 5'b00001;
assign A[16][200] = 5'b11110;
assign A[16][201] = 5'b00000;
assign A[16][202] = 5'b11101;
assign A[16][203] = 5'b11111;
assign A[16][204] = 5'b11110;
assign A[16][205] = 5'b11111;
assign A[16][206] = 5'b11111;
assign A[16][207] = 5'b00000;
assign A[16][208] = 5'b00000;
assign A[16][209] = 5'b00001;
assign A[16][210] = 5'b00000;
assign A[16][211] = 5'b00010;
assign A[16][212] = 5'b00001;
assign A[16][213] = 5'b11101;
assign A[16][214] = 5'b00010;
assign A[16][215] = 5'b00001;
assign A[16][216] = 5'b11110;
assign A[16][217] = 5'b11111;
assign A[16][218] = 5'b11110;
assign A[16][219] = 5'b00000;
assign A[16][220] = 5'b00001;
assign A[16][221] = 5'b00000;
assign A[16][222] = 5'b11111;
assign A[16][223] = 5'b11110;
assign A[16][224] = 5'b00000;
assign A[16][225] = 5'b00000;
assign A[16][226] = 5'b00000;
assign A[16][227] = 5'b00000;
assign A[16][228] = 5'b00000;
assign A[16][229] = 5'b00000;
assign A[16][230] = 5'b00010;
assign A[16][231] = 5'b00001;
assign A[16][232] = 5'b00000;
assign A[16][233] = 5'b11110;
assign A[16][234] = 5'b00010;
assign A[16][235] = 5'b11111;
assign A[16][236] = 5'b11111;
assign A[16][237] = 5'b00000;
assign A[16][238] = 5'b00000;
assign A[16][239] = 5'b11101;
assign A[16][240] = 5'b00000;
assign A[16][241] = 5'b11110;
assign A[16][242] = 5'b11110;
assign A[16][243] = 5'b11111;
assign A[16][244] = 5'b11111;
assign A[16][245] = 5'b11110;
assign A[16][246] = 5'b00001;
assign A[16][247] = 5'b00001;
assign A[16][248] = 5'b00000;
assign A[16][249] = 5'b00010;
assign A[16][250] = 5'b00000;
assign A[16][251] = 5'b00010;
assign A[16][252] = 5'b00010;
assign A[16][253] = 5'b00001;
assign A[16][254] = 5'b00001;
assign A[16][255] = 5'b00000;
assign A[17][0] = 5'b11111;
assign A[17][1] = 5'b11101;
assign A[17][2] = 5'b00010;
assign A[17][3] = 5'b00001;
assign A[17][4] = 5'b11101;
assign A[17][5] = 5'b11100;
assign A[17][6] = 5'b00010;
assign A[17][7] = 5'b00110;
assign A[17][8] = 5'b00000;
assign A[17][9] = 5'b11110;
assign A[17][10] = 5'b00000;
assign A[17][11] = 5'b11101;
assign A[17][12] = 5'b11101;
assign A[17][13] = 5'b11111;
assign A[17][14] = 5'b11110;
assign A[17][15] = 5'b11011;
assign A[17][16] = 5'b00000;
assign A[17][17] = 5'b00000;
assign A[17][18] = 5'b00010;
assign A[17][19] = 5'b11111;
assign A[17][20] = 5'b00000;
assign A[17][21] = 5'b00001;
assign A[17][22] = 5'b00010;
assign A[17][23] = 5'b00001;
assign A[17][24] = 5'b11110;
assign A[17][25] = 5'b00001;
assign A[17][26] = 5'b00001;
assign A[17][27] = 5'b00010;
assign A[17][28] = 5'b11110;
assign A[17][29] = 5'b00001;
assign A[17][30] = 5'b00010;
assign A[17][31] = 5'b11111;
assign A[17][32] = 5'b11111;
assign A[17][33] = 5'b11111;
assign A[17][34] = 5'b00000;
assign A[17][35] = 5'b11111;
assign A[17][36] = 5'b11110;
assign A[17][37] = 5'b11111;
assign A[17][38] = 5'b00000;
assign A[17][39] = 5'b11111;
assign A[17][40] = 5'b00000;
assign A[17][41] = 5'b11111;
assign A[17][42] = 5'b00010;
assign A[17][43] = 5'b11110;
assign A[17][44] = 5'b00001;
assign A[17][45] = 5'b11101;
assign A[17][46] = 5'b00001;
assign A[17][47] = 5'b00101;
assign A[17][48] = 5'b11111;
assign A[17][49] = 5'b11101;
assign A[17][50] = 5'b00001;
assign A[17][51] = 5'b11110;
assign A[17][52] = 5'b11110;
assign A[17][53] = 5'b11110;
assign A[17][54] = 5'b11111;
assign A[17][55] = 5'b00100;
assign A[17][56] = 5'b00000;
assign A[17][57] = 5'b00010;
assign A[17][58] = 5'b11111;
assign A[17][59] = 5'b00001;
assign A[17][60] = 5'b00001;
assign A[17][61] = 5'b11111;
assign A[17][62] = 5'b00010;
assign A[17][63] = 5'b00011;
assign A[17][64] = 5'b00000;
assign A[17][65] = 5'b11100;
assign A[17][66] = 5'b11101;
assign A[17][67] = 5'b00010;
assign A[17][68] = 5'b00000;
assign A[17][69] = 5'b00001;
assign A[17][70] = 5'b00001;
assign A[17][71] = 5'b00001;
assign A[17][72] = 5'b11110;
assign A[17][73] = 5'b11111;
assign A[17][74] = 5'b00010;
assign A[17][75] = 5'b00000;
assign A[17][76] = 5'b00101;
assign A[17][77] = 5'b11111;
assign A[17][78] = 5'b00100;
assign A[17][79] = 5'b00000;
assign A[17][80] = 5'b11111;
assign A[17][81] = 5'b11110;
assign A[17][82] = 5'b00000;
assign A[17][83] = 5'b11111;
assign A[17][84] = 5'b11110;
assign A[17][85] = 5'b00001;
assign A[17][86] = 5'b00001;
assign A[17][87] = 5'b11111;
assign A[17][88] = 5'b00100;
assign A[17][89] = 5'b00001;
assign A[17][90] = 5'b00000;
assign A[17][91] = 5'b00000;
assign A[17][92] = 5'b11110;
assign A[17][93] = 5'b00001;
assign A[17][94] = 5'b11110;
assign A[17][95] = 5'b00000;
assign A[17][96] = 5'b00000;
assign A[17][97] = 5'b00000;
assign A[17][98] = 5'b00010;
assign A[17][99] = 5'b11110;
assign A[17][100] = 5'b00010;
assign A[17][101] = 5'b11101;
assign A[17][102] = 5'b11101;
assign A[17][103] = 5'b00000;
assign A[17][104] = 5'b00010;
assign A[17][105] = 5'b11111;
assign A[17][106] = 5'b00000;
assign A[17][107] = 5'b00000;
assign A[17][108] = 5'b00010;
assign A[17][109] = 5'b11110;
assign A[17][110] = 5'b11110;
assign A[17][111] = 5'b00000;
assign A[17][112] = 5'b11100;
assign A[17][113] = 5'b11110;
assign A[17][114] = 5'b00000;
assign A[17][115] = 5'b11111;
assign A[17][116] = 5'b00000;
assign A[17][117] = 5'b11110;
assign A[17][118] = 5'b11111;
assign A[17][119] = 5'b00010;
assign A[17][120] = 5'b11101;
assign A[17][121] = 5'b00001;
assign A[17][122] = 5'b11111;
assign A[17][123] = 5'b00000;
assign A[17][124] = 5'b11111;
assign A[17][125] = 5'b11101;
assign A[17][126] = 5'b11110;
assign A[17][127] = 5'b11110;
assign A[17][128] = 5'b11110;
assign A[17][129] = 5'b11111;
assign A[17][130] = 5'b00001;
assign A[17][131] = 5'b00001;
assign A[17][132] = 5'b00010;
assign A[17][133] = 5'b11110;
assign A[17][134] = 5'b11111;
assign A[17][135] = 5'b00000;
assign A[17][136] = 5'b11111;
assign A[17][137] = 5'b00010;
assign A[17][138] = 5'b00000;
assign A[17][139] = 5'b11110;
assign A[17][140] = 5'b00001;
assign A[17][141] = 5'b00000;
assign A[17][142] = 5'b11111;
assign A[17][143] = 5'b11110;
assign A[17][144] = 5'b00000;
assign A[17][145] = 5'b11110;
assign A[17][146] = 5'b11111;
assign A[17][147] = 5'b00000;
assign A[17][148] = 5'b11011;
assign A[17][149] = 5'b11111;
assign A[17][150] = 5'b00001;
assign A[17][151] = 5'b00010;
assign A[17][152] = 5'b11110;
assign A[17][153] = 5'b00001;
assign A[17][154] = 5'b11111;
assign A[17][155] = 5'b00000;
assign A[17][156] = 5'b11100;
assign A[17][157] = 5'b00001;
assign A[17][158] = 5'b11110;
assign A[17][159] = 5'b11111;
assign A[17][160] = 5'b00000;
assign A[17][161] = 5'b00001;
assign A[17][162] = 5'b00010;
assign A[17][163] = 5'b00011;
assign A[17][164] = 5'b00001;
assign A[17][165] = 5'b00010;
assign A[17][166] = 5'b11111;
assign A[17][167] = 5'b00000;
assign A[17][168] = 5'b11110;
assign A[17][169] = 5'b11111;
assign A[17][170] = 5'b00001;
assign A[17][171] = 5'b11100;
assign A[17][172] = 5'b11110;
assign A[17][173] = 5'b00000;
assign A[17][174] = 5'b00001;
assign A[17][175] = 5'b11111;
assign A[17][176] = 5'b00000;
assign A[17][177] = 5'b11101;
assign A[17][178] = 5'b00001;
assign A[17][179] = 5'b00000;
assign A[17][180] = 5'b11111;
assign A[17][181] = 5'b00001;
assign A[17][182] = 5'b00011;
assign A[17][183] = 5'b00001;
assign A[17][184] = 5'b00000;
assign A[17][185] = 5'b11111;
assign A[17][186] = 5'b11101;
assign A[17][187] = 5'b11111;
assign A[17][188] = 5'b11110;
assign A[17][189] = 5'b00001;
assign A[17][190] = 5'b00000;
assign A[17][191] = 5'b00010;
assign A[17][192] = 5'b00001;
assign A[17][193] = 5'b00000;
assign A[17][194] = 5'b11111;
assign A[17][195] = 5'b00001;
assign A[17][196] = 5'b11111;
assign A[17][197] = 5'b00000;
assign A[17][198] = 5'b00000;
assign A[17][199] = 5'b11101;
assign A[17][200] = 5'b11110;
assign A[17][201] = 5'b11111;
assign A[17][202] = 5'b00000;
assign A[17][203] = 5'b00010;
assign A[17][204] = 5'b00010;
assign A[17][205] = 5'b00000;
assign A[17][206] = 5'b00000;
assign A[17][207] = 5'b00001;
assign A[17][208] = 5'b00101;
assign A[17][209] = 5'b11111;
assign A[17][210] = 5'b00000;
assign A[17][211] = 5'b11111;
assign A[17][212] = 5'b00010;
assign A[17][213] = 5'b11110;
assign A[17][214] = 5'b00000;
assign A[17][215] = 5'b11111;
assign A[17][216] = 5'b00000;
assign A[17][217] = 5'b00000;
assign A[17][218] = 5'b00000;
assign A[17][219] = 5'b00011;
assign A[17][220] = 5'b11110;
assign A[17][221] = 5'b00001;
assign A[17][222] = 5'b00101;
assign A[17][223] = 5'b11111;
assign A[17][224] = 5'b00001;
assign A[17][225] = 5'b11110;
assign A[17][226] = 5'b00000;
assign A[17][227] = 5'b00000;
assign A[17][228] = 5'b00000;
assign A[17][229] = 5'b00010;
assign A[17][230] = 5'b11101;
assign A[17][231] = 5'b00001;
assign A[17][232] = 5'b00001;
assign A[17][233] = 5'b00010;
assign A[17][234] = 5'b00001;
assign A[17][235] = 5'b00010;
assign A[17][236] = 5'b00001;
assign A[17][237] = 5'b00100;
assign A[17][238] = 5'b11110;
assign A[17][239] = 5'b00001;
assign A[17][240] = 5'b00010;
assign A[17][241] = 5'b00001;
assign A[17][242] = 5'b00000;
assign A[17][243] = 5'b00000;
assign A[17][244] = 5'b00000;
assign A[17][245] = 5'b11111;
assign A[17][246] = 5'b11110;
assign A[17][247] = 5'b00000;
assign A[17][248] = 5'b11110;
assign A[17][249] = 5'b11100;
assign A[17][250] = 5'b00010;
assign A[17][251] = 5'b00011;
assign A[17][252] = 5'b00001;
assign A[17][253] = 5'b00010;
assign A[17][254] = 5'b00001;
assign A[17][255] = 5'b11111;
assign A[18][0] = 5'b00001;
assign A[18][1] = 5'b00011;
assign A[18][2] = 5'b00001;
assign A[18][3] = 5'b00001;
assign A[18][4] = 5'b00000;
assign A[18][5] = 5'b00000;
assign A[18][6] = 5'b00000;
assign A[18][7] = 5'b11111;
assign A[18][8] = 5'b00000;
assign A[18][9] = 5'b00001;
assign A[18][10] = 5'b00010;
assign A[18][11] = 5'b00000;
assign A[18][12] = 5'b00010;
assign A[18][13] = 5'b11111;
assign A[18][14] = 5'b11110;
assign A[18][15] = 5'b00001;
assign A[18][16] = 5'b11101;
assign A[18][17] = 5'b00010;
assign A[18][18] = 5'b11111;
assign A[18][19] = 5'b00010;
assign A[18][20] = 5'b00000;
assign A[18][21] = 5'b00001;
assign A[18][22] = 5'b11111;
assign A[18][23] = 5'b00000;
assign A[18][24] = 5'b00010;
assign A[18][25] = 5'b00011;
assign A[18][26] = 5'b00000;
assign A[18][27] = 5'b00000;
assign A[18][28] = 5'b11111;
assign A[18][29] = 5'b00000;
assign A[18][30] = 5'b00100;
assign A[18][31] = 5'b11110;
assign A[18][32] = 5'b11111;
assign A[18][33] = 5'b11101;
assign A[18][34] = 5'b11111;
assign A[18][35] = 5'b11111;
assign A[18][36] = 5'b11110;
assign A[18][37] = 5'b11101;
assign A[18][38] = 5'b00000;
assign A[18][39] = 5'b00000;
assign A[18][40] = 5'b11111;
assign A[18][41] = 5'b11110;
assign A[18][42] = 5'b00010;
assign A[18][43] = 5'b00010;
assign A[18][44] = 5'b00001;
assign A[18][45] = 5'b00001;
assign A[18][46] = 5'b00000;
assign A[18][47] = 5'b00100;
assign A[18][48] = 5'b00011;
assign A[18][49] = 5'b00000;
assign A[18][50] = 5'b11110;
assign A[18][51] = 5'b00001;
assign A[18][52] = 5'b11111;
assign A[18][53] = 5'b00000;
assign A[18][54] = 5'b11110;
assign A[18][55] = 5'b11111;
assign A[18][56] = 5'b00001;
assign A[18][57] = 5'b00001;
assign A[18][58] = 5'b00100;
assign A[18][59] = 5'b00000;
assign A[18][60] = 5'b00001;
assign A[18][61] = 5'b00001;
assign A[18][62] = 5'b00001;
assign A[18][63] = 5'b00001;
assign A[18][64] = 5'b11110;
assign A[18][65] = 5'b11111;
assign A[18][66] = 5'b11100;
assign A[18][67] = 5'b00000;
assign A[18][68] = 5'b00001;
assign A[18][69] = 5'b00001;
assign A[18][70] = 5'b00000;
assign A[18][71] = 5'b11111;
assign A[18][72] = 5'b11111;
assign A[18][73] = 5'b11110;
assign A[18][74] = 5'b00000;
assign A[18][75] = 5'b11111;
assign A[18][76] = 5'b00001;
assign A[18][77] = 5'b11111;
assign A[18][78] = 5'b00010;
assign A[18][79] = 5'b11111;
assign A[18][80] = 5'b00001;
assign A[18][81] = 5'b00001;
assign A[18][82] = 5'b00000;
assign A[18][83] = 5'b11111;
assign A[18][84] = 5'b11111;
assign A[18][85] = 5'b00000;
assign A[18][86] = 5'b00001;
assign A[18][87] = 5'b00000;
assign A[18][88] = 5'b11110;
assign A[18][89] = 5'b11100;
assign A[18][90] = 5'b11111;
assign A[18][91] = 5'b11101;
assign A[18][92] = 5'b11110;
assign A[18][93] = 5'b11110;
assign A[18][94] = 5'b00000;
assign A[18][95] = 5'b00011;
assign A[18][96] = 5'b11111;
assign A[18][97] = 5'b00001;
assign A[18][98] = 5'b11111;
assign A[18][99] = 5'b11110;
assign A[18][100] = 5'b11111;
assign A[18][101] = 5'b00000;
assign A[18][102] = 5'b00000;
assign A[18][103] = 5'b11101;
assign A[18][104] = 5'b11110;
assign A[18][105] = 5'b11110;
assign A[18][106] = 5'b00001;
assign A[18][107] = 5'b00000;
assign A[18][108] = 5'b11111;
assign A[18][109] = 5'b00000;
assign A[18][110] = 5'b00011;
assign A[18][111] = 5'b00001;
assign A[18][112] = 5'b00011;
assign A[18][113] = 5'b00001;
assign A[18][114] = 5'b11110;
assign A[18][115] = 5'b00000;
assign A[18][116] = 5'b00001;
assign A[18][117] = 5'b11110;
assign A[18][118] = 5'b11111;
assign A[18][119] = 5'b00000;
assign A[18][120] = 5'b00000;
assign A[18][121] = 5'b00000;
assign A[18][122] = 5'b11101;
assign A[18][123] = 5'b11110;
assign A[18][124] = 5'b11110;
assign A[18][125] = 5'b00010;
assign A[18][126] = 5'b00101;
assign A[18][127] = 5'b11111;
assign A[18][128] = 5'b11111;
assign A[18][129] = 5'b00011;
assign A[18][130] = 5'b00001;
assign A[18][131] = 5'b11101;
assign A[18][132] = 5'b11101;
assign A[18][133] = 5'b11111;
assign A[18][134] = 5'b11111;
assign A[18][135] = 5'b11111;
assign A[18][136] = 5'b00001;
assign A[18][137] = 5'b11111;
assign A[18][138] = 5'b11111;
assign A[18][139] = 5'b11111;
assign A[18][140] = 5'b00000;
assign A[18][141] = 5'b11111;
assign A[18][142] = 5'b00001;
assign A[18][143] = 5'b00001;
assign A[18][144] = 5'b00001;
assign A[18][145] = 5'b00001;
assign A[18][146] = 5'b11111;
assign A[18][147] = 5'b00000;
assign A[18][148] = 5'b00001;
assign A[18][149] = 5'b11111;
assign A[18][150] = 5'b00000;
assign A[18][151] = 5'b11101;
assign A[18][152] = 5'b11110;
assign A[18][153] = 5'b00011;
assign A[18][154] = 5'b00000;
assign A[18][155] = 5'b00010;
assign A[18][156] = 5'b11111;
assign A[18][157] = 5'b00001;
assign A[18][158] = 5'b00001;
assign A[18][159] = 5'b00100;
assign A[18][160] = 5'b00010;
assign A[18][161] = 5'b00000;
assign A[18][162] = 5'b00010;
assign A[18][163] = 5'b11110;
assign A[18][164] = 5'b00000;
assign A[18][165] = 5'b11101;
assign A[18][166] = 5'b11111;
assign A[18][167] = 5'b11101;
assign A[18][168] = 5'b00000;
assign A[18][169] = 5'b00000;
assign A[18][170] = 5'b00000;
assign A[18][171] = 5'b11101;
assign A[18][172] = 5'b11111;
assign A[18][173] = 5'b11111;
assign A[18][174] = 5'b00000;
assign A[18][175] = 5'b00001;
assign A[18][176] = 5'b11111;
assign A[18][177] = 5'b11101;
assign A[18][178] = 5'b00000;
assign A[18][179] = 5'b00001;
assign A[18][180] = 5'b00011;
assign A[18][181] = 5'b00010;
assign A[18][182] = 5'b00000;
assign A[18][183] = 5'b11110;
assign A[18][184] = 5'b00000;
assign A[18][185] = 5'b00010;
assign A[18][186] = 5'b00011;
assign A[18][187] = 5'b00000;
assign A[18][188] = 5'b11111;
assign A[18][189] = 5'b11111;
assign A[18][190] = 5'b00001;
assign A[18][191] = 5'b11111;
assign A[18][192] = 5'b00011;
assign A[18][193] = 5'b00000;
assign A[18][194] = 5'b11111;
assign A[18][195] = 5'b00000;
assign A[18][196] = 5'b00000;
assign A[18][197] = 5'b00001;
assign A[18][198] = 5'b00001;
assign A[18][199] = 5'b00001;
assign A[18][200] = 5'b00000;
assign A[18][201] = 5'b00001;
assign A[18][202] = 5'b00001;
assign A[18][203] = 5'b00010;
assign A[18][204] = 5'b00010;
assign A[18][205] = 5'b00001;
assign A[18][206] = 5'b11111;
assign A[18][207] = 5'b11111;
assign A[18][208] = 5'b00001;
assign A[18][209] = 5'b00011;
assign A[18][210] = 5'b00001;
assign A[18][211] = 5'b00010;
assign A[18][212] = 5'b00011;
assign A[18][213] = 5'b00000;
assign A[18][214] = 5'b11111;
assign A[18][215] = 5'b00011;
assign A[18][216] = 5'b00000;
assign A[18][217] = 5'b11111;
assign A[18][218] = 5'b00000;
assign A[18][219] = 5'b11110;
assign A[18][220] = 5'b00000;
assign A[18][221] = 5'b11111;
assign A[18][222] = 5'b00000;
assign A[18][223] = 5'b11110;
assign A[18][224] = 5'b00010;
assign A[18][225] = 5'b00010;
assign A[18][226] = 5'b00001;
assign A[18][227] = 5'b00000;
assign A[18][228] = 5'b11111;
assign A[18][229] = 5'b00010;
assign A[18][230] = 5'b11111;
assign A[18][231] = 5'b00011;
assign A[18][232] = 5'b00000;
assign A[18][233] = 5'b00010;
assign A[18][234] = 5'b00000;
assign A[18][235] = 5'b11110;
assign A[18][236] = 5'b00000;
assign A[18][237] = 5'b11110;
assign A[18][238] = 5'b11111;
assign A[18][239] = 5'b11111;
assign A[18][240] = 5'b00001;
assign A[18][241] = 5'b00010;
assign A[18][242] = 5'b00001;
assign A[18][243] = 5'b00000;
assign A[18][244] = 5'b11110;
assign A[18][245] = 5'b11111;
assign A[18][246] = 5'b00011;
assign A[18][247] = 5'b00010;
assign A[18][248] = 5'b00000;
assign A[18][249] = 5'b00000;
assign A[18][250] = 5'b11111;
assign A[18][251] = 5'b00001;
assign A[18][252] = 5'b00000;
assign A[18][253] = 5'b11111;
assign A[18][254] = 5'b11111;
assign A[18][255] = 5'b00001;
assign A[19][0] = 5'b00100;
assign A[19][1] = 5'b11111;
assign A[19][2] = 5'b00011;
assign A[19][3] = 5'b00001;
assign A[19][4] = 5'b11111;
assign A[19][5] = 5'b00001;
assign A[19][6] = 5'b00100;
assign A[19][7] = 5'b00010;
assign A[19][8] = 5'b00000;
assign A[19][9] = 5'b00000;
assign A[19][10] = 5'b00000;
assign A[19][11] = 5'b00010;
assign A[19][12] = 5'b00011;
assign A[19][13] = 5'b00001;
assign A[19][14] = 5'b00000;
assign A[19][15] = 5'b00100;
assign A[19][16] = 5'b00001;
assign A[19][17] = 5'b11110;
assign A[19][18] = 5'b00001;
assign A[19][19] = 5'b00001;
assign A[19][20] = 5'b00000;
assign A[19][21] = 5'b00010;
assign A[19][22] = 5'b00010;
assign A[19][23] = 5'b11111;
assign A[19][24] = 5'b00001;
assign A[19][25] = 5'b00010;
assign A[19][26] = 5'b11100;
assign A[19][27] = 5'b00010;
assign A[19][28] = 5'b11111;
assign A[19][29] = 5'b11111;
assign A[19][30] = 5'b00001;
assign A[19][31] = 5'b11101;
assign A[19][32] = 5'b00001;
assign A[19][33] = 5'b11111;
assign A[19][34] = 5'b11111;
assign A[19][35] = 5'b00000;
assign A[19][36] = 5'b00001;
assign A[19][37] = 5'b11101;
assign A[19][38] = 5'b00000;
assign A[19][39] = 5'b00100;
assign A[19][40] = 5'b00000;
assign A[19][41] = 5'b11111;
assign A[19][42] = 5'b00000;
assign A[19][43] = 5'b00000;
assign A[19][44] = 5'b11101;
assign A[19][45] = 5'b00010;
assign A[19][46] = 5'b11100;
assign A[19][47] = 5'b11110;
assign A[19][48] = 5'b11110;
assign A[19][49] = 5'b11110;
assign A[19][50] = 5'b00000;
assign A[19][51] = 5'b00000;
assign A[19][52] = 5'b11111;
assign A[19][53] = 5'b00000;
assign A[19][54] = 5'b11110;
assign A[19][55] = 5'b00000;
assign A[19][56] = 5'b11101;
assign A[19][57] = 5'b11100;
assign A[19][58] = 5'b11110;
assign A[19][59] = 5'b11010;
assign A[19][60] = 5'b11100;
assign A[19][61] = 5'b11110;
assign A[19][62] = 5'b11110;
assign A[19][63] = 5'b00000;
assign A[19][64] = 5'b00000;
assign A[19][65] = 5'b11111;
assign A[19][66] = 5'b11111;
assign A[19][67] = 5'b00000;
assign A[19][68] = 5'b11111;
assign A[19][69] = 5'b11111;
assign A[19][70] = 5'b11111;
assign A[19][71] = 5'b11111;
assign A[19][72] = 5'b11111;
assign A[19][73] = 5'b11101;
assign A[19][74] = 5'b00010;
assign A[19][75] = 5'b11111;
assign A[19][76] = 5'b11101;
assign A[19][77] = 5'b11011;
assign A[19][78] = 5'b11001;
assign A[19][79] = 5'b11011;
assign A[19][80] = 5'b11110;
assign A[19][81] = 5'b11111;
assign A[19][82] = 5'b11100;
assign A[19][83] = 5'b11110;
assign A[19][84] = 5'b00001;
assign A[19][85] = 5'b11111;
assign A[19][86] = 5'b00010;
assign A[19][87] = 5'b11011;
assign A[19][88] = 5'b11111;
assign A[19][89] = 5'b00000;
assign A[19][90] = 5'b11111;
assign A[19][91] = 5'b11110;
assign A[19][92] = 5'b11111;
assign A[19][93] = 5'b11110;
assign A[19][94] = 5'b11000;
assign A[19][95] = 5'b11100;
assign A[19][96] = 5'b11111;
assign A[19][97] = 5'b00001;
assign A[19][98] = 5'b00000;
assign A[19][99] = 5'b00000;
assign A[19][100] = 5'b11110;
assign A[19][101] = 5'b00000;
assign A[19][102] = 5'b11111;
assign A[19][103] = 5'b00000;
assign A[19][104] = 5'b11111;
assign A[19][105] = 5'b00000;
assign A[19][106] = 5'b11111;
assign A[19][107] = 5'b00000;
assign A[19][108] = 5'b11111;
assign A[19][109] = 5'b00000;
assign A[19][110] = 5'b11100;
assign A[19][111] = 5'b11001;
assign A[19][112] = 5'b00000;
assign A[19][113] = 5'b00000;
assign A[19][114] = 5'b00001;
assign A[19][115] = 5'b11111;
assign A[19][116] = 5'b00000;
assign A[19][117] = 5'b00001;
assign A[19][118] = 5'b11111;
assign A[19][119] = 5'b11110;
assign A[19][120] = 5'b11110;
assign A[19][121] = 5'b00000;
assign A[19][122] = 5'b00000;
assign A[19][123] = 5'b11111;
assign A[19][124] = 5'b00000;
assign A[19][125] = 5'b00001;
assign A[19][126] = 5'b00000;
assign A[19][127] = 5'b11111;
assign A[19][128] = 5'b11101;
assign A[19][129] = 5'b00000;
assign A[19][130] = 5'b00001;
assign A[19][131] = 5'b00001;
assign A[19][132] = 5'b11110;
assign A[19][133] = 5'b11111;
assign A[19][134] = 5'b11110;
assign A[19][135] = 5'b00000;
assign A[19][136] = 5'b11110;
assign A[19][137] = 5'b00000;
assign A[19][138] = 5'b00011;
assign A[19][139] = 5'b11111;
assign A[19][140] = 5'b00001;
assign A[19][141] = 5'b11111;
assign A[19][142] = 5'b00000;
assign A[19][143] = 5'b11111;
assign A[19][144] = 5'b11011;
assign A[19][145] = 5'b11101;
assign A[19][146] = 5'b00001;
assign A[19][147] = 5'b11110;
assign A[19][148] = 5'b00000;
assign A[19][149] = 5'b00000;
assign A[19][150] = 5'b00001;
assign A[19][151] = 5'b11111;
assign A[19][152] = 5'b11111;
assign A[19][153] = 5'b00000;
assign A[19][154] = 5'b11111;
assign A[19][155] = 5'b11111;
assign A[19][156] = 5'b00000;
assign A[19][157] = 5'b11111;
assign A[19][158] = 5'b00000;
assign A[19][159] = 5'b00000;
assign A[19][160] = 5'b11110;
assign A[19][161] = 5'b11110;
assign A[19][162] = 5'b11111;
assign A[19][163] = 5'b00000;
assign A[19][164] = 5'b00000;
assign A[19][165] = 5'b00001;
assign A[19][166] = 5'b00000;
assign A[19][167] = 5'b00000;
assign A[19][168] = 5'b11111;
assign A[19][169] = 5'b00000;
assign A[19][170] = 5'b00001;
assign A[19][171] = 5'b00000;
assign A[19][172] = 5'b00000;
assign A[19][173] = 5'b11101;
assign A[19][174] = 5'b11110;
assign A[19][175] = 5'b00000;
assign A[19][176] = 5'b11110;
assign A[19][177] = 5'b00000;
assign A[19][178] = 5'b11110;
assign A[19][179] = 5'b11110;
assign A[19][180] = 5'b00000;
assign A[19][181] = 5'b11111;
assign A[19][182] = 5'b11111;
assign A[19][183] = 5'b11111;
assign A[19][184] = 5'b11101;
assign A[19][185] = 5'b00000;
assign A[19][186] = 5'b00000;
assign A[19][187] = 5'b00010;
assign A[19][188] = 5'b11110;
assign A[19][189] = 5'b00001;
assign A[19][190] = 5'b00010;
assign A[19][191] = 5'b00010;
assign A[19][192] = 5'b00010;
assign A[19][193] = 5'b00001;
assign A[19][194] = 5'b00000;
assign A[19][195] = 5'b11101;
assign A[19][196] = 5'b00000;
assign A[19][197] = 5'b11111;
assign A[19][198] = 5'b00010;
assign A[19][199] = 5'b11111;
assign A[19][200] = 5'b00000;
assign A[19][201] = 5'b11100;
assign A[19][202] = 5'b11110;
assign A[19][203] = 5'b00000;
assign A[19][204] = 5'b00001;
assign A[19][205] = 5'b00010;
assign A[19][206] = 5'b11111;
assign A[19][207] = 5'b00010;
assign A[19][208] = 5'b11111;
assign A[19][209] = 5'b00000;
assign A[19][210] = 5'b11110;
assign A[19][211] = 5'b00010;
assign A[19][212] = 5'b00001;
assign A[19][213] = 5'b00001;
assign A[19][214] = 5'b11110;
assign A[19][215] = 5'b00011;
assign A[19][216] = 5'b00000;
assign A[19][217] = 5'b00001;
assign A[19][218] = 5'b11111;
assign A[19][219] = 5'b11110;
assign A[19][220] = 5'b00000;
assign A[19][221] = 5'b11111;
assign A[19][222] = 5'b11111;
assign A[19][223] = 5'b00000;
assign A[19][224] = 5'b11110;
assign A[19][225] = 5'b00000;
assign A[19][226] = 5'b00000;
assign A[19][227] = 5'b00011;
assign A[19][228] = 5'b00000;
assign A[19][229] = 5'b11110;
assign A[19][230] = 5'b00000;
assign A[19][231] = 5'b00010;
assign A[19][232] = 5'b11101;
assign A[19][233] = 5'b00001;
assign A[19][234] = 5'b00010;
assign A[19][235] = 5'b11111;
assign A[19][236] = 5'b00001;
assign A[19][237] = 5'b00001;
assign A[19][238] = 5'b11101;
assign A[19][239] = 5'b00000;
assign A[19][240] = 5'b00000;
assign A[19][241] = 5'b00000;
assign A[19][242] = 5'b00010;
assign A[19][243] = 5'b00000;
assign A[19][244] = 5'b11110;
assign A[19][245] = 5'b00000;
assign A[19][246] = 5'b00001;
assign A[19][247] = 5'b00000;
assign A[19][248] = 5'b11101;
assign A[19][249] = 5'b00000;
assign A[19][250] = 5'b00001;
assign A[19][251] = 5'b00000;
assign A[19][252] = 5'b00001;
assign A[19][253] = 5'b11110;
assign A[19][254] = 5'b11111;
assign A[19][255] = 5'b00000;




    // reg [6:0] biases_l1 [0:19];
    // initial begin
    //     $readmemb("b1.mem", biases_l1);
    // end

wire [6:0] biases_l1 [0:19];
assign biases_l1[0] = 7'b1110011;
assign biases_l1[1] = 7'b1111001;
assign biases_l1[2] = 7'b0010011;
assign biases_l1[3] = 7'b1111000;
assign biases_l1[4] = 7'b0001011;
assign biases_l1[5] = 7'b0000101;
assign biases_l1[6] = 7'b0000011;
assign biases_l1[7] = 7'b0001001;
assign biases_l1[8] = 7'b0011101;
assign biases_l1[9] = 7'b0010110;
assign biases_l1[10] = 7'b1100111;
assign biases_l1[11] = 7'b0000101;
assign biases_l1[12] = 7'b1101100;
assign biases_l1[13] = 7'b1100000;
assign biases_l1[14] = 7'b1101101;
assign biases_l1[15] = 7'b1011101;
assign biases_l1[16] = 7'b1101110;
assign biases_l1[17] = 7'b0010010;
assign biases_l1[18] = 7'b1111010;
assign biases_l1[19] = 7'b0101001;


    wire [9:0] biases_l1_ext [0:19];
    wire [5:0] level_1_sums [0:19][0:127]; // 128 outputs, each 6 bits wide
    wire [6:0] level_2_sums [0:19][0:63];  // 64 outputs, each 7 bits wide
    wire [7:0] level_3_sums [0:19][0:31];  // 32 outputs, each 8 bits wide
    wire [8:0] level_4_sums [0:19][0:15];  // 16 outputs, each 9 bits wide
    wire [9:0] level_5_sums [0:19][0:7];   // 8 outputs, each 10 bits wide
    wire [9:0] level_6_sums [0:19][0:3];   // 4 outputs, each 10 bits wide
    wire [9:0] level_7_sums [0:19][0:1];   // 2 outputs, each 10 bits wide
    wire [9:0] level_8_sums [0:19];        // 1 output, 10 bits wide
    wire [9:0] final_sums [0:19];          // Final output, 10 bits wide

    reg [8:0] out_reg [0:19];
    wire [8:0] out_sig [0:19];
    
    always @ (posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            B <= 256'd0;
        end

        else begin
            if(!updown) begin
                B <= {in, B[128:255]};
            end
            else begin
                B <= {B[0:127], in};
            end
        end
    end


    // --- Generate 20 Parallel Dot-Product Units ---
    genvar i, j;
    generate
        for (i = 0; i < 20; i = i + 1) begin : dot_product_and_ReLU
            assign biases_l1_ext[i] = { {3{biases_l1[i][6]}}, biases_l1[i] }; // Sign-extend 7-bit bias to 9 bits
            wire [4:0] product_terms [0:255]; // 256 products, each 5 bits wide            
            for (j = 0; j < 256; j = j + 1) begin : product_terms_gen
                assign product_terms[j] = B[j] ? A[i][j] : {5{1'b0}};
                if (j%2 == 1) begin : adder_pairs
                    // assign level_1_sums[i][j/2] = product_terms[j] + product_terms[j-1];
                    adder_5to6 adder_inst (
                        .a(product_terms[j-1]),
                        .b(product_terms[j]),
                        .sum(level_1_sums[i][j/2])
                    );
                end
                if (j%4 == 3) begin : adder_quads
                    adder_6to7 adder_inst (
                        .a(level_1_sums[i][(j-1)/2]),
                        .b(level_1_sums[i][(j-3)/2]),
                        .sum(level_2_sums[i][j/4])
                    );
                end
                if (j%8 == 7) begin : adder_octets
                    adder_7to8 adder_inst (
                        .a(level_2_sums[i][(j-1)/4]),
                        .b(level_2_sums[i][(j-7)/4]),
                        .sum(level_3_sums[i][j/8])
                    );
                end
                if (j%16 == 15) begin : adder_16s
                    adder_8to9 adder_inst (
                        .a(level_3_sums[i][(j-1)/8]),
                        .b(level_3_sums[i][(j-15)/8]),
                        .sum(level_4_sums[i][j/16])
                    );
                end
                if (j%32 == 31) begin : adder_32s
                    adder_9to10 adder_inst (
                        .a(level_4_sums[i][(j-1)/16]),
                        .b(level_4_sums[i][(j-31)/16]),
                        .sum(level_5_sums[i][j/32])
                    );
                end
                if (j%64 == 63) begin : adder_64s
                    adder_10to10 adder_inst (
                        .a(level_5_sums[i][(j-1)/32]),
                        .b(level_5_sums[i][(j-63)/32]),
                        .sum(level_6_sums[i][j/64])
                    );
                end
                if (j%128 == 127) begin : adder_128s
                    adder_10to10 adder_inst (
                        .a(level_6_sums[i][(j-1)/64]),
                        .b(level_6_sums[i][(j-127)/64]),
                        .sum(level_7_sums[i][j/128])
                    );
                end
                if (j == 255) begin : final_adder
                    adder_10to10 adder_inst (
                        .a(level_7_sums[i][0]),
                        .b(level_7_sums[i][1]),
                        .sum(level_8_sums[i])
                    );
                end    
            end 
            assign final_sums[i] = level_8_sums[i] + biases_l1_ext[i];
            // Apply ReLU activation
            ReLU_10bit relu_inst (
                //.clk(clk),
                //.rst_n(rst_n),
                .in_data(final_sums[i]),
                .out_data(out_sig[i])
            );  
        end        
    endgenerate
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            
    out_reg[0]  <= 9'd0;
    out_reg[1]  <= 9'd0;
    out_reg[2]  <= 9'd0;
    out_reg[3]  <= 9'd0;
    out_reg[4]  <= 9'd0;
    out_reg[5]  <= 9'd0;
    out_reg[6]  <= 9'd0;
    out_reg[7]  <= 9'd0;
    out_reg[8]  <= 9'd0;
    out_reg[9]  <= 9'd0;
    out_reg[10] <= 9'd0;
    out_reg[11] <= 9'd0;
    out_reg[12] <= 9'd0;
    out_reg[13] <= 9'd0;
    out_reg[14] <= 9'd0;
    out_reg[15] <= 9'd0;
    out_reg[16] <= 9'd0;
    out_reg[17] <= 9'd0;
    out_reg[18] <= 9'd0;
    out_reg[19] <= 9'd0;

        end else begin
            // for (integer i = 0; i < 20; i++) begin
            //     out_reg[i] <= out_sig[i];
            // end
out_reg[0]  <= out_sig[0];
out_reg[1]  <= out_sig[1];
out_reg[2]  <= out_sig[2];
out_reg[3]  <= out_sig[3];
out_reg[4]  <= out_sig[4];
out_reg[5]  <= out_sig[5];
out_reg[6]  <= out_sig[6];
out_reg[7]  <= out_sig[7];
out_reg[8]  <= out_sig[8];
out_reg[9]  <= out_sig[9];
out_reg[10] <= out_sig[10];
out_reg[11] <= out_sig[11];
out_reg[12] <= out_sig[12];
out_reg[13] <= out_sig[13];
out_reg[14] <= out_sig[14];
out_reg[15] <= out_sig[15];
out_reg[16] <= out_sig[16];
out_reg[17] <= out_sig[17];
out_reg[18] <= out_sig[18];
out_reg[19] <= out_sig[19];

        end
    end

    genvar m;
    generate
        for (m = 0; m < 20; m = m + 1) begin : output_assign
            assign out[(m+1)*9-1:m*9] = out_reg[m];
        end
    endgenerate
endmodule

module layer2(
    input  wire         clk,
    input  wire         rst_n,
    input  wire [179:0] in, // 180-bit input
    output wire  [179:0]  out // 180-bit final output
);

    // reg signed [4:0] w2 [0:9][0:19];
    // initial begin
    //     $readmemb("w2.mem", w2);
    // end

wire signed [4:0] w2 [0:9][0:19];
assign w2[0][0] = 5'b11110;
assign w2[0][1] = 5'b00011;
assign w2[0][2] = 5'b11101;
assign w2[0][3] = 5'b11101;
assign w2[0][4] = 5'b11010;
assign w2[0][5] = 5'b11101;
assign w2[0][6] = 5'b00001;
assign w2[0][7] = 5'b11110;
assign w2[0][8] = 5'b00000;
assign w2[0][9] = 5'b10111;
assign w2[0][10] = 5'b11110;
assign w2[0][11] = 5'b11111;
assign w2[0][12] = 5'b00001;
assign w2[0][13] = 5'b00001;
assign w2[0][14] = 5'b00011;
assign w2[0][15] = 5'b00010;
assign w2[0][16] = 5'b11111;
assign w2[0][17] = 5'b11101;
assign w2[0][18] = 5'b00100;
assign w2[0][19] = 5'b11011;
assign w2[1][0] = 5'b00100;
assign w2[1][1] = 5'b11101;
assign w2[1][2] = 5'b01001;
assign w2[1][3] = 5'b00101;
assign w2[1][4] = 5'b00101;
assign w2[1][5] = 5'b01010;
assign w2[1][6] = 5'b10111;
assign w2[1][7] = 5'b11110;
assign w2[1][8] = 5'b11110;
assign w2[1][9] = 5'b11110;
assign w2[1][10] = 5'b00101;
assign w2[1][11] = 5'b10110;
assign w2[1][12] = 5'b00100;
assign w2[1][13] = 5'b11011;
assign w2[1][14] = 5'b10011;
assign w2[1][15] = 5'b00111;
assign w2[1][16] = 5'b00111;
assign w2[1][17] = 5'b11101;
assign w2[1][18] = 5'b00010;
assign w2[1][19] = 5'b11100;
assign w2[2][0] = 5'b11011;
assign w2[2][1] = 5'b11111;
assign w2[2][2] = 5'b11000;
assign w2[2][3] = 5'b11111;
assign w2[2][4] = 5'b00010;
assign w2[2][5] = 5'b11110;
assign w2[2][6] = 5'b11010;
assign w2[2][7] = 5'b11110;
assign w2[2][8] = 5'b00101;
assign w2[2][9] = 5'b11100;
assign w2[2][10] = 5'b00101;
assign w2[2][11] = 5'b10101;
assign w2[2][12] = 5'b00000;
assign w2[2][13] = 5'b00111;
assign w2[2][14] = 5'b00001;
assign w2[2][15] = 5'b00000;
assign w2[2][16] = 5'b01011;
assign w2[2][17] = 5'b00100;
assign w2[2][18] = 5'b00000;
assign w2[2][19] = 5'b00001;
assign w2[3][0] = 5'b00001;
assign w2[3][1] = 5'b11100;
assign w2[3][2] = 5'b11000;
assign w2[3][3] = 5'b11000;
assign w2[3][4] = 5'b00010;
assign w2[3][5] = 5'b00010;
assign w2[3][6] = 5'b11100;
assign w2[3][7] = 5'b00011;
assign w2[3][8] = 5'b10111;
assign w2[3][9] = 5'b00011;
assign w2[3][10] = 5'b00000;
assign w2[3][11] = 5'b00010;
assign w2[3][12] = 5'b11100;
assign w2[3][13] = 5'b00000;
assign w2[3][14] = 5'b00101;
assign w2[3][15] = 5'b00000;
assign w2[3][16] = 5'b00001;
assign w2[3][17] = 5'b00101;
assign w2[3][18] = 5'b00111;
assign w2[3][19] = 5'b00100;
assign w2[4][0] = 5'b00000;
assign w2[4][1] = 5'b00010;
assign w2[4][2] = 5'b01010;
assign w2[4][3] = 5'b11101;
assign w2[4][4] = 5'b00100;
assign w2[4][5] = 5'b00010;
assign w2[4][6] = 5'b00101;
assign w2[4][7] = 5'b11100;
assign w2[4][8] = 5'b00001;
assign w2[4][9] = 5'b11110;
assign w2[4][10] = 5'b00000;
assign w2[4][11] = 5'b00101;
assign w2[4][12] = 5'b11001;
assign w2[4][13] = 5'b00001;
assign w2[4][14] = 5'b11111;
assign w2[4][15] = 5'b00010;
assign w2[4][16] = 5'b11110;
assign w2[4][17] = 5'b11111;
assign w2[4][18] = 5'b11100;
assign w2[4][19] = 5'b00010;
assign w2[5][0] = 5'b01000;
assign w2[5][1] = 5'b00010;
assign w2[5][2] = 5'b00001;
assign w2[5][3] = 5'b11111;
assign w2[5][4] = 5'b11100;
assign w2[5][5] = 5'b11100;
assign w2[5][6] = 5'b00010;
assign w2[5][7] = 5'b00000;
assign w2[5][8] = 5'b11110;
assign w2[5][9] = 5'b11100;
assign w2[5][10] = 5'b00100;
assign w2[5][11] = 5'b11100;
assign w2[5][12] = 5'b11101;
assign w2[5][13] = 5'b11100;
assign w2[5][14] = 5'b00011;
assign w2[5][15] = 5'b00111;
assign w2[5][16] = 5'b11110;
assign w2[5][17] = 5'b10110;
assign w2[5][18] = 5'b11100;
assign w2[5][19] = 5'b00111;
assign w2[6][0] = 5'b00010;
assign w2[6][1] = 5'b01001;
assign w2[6][2] = 5'b10110;
assign w2[6][3] = 5'b00001;
assign w2[6][4] = 5'b00001;
assign w2[6][5] = 5'b10110;
assign w2[6][6] = 5'b00000;
assign w2[6][7] = 5'b00011;
assign w2[6][8] = 5'b00011;
assign w2[6][9] = 5'b11100;
assign w2[6][10] = 5'b10111;
assign w2[6][11] = 5'b00110;
assign w2[6][12] = 5'b11001;
assign w2[6][13] = 5'b00011;
assign w2[6][14] = 5'b11100;
assign w2[6][15] = 5'b10011;
assign w2[6][16] = 5'b11111;
assign w2[6][17] = 5'b11110;
assign w2[6][18] = 5'b00001;
assign w2[6][19] = 5'b00001;
assign w2[7][0] = 5'b00000;
assign w2[7][1] = 5'b01001;
assign w2[7][2] = 5'b11111;
assign w2[7][3] = 5'b10111;
assign w2[7][4] = 5'b11001;
assign w2[7][5] = 5'b11001;
assign w2[7][6] = 5'b11010;
assign w2[7][7] = 5'b11111;
assign w2[7][8] = 5'b00101;
assign w2[7][9] = 5'b01001;
assign w2[7][10] = 5'b00000;
assign w2[7][11] = 5'b11110;
assign w2[7][12] = 5'b00110;
assign w2[7][13] = 5'b00000;
assign w2[7][14] = 5'b00001;
assign w2[7][15] = 5'b10111;
assign w2[7][16] = 5'b00100;
assign w2[7][17] = 5'b10111;
assign w2[7][18] = 5'b00011;
assign w2[7][19] = 5'b00000;
assign w2[8][0] = 5'b11001;
assign w2[8][1] = 5'b00100;
assign w2[8][2] = 5'b11100;
assign w2[8][3] = 5'b00010;
assign w2[8][4] = 5'b00000;
assign w2[8][5] = 5'b00001;
assign w2[8][6] = 5'b00010;
assign w2[8][7] = 5'b01010;
assign w2[8][8] = 5'b00011;
assign w2[8][9] = 5'b00001;
assign w2[8][10] = 5'b00000;
assign w2[8][11] = 5'b10100;
assign w2[8][12] = 5'b00000;
assign w2[8][13] = 5'b00010;
assign w2[8][14] = 5'b11101;
assign w2[8][15] = 5'b00110;
assign w2[8][16] = 5'b11111;
assign w2[8][17] = 5'b11111;
assign w2[8][18] = 5'b11010;
assign w2[8][19] = 5'b10011;
assign w2[9][0] = 5'b11000;
assign w2[9][1] = 5'b00110;
assign w2[9][2] = 5'b10111;
assign w2[9][3] = 5'b01001;
assign w2[9][4] = 5'b10111;
assign w2[9][5] = 5'b11111;
assign w2[9][6] = 5'b00100;
assign w2[9][7] = 5'b11100;
assign w2[9][8] = 5'b11011;
assign w2[9][9] = 5'b00001;
assign w2[9][10] = 5'b00010;
assign w2[9][11] = 5'b00000;
assign w2[9][12] = 5'b10111;
assign w2[9][13] = 5'b11110;
assign w2[9][14] = 5'b00101;
assign w2[9][15] = 5'b01001;
assign w2[9][16] = 5'b01010;
assign w2[9][17] = 5'b00011;
assign w2[9][18] = 5'b10111;
assign w2[9][19] = 5'b11011;


    // reg [5:0] biases_l2 [0:9];
    // initial begin
    //     $readmemb("b2.mem", biases_l2);
    // end

wire [5:0] biases_l2 [0:9];
assign biases_l2[0] = 6'b001001;
assign biases_l2[1] = 6'b001101;
assign biases_l2[2] = 6'b111110;
assign biases_l2[3] = 6'b111001;
assign biases_l2[4] = 6'b110001;
assign biases_l2[5] = 6'b000010;
assign biases_l2[6] = 6'b101101;
assign biases_l2[7] = 6'b110110;
assign biases_l2[8] = 6'b110001;
assign biases_l2[9] = 6'b000110;
    
    wire signed [13:0] prod_terms[0:9][0:19];
    wire signed [13:0] b2_extended [0:9];
    
    wire signed [18:0] row_sums [0:9];

    wire [17:0] row_output [0:9]; 
    reg [17:0] out_reg [0:9];

    
    genvar i,j;
    generate
        for (i = 0; i < 10; i = i + 1) begin : row_iteration

            assign b2_extended[i] = { {4{biases_l2[i][5]}}, biases_l2[i], 4'd0 };

            for (j = 0; j < 20; j = j + 1) begin : prod_calc
                //assign prod_terms[i][j] = $signed(in[(j+1)*9-1:j*9]) * w2[i][j]; 
                multiplier9514 mult_inst (.prod(prod_terms[i][j]), .num1($signed(in[(j+1)*9-1:j*9])), .num2(w2[i][j]));
            end
            
            assign row_sums[i] = prod_terms[i][0]  + prod_terms[i][1] + prod_terms[i][2]  +
                             prod_terms[i][3]  + prod_terms[i][4]  + prod_terms[i][5]  +
                             prod_terms[i][6]  + prod_terms[i][7]  + prod_terms[i][8]  +
                             prod_terms[i][9]  + prod_terms[i][10] + prod_terms[i][11] +
                             prod_terms[i][12] + prod_terms[i][13] + prod_terms[i][14] +
                             prod_terms[i][15] + prod_terms[i][16] + prod_terms[i][17] +
                             prod_terms[i][18] + prod_terms[i][19] + b2_extended[i];        
            //apply ReLU
            ReLU_19bit relu_inst (
                //.clk(clk),
                //.rst_n(rst_n),
                .in_data(row_sums[i]),
                .out_data(row_output[i])
            );  
        end
    endgenerate

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // for (integer i = 0; i < 10; i++) begin
            //     out_reg[i] <= 18'd0;
            // end
out_reg[0] <= 18'd0;
out_reg[1] <= 18'd0;
out_reg[2] <= 18'd0;
out_reg[3] <= 18'd0;
out_reg[4] <= 18'd0;
out_reg[5] <= 18'd0;
out_reg[6] <= 18'd0;
out_reg[7] <= 18'd0;
out_reg[8] <= 18'd0;
out_reg[9] <= 18'd0;

        end else begin
            // for (integer i = 0; i < 10; i++) begin
            //     out_reg[i] <= row_output[i];
            // end
out_reg[0] <= row_output[0];
out_reg[1] <= row_output[1];
out_reg[2] <= row_output[2];
out_reg[3] <= row_output[3];
out_reg[4] <= row_output[4];
out_reg[5] <= row_output[5];
out_reg[6] <= row_output[6];
out_reg[7] <= row_output[7];
out_reg[8] <= row_output[8];
out_reg[9] <= row_output[9];

        end
    end

    genvar m;
    generate
        for (m = 0; m < 10; m = m + 1) begin : output_assign
            assign out[(m+1)*18-1:m*18] = out_reg[m];
        end
    endgenerate

endmodule

module mytop (
input wire [127:0] in,
input wire clk, 
input wire rst_n,
input wire updown,
//output wire [3:0] out,
output wire [0:9] out_activehigh,
output reg done
//output wire [17:0] max
);

wire [179:0] layer1_out;

reg [1:0] counter;

always @ (posedge clk or negedge updown) begin
if(!updown)begin
    counter <= 0;
    done <= 0;
end

else begin
    
    if (counter < 3) begin
        //done <=1;
        counter <= counter + 1;
        //counter <= 0;
    end    
    else begin
        done <=1;
    end

end
end


layer1 instanceL1 (
        .clk(clk),
        .rst_n(rst_n),
        .updown(updown),
        .in(in),
        .out(layer1_out)
    );

wire [179:0] layer2_out;

layer2 instanceL2 (
        .clk(clk),
        .rst_n(rst_n),
        .in(layer1_out),
        .out(layer2_out)
    );

wire [3:0] out;
wire [17:0] max;

find_max_index uut (
        .data_in(layer2_out),
        .clk(clk),
        .rst_n(rst_n),
        .max_index(out),
        .max_value(max)
    );

decoder_4_to_10 dut (
        .in_val(out),
        .out_activehigh(out_activehigh)
    );
endmodule

